// This is the unpowered netlist.
module wrapped_as1802 (clk,
    io_oeb,
    rst,
    io_in,
    io_out);
 input clk;
 output io_oeb;
 input rst;
 input [12:0] io_in;
 output [26:0] io_out;

 wire net285;
 wire net286;
 wire net287;
 wire net283;
 wire net284;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire \as1802.DF ;
 wire \as1802.D[0] ;
 wire \as1802.D[1] ;
 wire \as1802.D[2] ;
 wire \as1802.D[3] ;
 wire \as1802.D[4] ;
 wire \as1802.D[5] ;
 wire \as1802.D[6] ;
 wire \as1802.D[7] ;
 wire \as1802.EF_l[0] ;
 wire \as1802.EF_l[1] ;
 wire \as1802.EF_l[2] ;
 wire \as1802.EF_l[3] ;
 wire \as1802.IE ;
 wire \as1802.P[0] ;
 wire \as1802.P[1] ;
 wire \as1802.P[2] ;
 wire \as1802.P[3] ;
 wire \as1802.T[0] ;
 wire \as1802.T[1] ;
 wire \as1802.T[2] ;
 wire \as1802.T[3] ;
 wire \as1802.T[4] ;
 wire \as1802.T[5] ;
 wire \as1802.T[6] ;
 wire \as1802.T[7] ;
 wire \as1802.X[0] ;
 wire \as1802.X[1] ;
 wire \as1802.X[2] ;
 wire \as1802.X[3] ;
 wire \as1802.addr_buff[0] ;
 wire \as1802.addr_buff[10] ;
 wire \as1802.addr_buff[11] ;
 wire \as1802.addr_buff[12] ;
 wire \as1802.addr_buff[13] ;
 wire \as1802.addr_buff[14] ;
 wire \as1802.addr_buff[15] ;
 wire \as1802.addr_buff[1] ;
 wire \as1802.addr_buff[2] ;
 wire \as1802.addr_buff[3] ;
 wire \as1802.addr_buff[4] ;
 wire \as1802.addr_buff[5] ;
 wire \as1802.addr_buff[6] ;
 wire \as1802.addr_buff[7] ;
 wire \as1802.addr_buff[8] ;
 wire \as1802.addr_buff[9] ;
 wire \as1802.cond_inv ;
 wire \as1802.idle ;
 wire \as1802.instr_cycle[0] ;
 wire \as1802.instr_cycle[1] ;
 wire \as1802.instr_cycle[2] ;
 wire \as1802.instr_cycle[3] ;
 wire \as1802.instr_latch[0] ;
 wire \as1802.instr_latch[1] ;
 wire \as1802.instr_latch[2] ;
 wire \as1802.instr_latch[4] ;
 wire \as1802.instr_latch[5] ;
 wire \as1802.instr_latch[6] ;
 wire \as1802.instr_latch[7] ;
 wire \as1802.last_hi_addr[0] ;
 wire \as1802.last_hi_addr[1] ;
 wire \as1802.last_hi_addr[2] ;
 wire \as1802.last_hi_addr[3] ;
 wire \as1802.last_hi_addr[4] ;
 wire \as1802.last_hi_addr[5] ;
 wire \as1802.last_hi_addr[6] ;
 wire \as1802.last_hi_addr[7] ;
 wire \as1802.lda ;
 wire \as1802.mem_cycle[0] ;
 wire \as1802.mem_cycle[1] ;
 wire \as1802.mem_cycle[2] ;
 wire \as1802.mem_write ;
 wire \as1802.regs[0][0] ;
 wire \as1802.regs[0][10] ;
 wire \as1802.regs[0][11] ;
 wire \as1802.regs[0][12] ;
 wire \as1802.regs[0][13] ;
 wire \as1802.regs[0][14] ;
 wire \as1802.regs[0][15] ;
 wire \as1802.regs[0][1] ;
 wire \as1802.regs[0][2] ;
 wire \as1802.regs[0][3] ;
 wire \as1802.regs[0][4] ;
 wire \as1802.regs[0][5] ;
 wire \as1802.regs[0][6] ;
 wire \as1802.regs[0][7] ;
 wire \as1802.regs[0][8] ;
 wire \as1802.regs[0][9] ;
 wire \as1802.regs[10][0] ;
 wire \as1802.regs[10][10] ;
 wire \as1802.regs[10][11] ;
 wire \as1802.regs[10][12] ;
 wire \as1802.regs[10][13] ;
 wire \as1802.regs[10][14] ;
 wire \as1802.regs[10][15] ;
 wire \as1802.regs[10][1] ;
 wire \as1802.regs[10][2] ;
 wire \as1802.regs[10][3] ;
 wire \as1802.regs[10][4] ;
 wire \as1802.regs[10][5] ;
 wire \as1802.regs[10][6] ;
 wire \as1802.regs[10][7] ;
 wire \as1802.regs[10][8] ;
 wire \as1802.regs[10][9] ;
 wire \as1802.regs[11][0] ;
 wire \as1802.regs[11][10] ;
 wire \as1802.regs[11][11] ;
 wire \as1802.regs[11][12] ;
 wire \as1802.regs[11][13] ;
 wire \as1802.regs[11][14] ;
 wire \as1802.regs[11][15] ;
 wire \as1802.regs[11][1] ;
 wire \as1802.regs[11][2] ;
 wire \as1802.regs[11][3] ;
 wire \as1802.regs[11][4] ;
 wire \as1802.regs[11][5] ;
 wire \as1802.regs[11][6] ;
 wire \as1802.regs[11][7] ;
 wire \as1802.regs[11][8] ;
 wire \as1802.regs[11][9] ;
 wire \as1802.regs[12][0] ;
 wire \as1802.regs[12][10] ;
 wire \as1802.regs[12][11] ;
 wire \as1802.regs[12][12] ;
 wire \as1802.regs[12][13] ;
 wire \as1802.regs[12][14] ;
 wire \as1802.regs[12][15] ;
 wire \as1802.regs[12][1] ;
 wire \as1802.regs[12][2] ;
 wire \as1802.regs[12][3] ;
 wire \as1802.regs[12][4] ;
 wire \as1802.regs[12][5] ;
 wire \as1802.regs[12][6] ;
 wire \as1802.regs[12][7] ;
 wire \as1802.regs[12][8] ;
 wire \as1802.regs[12][9] ;
 wire \as1802.regs[13][0] ;
 wire \as1802.regs[13][10] ;
 wire \as1802.regs[13][11] ;
 wire \as1802.regs[13][12] ;
 wire \as1802.regs[13][13] ;
 wire \as1802.regs[13][14] ;
 wire \as1802.regs[13][15] ;
 wire \as1802.regs[13][1] ;
 wire \as1802.regs[13][2] ;
 wire \as1802.regs[13][3] ;
 wire \as1802.regs[13][4] ;
 wire \as1802.regs[13][5] ;
 wire \as1802.regs[13][6] ;
 wire \as1802.regs[13][7] ;
 wire \as1802.regs[13][8] ;
 wire \as1802.regs[13][9] ;
 wire \as1802.regs[14][0] ;
 wire \as1802.regs[14][10] ;
 wire \as1802.regs[14][11] ;
 wire \as1802.regs[14][12] ;
 wire \as1802.regs[14][13] ;
 wire \as1802.regs[14][14] ;
 wire \as1802.regs[14][15] ;
 wire \as1802.regs[14][1] ;
 wire \as1802.regs[14][2] ;
 wire \as1802.regs[14][3] ;
 wire \as1802.regs[14][4] ;
 wire \as1802.regs[14][5] ;
 wire \as1802.regs[14][6] ;
 wire \as1802.regs[14][7] ;
 wire \as1802.regs[14][8] ;
 wire \as1802.regs[14][9] ;
 wire \as1802.regs[15][0] ;
 wire \as1802.regs[15][10] ;
 wire \as1802.regs[15][11] ;
 wire \as1802.regs[15][12] ;
 wire \as1802.regs[15][13] ;
 wire \as1802.regs[15][14] ;
 wire \as1802.regs[15][15] ;
 wire \as1802.regs[15][1] ;
 wire \as1802.regs[15][2] ;
 wire \as1802.regs[15][3] ;
 wire \as1802.regs[15][4] ;
 wire \as1802.regs[15][5] ;
 wire \as1802.regs[15][6] ;
 wire \as1802.regs[15][7] ;
 wire \as1802.regs[15][8] ;
 wire \as1802.regs[15][9] ;
 wire \as1802.regs[1][0] ;
 wire \as1802.regs[1][10] ;
 wire \as1802.regs[1][11] ;
 wire \as1802.regs[1][12] ;
 wire \as1802.regs[1][13] ;
 wire \as1802.regs[1][14] ;
 wire \as1802.regs[1][15] ;
 wire \as1802.regs[1][1] ;
 wire \as1802.regs[1][2] ;
 wire \as1802.regs[1][3] ;
 wire \as1802.regs[1][4] ;
 wire \as1802.regs[1][5] ;
 wire \as1802.regs[1][6] ;
 wire \as1802.regs[1][7] ;
 wire \as1802.regs[1][8] ;
 wire \as1802.regs[1][9] ;
 wire \as1802.regs[2][0] ;
 wire \as1802.regs[2][10] ;
 wire \as1802.regs[2][11] ;
 wire \as1802.regs[2][12] ;
 wire \as1802.regs[2][13] ;
 wire \as1802.regs[2][14] ;
 wire \as1802.regs[2][15] ;
 wire \as1802.regs[2][1] ;
 wire \as1802.regs[2][2] ;
 wire \as1802.regs[2][3] ;
 wire \as1802.regs[2][4] ;
 wire \as1802.regs[2][5] ;
 wire \as1802.regs[2][6] ;
 wire \as1802.regs[2][7] ;
 wire \as1802.regs[2][8] ;
 wire \as1802.regs[2][9] ;
 wire \as1802.regs[3][0] ;
 wire \as1802.regs[3][10] ;
 wire \as1802.regs[3][11] ;
 wire \as1802.regs[3][12] ;
 wire \as1802.regs[3][13] ;
 wire \as1802.regs[3][14] ;
 wire \as1802.regs[3][15] ;
 wire \as1802.regs[3][1] ;
 wire \as1802.regs[3][2] ;
 wire \as1802.regs[3][3] ;
 wire \as1802.regs[3][4] ;
 wire \as1802.regs[3][5] ;
 wire \as1802.regs[3][6] ;
 wire \as1802.regs[3][7] ;
 wire \as1802.regs[3][8] ;
 wire \as1802.regs[3][9] ;
 wire \as1802.regs[4][0] ;
 wire \as1802.regs[4][10] ;
 wire \as1802.regs[4][11] ;
 wire \as1802.regs[4][12] ;
 wire \as1802.regs[4][13] ;
 wire \as1802.regs[4][14] ;
 wire \as1802.regs[4][15] ;
 wire \as1802.regs[4][1] ;
 wire \as1802.regs[4][2] ;
 wire \as1802.regs[4][3] ;
 wire \as1802.regs[4][4] ;
 wire \as1802.regs[4][5] ;
 wire \as1802.regs[4][6] ;
 wire \as1802.regs[4][7] ;
 wire \as1802.regs[4][8] ;
 wire \as1802.regs[4][9] ;
 wire \as1802.regs[5][0] ;
 wire \as1802.regs[5][10] ;
 wire \as1802.regs[5][11] ;
 wire \as1802.regs[5][12] ;
 wire \as1802.regs[5][13] ;
 wire \as1802.regs[5][14] ;
 wire \as1802.regs[5][15] ;
 wire \as1802.regs[5][1] ;
 wire \as1802.regs[5][2] ;
 wire \as1802.regs[5][3] ;
 wire \as1802.regs[5][4] ;
 wire \as1802.regs[5][5] ;
 wire \as1802.regs[5][6] ;
 wire \as1802.regs[5][7] ;
 wire \as1802.regs[5][8] ;
 wire \as1802.regs[5][9] ;
 wire \as1802.regs[6][0] ;
 wire \as1802.regs[6][10] ;
 wire \as1802.regs[6][11] ;
 wire \as1802.regs[6][12] ;
 wire \as1802.regs[6][13] ;
 wire \as1802.regs[6][14] ;
 wire \as1802.regs[6][15] ;
 wire \as1802.regs[6][1] ;
 wire \as1802.regs[6][2] ;
 wire \as1802.regs[6][3] ;
 wire \as1802.regs[6][4] ;
 wire \as1802.regs[6][5] ;
 wire \as1802.regs[6][6] ;
 wire \as1802.regs[6][7] ;
 wire \as1802.regs[6][8] ;
 wire \as1802.regs[6][9] ;
 wire \as1802.regs[7][0] ;
 wire \as1802.regs[7][10] ;
 wire \as1802.regs[7][11] ;
 wire \as1802.regs[7][12] ;
 wire \as1802.regs[7][13] ;
 wire \as1802.regs[7][14] ;
 wire \as1802.regs[7][15] ;
 wire \as1802.regs[7][1] ;
 wire \as1802.regs[7][2] ;
 wire \as1802.regs[7][3] ;
 wire \as1802.regs[7][4] ;
 wire \as1802.regs[7][5] ;
 wire \as1802.regs[7][6] ;
 wire \as1802.regs[7][7] ;
 wire \as1802.regs[7][8] ;
 wire \as1802.regs[7][9] ;
 wire \as1802.regs[8][0] ;
 wire \as1802.regs[8][10] ;
 wire \as1802.regs[8][11] ;
 wire \as1802.regs[8][12] ;
 wire \as1802.regs[8][13] ;
 wire \as1802.regs[8][14] ;
 wire \as1802.regs[8][15] ;
 wire \as1802.regs[8][1] ;
 wire \as1802.regs[8][2] ;
 wire \as1802.regs[8][3] ;
 wire \as1802.regs[8][4] ;
 wire \as1802.regs[8][5] ;
 wire \as1802.regs[8][6] ;
 wire \as1802.regs[8][7] ;
 wire \as1802.regs[8][8] ;
 wire \as1802.regs[8][9] ;
 wire \as1802.regs[9][0] ;
 wire \as1802.regs[9][10] ;
 wire \as1802.regs[9][11] ;
 wire \as1802.regs[9][12] ;
 wire \as1802.regs[9][13] ;
 wire \as1802.regs[9][14] ;
 wire \as1802.regs[9][15] ;
 wire \as1802.regs[9][1] ;
 wire \as1802.regs[9][2] ;
 wire \as1802.regs[9][3] ;
 wire \as1802.regs[9][4] ;
 wire \as1802.regs[9][5] ;
 wire \as1802.regs[9][6] ;
 wire \as1802.regs[9][7] ;
 wire \as1802.regs[9][8] ;
 wire \as1802.regs[9][9] ;
 wire \as1802.will_interrupt ;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_opt_1_0_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1928_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_1928_));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _2176_ (.A(\as1802.X[3] ),
    .Y(_1909_));
 sky130_fd_sc_hd__inv_2 _2177_ (.A(\as1802.X[2] ),
    .Y(_1910_));
 sky130_fd_sc_hd__clkinv_4 _2178_ (.A(\as1802.DF ),
    .Y(_1911_));
 sky130_fd_sc_hd__inv_2 _2179_ (.A(net272),
    .Y(_1912_));
 sky130_fd_sc_hd__inv_2 _2180_ (.A(net26),
    .Y(_1913_));
 sky130_fd_sc_hd__inv_2 _2181_ (.A(\as1802.last_hi_addr[7] ),
    .Y(_1914_));
 sky130_fd_sc_hd__inv_2 _2182_ (.A(\as1802.addr_buff[15] ),
    .Y(_1915_));
 sky130_fd_sc_hd__inv_2 _2183_ (.A(\as1802.last_hi_addr[5] ),
    .Y(_1916_));
 sky130_fd_sc_hd__inv_2 _2184_ (.A(\as1802.addr_buff[13] ),
    .Y(_1917_));
 sky130_fd_sc_hd__inv_2 _2185_ (.A(\as1802.last_hi_addr[0] ),
    .Y(_1918_));
 sky130_fd_sc_hd__inv_2 _2186_ (.A(\as1802.addr_buff[8] ),
    .Y(_1919_));
 sky130_fd_sc_hd__clkinv_4 _2187_ (.A(\as1802.mem_cycle[2] ),
    .Y(_1920_));
 sky130_fd_sc_hd__inv_2 _2188_ (.A(\as1802.mem_cycle[0] ),
    .Y(_1921_));
 sky130_fd_sc_hd__inv_2 _2189_ (.A(\as1802.lda ),
    .Y(_1922_));
 sky130_fd_sc_hd__inv_2 _2190_ (.A(net224),
    .Y(_1923_));
 sky130_fd_sc_hd__inv_2 _2191_ (.A(net221),
    .Y(_1924_));
 sky130_fd_sc_hd__clkinv_4 _2192_ (.A(net237),
    .Y(_1925_));
 sky130_fd_sc_hd__clkinv_4 _2193_ (.A(net233),
    .Y(_1926_));
 sky130_fd_sc_hd__inv_2 _2194_ (.A(net226),
    .Y(_1927_));
 sky130_fd_sc_hd__inv_2 _2195_ (.A(net280),
    .Y(_1928_));
 sky130_fd_sc_hd__inv_2 _2196_ (.A(\as1802.D[6] ),
    .Y(_1929_));
 sky130_fd_sc_hd__inv_2 _2197_ (.A(\as1802.regs[2][0] ),
    .Y(_1930_));
 sky130_fd_sc_hd__clkinv_4 _2198_ (.A(net243),
    .Y(_1931_));
 sky130_fd_sc_hd__clkinv_4 _2199_ (.A(net239),
    .Y(_1932_));
 sky130_fd_sc_hd__inv_2 _2200_ (.A(net13),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _2201_ (.A(net2),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _2202_ (.A(net3),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _2203_ (.A(net4),
    .Y(_0011_));
 sky130_fd_sc_hd__nor3_1 _2204_ (.A(\as1802.mem_cycle[2] ),
    .B(net238),
    .C(\as1802.mem_cycle[0] ),
    .Y(_1933_));
 sky130_fd_sc_hd__or3_1 _2205_ (.A(\as1802.mem_cycle[2] ),
    .B(net238),
    .C(\as1802.mem_cycle[0] ),
    .X(_1934_));
 sky130_fd_sc_hd__and3_1 _2206_ (.A(net279),
    .B(\as1802.instr_cycle[3] ),
    .C(net192),
    .X(_1935_));
 sky130_fd_sc_hd__nor2_2 _2207_ (.A(net220),
    .B(net222),
    .Y(_1936_));
 sky130_fd_sc_hd__or2_4 _2208_ (.A(net221),
    .B(net222),
    .X(_1937_));
 sky130_fd_sc_hd__nand2_8 _2209_ (.A(net224),
    .B(\as1802.instr_latch[4] ),
    .Y(_1938_));
 sky130_fd_sc_hd__nand2b_4 _2210_ (.A_N(\as1802.instr_latch[4] ),
    .B(net224),
    .Y(_1939_));
 sky130_fd_sc_hd__nand2b_4 _2211_ (.A_N(net224),
    .B(\as1802.instr_latch[4] ),
    .Y(_1940_));
 sky130_fd_sc_hd__or2_4 _2212_ (.A(net224),
    .B(\as1802.instr_latch[4] ),
    .X(_1941_));
 sky130_fd_sc_hd__nor2_2 _2213_ (.A(net220),
    .B(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__nor2_4 _2214_ (.A(_1937_),
    .B(_1941_),
    .Y(_1943_));
 sky130_fd_sc_hd__or4_4 _2215_ (.A(net224),
    .B(\as1802.instr_latch[4] ),
    .C(net220),
    .D(net222),
    .X(_1944_));
 sky130_fd_sc_hd__a211o_4 _2216_ (.A1(net224),
    .A2(\as1802.instr_latch[4] ),
    .B1(net220),
    .C1(net223),
    .X(_1945_));
 sky130_fd_sc_hd__nand2_1 _2217_ (.A(net195),
    .B(_1945_),
    .Y(_1946_));
 sky130_fd_sc_hd__nor2_8 _2218_ (.A(net282),
    .B(net192),
    .Y(_1947_));
 sky130_fd_sc_hd__or4_4 _2219_ (.A(\as1802.mem_cycle[2] ),
    .B(net238),
    .C(\as1802.mem_cycle[0] ),
    .D(net280),
    .X(_1948_));
 sky130_fd_sc_hd__nand2_8 _2220_ (.A(net221),
    .B(net222),
    .Y(_1949_));
 sky130_fd_sc_hd__nor2_8 _2221_ (.A(_1941_),
    .B(_1949_),
    .Y(_1950_));
 sky130_fd_sc_hd__or2_4 _2222_ (.A(_1941_),
    .B(_1949_),
    .X(_1951_));
 sky130_fd_sc_hd__nor2_8 _2223_ (.A(net236),
    .B(net237),
    .Y(_1952_));
 sky130_fd_sc_hd__or2_4 _2224_ (.A(net235),
    .B(net237),
    .X(_1953_));
 sky130_fd_sc_hd__nor2_4 _2225_ (.A(net202),
    .B(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__nand2_4 _2226_ (.A(net232),
    .B(_1952_),
    .Y(_1955_));
 sky130_fd_sc_hd__o2111a_2 _2227_ (.A1(net229),
    .A2(_1955_),
    .B1(_1950_),
    .C1(_1947_),
    .D1(_1945_),
    .X(_1956_));
 sky130_fd_sc_hd__nor2_4 _2228_ (.A(net201),
    .B(_1953_),
    .Y(_1957_));
 sky130_fd_sc_hd__nor2_4 _2229_ (.A(net232),
    .B(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__or2_4 _2230_ (.A(net232),
    .B(_1957_),
    .X(_1959_));
 sky130_fd_sc_hd__a31o_1 _2231_ (.A1(\as1802.instr_cycle[1] ),
    .A2(_1956_),
    .A3(_1958_),
    .B1(_1935_),
    .X(_0007_));
 sky130_fd_sc_hd__a21o_2 _2232_ (.A1(\as1802.IE ),
    .A2(net12),
    .B1(\as1802.idle ),
    .X(_1960_));
 sky130_fd_sc_hd__nor3_4 _2233_ (.A(\as1802.will_interrupt ),
    .B(net203),
    .C(_1960_),
    .Y(_1961_));
 sky130_fd_sc_hd__and2_1 _2234_ (.A(net269),
    .B(net279),
    .X(_1962_));
 sky130_fd_sc_hd__a22o_1 _2235_ (.A1(_1947_),
    .A2(_1961_),
    .B1(_1962_),
    .B2(net192),
    .X(_0006_));
 sky130_fd_sc_hd__and2b_2 _2236_ (.A_N(net237),
    .B(net235),
    .X(_1963_));
 sky130_fd_sc_hd__nand2b_4 _2237_ (.A_N(net237),
    .B(net235),
    .Y(_1964_));
 sky130_fd_sc_hd__a2bb2o_4 _2238_ (.A1_N(net235),
    .A2_N(net229),
    .B1(_1964_),
    .B2(net232),
    .X(_1965_));
 sky130_fd_sc_hd__a21o_2 _2239_ (.A1(_1923_),
    .A2(_1936_),
    .B1(net192),
    .X(_1966_));
 sky130_fd_sc_hd__nand2_2 _2240_ (.A(_1924_),
    .B(net223),
    .Y(_1967_));
 sky130_fd_sc_hd__nor2_1 _2241_ (.A(_1938_),
    .B(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hd__or2_4 _2242_ (.A(_1938_),
    .B(_1967_),
    .X(_1969_));
 sky130_fd_sc_hd__nor2_1 _2243_ (.A(_1966_),
    .B(net173),
    .Y(_1970_));
 sky130_fd_sc_hd__or4_2 _2244_ (.A(net212),
    .B(net213),
    .C(net211),
    .D(\as1802.D[6] ),
    .X(_1971_));
 sky130_fd_sc_hd__or4_2 _2245_ (.A(net217),
    .B(net218),
    .C(net214),
    .D(net215),
    .X(_1972_));
 sky130_fd_sc_hd__and2_4 _2246_ (.A(net235),
    .B(\as1802.instr_latch[0] ),
    .X(_1973_));
 sky130_fd_sc_hd__nand2_2 _2247_ (.A(net235),
    .B(\as1802.instr_latch[0] ),
    .Y(_1974_));
 sky130_fd_sc_hd__nand2_1 _2248_ (.A(\as1802.DF ),
    .B(_1973_),
    .Y(_1975_));
 sky130_fd_sc_hd__nand2b_4 _2249_ (.A_N(net235),
    .B(\as1802.instr_latch[0] ),
    .Y(_1976_));
 sky130_fd_sc_hd__o32a_1 _2250_ (.A1(_1964_),
    .A2(_1971_),
    .A3(_1972_),
    .B1(_1976_),
    .B2(_1913_),
    .X(_1977_));
 sky130_fd_sc_hd__a21oi_1 _2251_ (.A1(_1975_),
    .A2(_1977_),
    .B1(net231),
    .Y(_1978_));
 sky130_fd_sc_hd__nor2_4 _2252_ (.A(net202),
    .B(_1974_),
    .Y(_1979_));
 sky130_fd_sc_hd__nand2_4 _2253_ (.A(net231),
    .B(_1973_),
    .Y(_1980_));
 sky130_fd_sc_hd__nor2_8 _2254_ (.A(net202),
    .B(_1976_),
    .Y(_1981_));
 sky130_fd_sc_hd__a22o_1 _2255_ (.A1(\as1802.EF_l[3] ),
    .A2(_1979_),
    .B1(_1981_),
    .B2(\as1802.EF_l[1] ),
    .X(_1982_));
 sky130_fd_sc_hd__nand2_1 _2256_ (.A(net232),
    .B(_1963_),
    .Y(_1983_));
 sky130_fd_sc_hd__and3_1 _2257_ (.A(net231),
    .B(\as1802.EF_l[2] ),
    .C(_1963_),
    .X(_1984_));
 sky130_fd_sc_hd__o21a_1 _2258_ (.A1(net202),
    .A2(\as1802.EF_l[0] ),
    .B1(_1952_),
    .X(_1985_));
 sky130_fd_sc_hd__nand2_8 _2259_ (.A(net202),
    .B(_1973_),
    .Y(_1986_));
 sky130_fd_sc_hd__inv_2 _2260_ (.A(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__nor2_2 _2261_ (.A(net231),
    .B(_1953_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_4 _2262_ (.A(_1926_),
    .B(_1952_),
    .Y(_1989_));
 sky130_fd_sc_hd__or4_4 _2263_ (.A(_1978_),
    .B(_1982_),
    .C(_1984_),
    .D(_1985_),
    .X(_1990_));
 sky130_fd_sc_hd__xnor2_4 _2264_ (.A(net201),
    .B(_1990_),
    .Y(_1991_));
 sky130_fd_sc_hd__inv_2 _2265_ (.A(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__nor2_4 _2266_ (.A(_1937_),
    .B(_1938_),
    .Y(_1993_));
 sky130_fd_sc_hd__or2_2 _2267_ (.A(_1937_),
    .B(_1938_),
    .X(_1994_));
 sky130_fd_sc_hd__and3_1 _2268_ (.A(net195),
    .B(_1991_),
    .C(_1993_),
    .X(_1995_));
 sky130_fd_sc_hd__a21o_1 _2269_ (.A1(_1965_),
    .A2(_1970_),
    .B1(_1995_),
    .X(_1996_));
 sky130_fd_sc_hd__and2_1 _2270_ (.A(net269),
    .B(_1983_),
    .X(_1997_));
 sky130_fd_sc_hd__or2_1 _2271_ (.A(_1938_),
    .B(_1949_),
    .X(_1998_));
 sky130_fd_sc_hd__and3b_2 _2272_ (.A_N(_1998_),
    .B(_1989_),
    .C(_1997_),
    .X(_1999_));
 sky130_fd_sc_hd__inv_2 _2273_ (.A(_1999_),
    .Y(_2000_));
 sky130_fd_sc_hd__and3_1 _2274_ (.A(net279),
    .B(\as1802.instr_cycle[1] ),
    .C(net192),
    .X(_2001_));
 sky130_fd_sc_hd__a31o_1 _2275_ (.A1(_1945_),
    .A2(_1947_),
    .A3(_1999_),
    .B1(_2001_),
    .X(_2002_));
 sky130_fd_sc_hd__nor2_2 _2276_ (.A(net232),
    .B(net229),
    .Y(_2003_));
 sky130_fd_sc_hd__or2_4 _2277_ (.A(net231),
    .B(net229),
    .X(_2004_));
 sky130_fd_sc_hd__nand2_8 _2278_ (.A(net231),
    .B(net229),
    .Y(_2005_));
 sky130_fd_sc_hd__a22o_2 _2279_ (.A1(_1975_),
    .A2(_1977_),
    .B1(_2004_),
    .B2(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__o21a_1 _2280_ (.A1(_1971_),
    .A2(_1972_),
    .B1(_1963_),
    .X(_2007_));
 sky130_fd_sc_hd__a2bb2o_1 _2281_ (.A1_N(_1976_),
    .A2_N(net26),
    .B1(_1911_),
    .B2(_1973_),
    .X(_2008_));
 sky130_fd_sc_hd__o211ai_4 _2282_ (.A1(_2007_),
    .A2(_2008_),
    .B1(_2004_),
    .C1(_2005_),
    .Y(_2009_));
 sky130_fd_sc_hd__a21oi_2 _2283_ (.A1(\as1802.IE ),
    .A2(_1957_),
    .B1(_1988_),
    .Y(_2010_));
 sky130_fd_sc_hd__and3_4 _2284_ (.A(_2006_),
    .B(_2009_),
    .C(_2010_),
    .X(_2011_));
 sky130_fd_sc_hd__nand2_2 _2285_ (.A(net268),
    .B(_1958_),
    .Y(_2012_));
 sky130_fd_sc_hd__and4b_1 _2286_ (.A_N(_2011_),
    .B(_1958_),
    .C(_1956_),
    .D(net269),
    .X(_2013_));
 sky130_fd_sc_hd__a211o_1 _2287_ (.A1(_1962_),
    .A2(_1996_),
    .B1(_2002_),
    .C1(_2013_),
    .X(_0005_));
 sky130_fd_sc_hd__nor2_1 _2288_ (.A(net269),
    .B(\as1802.instr_cycle[1] ),
    .Y(_2014_));
 sky130_fd_sc_hd__o311a_1 _2289_ (.A1(\as1802.instr_cycle[1] ),
    .A2(\as1802.instr_cycle[3] ),
    .A3(_1992_),
    .B1(_1993_),
    .C1(net195),
    .X(_2015_));
 sky130_fd_sc_hd__nand2_2 _2290_ (.A(net223),
    .B(_1942_),
    .Y(_2016_));
 sky130_fd_sc_hd__or3b_1 _2291_ (.A(net193),
    .B(_1936_),
    .C_N(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__nand2b_4 _2292_ (.A_N(net222),
    .B(net221),
    .Y(_2018_));
 sky130_fd_sc_hd__or3_1 _2293_ (.A(_1938_),
    .B(_2017_),
    .C(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__and2_4 _2294_ (.A(net268),
    .B(_1965_),
    .X(_2020_));
 sky130_fd_sc_hd__nand2_8 _2295_ (.A(net268),
    .B(_1965_),
    .Y(_2021_));
 sky130_fd_sc_hd__nand2_8 _2296_ (.A(net176),
    .B(_2021_),
    .Y(_2022_));
 sky130_fd_sc_hd__or2_4 _2297_ (.A(_1939_),
    .B(_1967_),
    .X(_2023_));
 sky130_fd_sc_hd__and2_2 _2298_ (.A(_2022_),
    .B(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__or2_2 _2299_ (.A(_1989_),
    .B(_1998_),
    .X(_2025_));
 sky130_fd_sc_hd__or3_4 _2300_ (.A(_1988_),
    .B(_1997_),
    .C(_1998_),
    .X(_2026_));
 sky130_fd_sc_hd__a21o_1 _2301_ (.A1(_1939_),
    .A2(_1940_),
    .B1(_1924_),
    .X(_2027_));
 sky130_fd_sc_hd__or2_1 _2302_ (.A(_1941_),
    .B(_2018_),
    .X(_2028_));
 sky130_fd_sc_hd__nor2_2 _2303_ (.A(\as1802.instr_latch[5] ),
    .B(_1967_),
    .Y(_2029_));
 sky130_fd_sc_hd__nand2_1 _2304_ (.A(\as1802.instr_cycle[3] ),
    .B(_1950_),
    .Y(_2030_));
 sky130_fd_sc_hd__o311a_1 _2305_ (.A1(net190),
    .A2(_1958_),
    .A3(_2014_),
    .B1(_2027_),
    .C1(_1945_),
    .X(_2031_));
 sky130_fd_sc_hd__and4_1 _2306_ (.A(_2024_),
    .B(_2025_),
    .C(_2026_),
    .D(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__and4b_1 _2307_ (.A_N(_2029_),
    .B(_2032_),
    .C(_2030_),
    .D(net187),
    .X(_2033_));
 sky130_fd_sc_hd__o21ai_1 _2308_ (.A1(net192),
    .A2(_2033_),
    .B1(_2019_),
    .Y(_2034_));
 sky130_fd_sc_hd__nor2_4 _2309_ (.A(_1940_),
    .B(_2018_),
    .Y(_2035_));
 sky130_fd_sc_hd__or4bb_4 _2310_ (.A(net224),
    .B(net222),
    .C_N(net221),
    .D_N(\as1802.instr_latch[4] ),
    .X(_2036_));
 sky130_fd_sc_hd__o32a_1 _2311_ (.A1(net268),
    .A2(\as1802.instr_cycle[1] ),
    .A3(\as1802.instr_cycle[3] ),
    .B1(_2015_),
    .B2(_2034_),
    .X(_2037_));
 sky130_fd_sc_hd__or2_1 _2312_ (.A(\as1802.will_interrupt ),
    .B(net193),
    .X(_2038_));
 sky130_fd_sc_hd__o21a_1 _2313_ (.A1(_1960_),
    .A2(_2038_),
    .B1(net272),
    .X(_2039_));
 sky130_fd_sc_hd__a41o_1 _2314_ (.A1(net269),
    .A2(_1956_),
    .A3(_1958_),
    .A4(_2011_),
    .B1(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__a21o_1 _2315_ (.A1(net231),
    .A2(_1953_),
    .B1(_1957_),
    .X(_2041_));
 sky130_fd_sc_hd__or3_1 _2316_ (.A(net280),
    .B(_2037_),
    .C(_2040_),
    .X(_0004_));
 sky130_fd_sc_hd__a31oi_4 _2317_ (.A1(_2006_),
    .A2(_2009_),
    .A3(_2010_),
    .B1(_2041_),
    .Y(_2042_));
 sky130_fd_sc_hd__nand2_4 _2318_ (.A(net203),
    .B(_1950_),
    .Y(_2043_));
 sky130_fd_sc_hd__nand2_4 _2319_ (.A(net203),
    .B(net195),
    .Y(_2044_));
 sky130_fd_sc_hd__nor2_4 _2320_ (.A(net270),
    .B(_1948_),
    .Y(_2045_));
 sky130_fd_sc_hd__or2_4 _2321_ (.A(net270),
    .B(_1948_),
    .X(_2046_));
 sky130_fd_sc_hd__nand2_2 _2322_ (.A(_1950_),
    .B(_2045_),
    .Y(_2047_));
 sky130_fd_sc_hd__a211oi_4 _2323_ (.A1(_2011_),
    .A2(_2012_),
    .B1(_2042_),
    .C1(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__a211o_4 _2324_ (.A1(_2011_),
    .A2(_2012_),
    .B1(_2042_),
    .C1(_2047_),
    .X(_2049_));
 sky130_fd_sc_hd__or2_4 _2325_ (.A(net271),
    .B(_2025_),
    .X(_2050_));
 sky130_fd_sc_hd__or3b_1 _2326_ (.A(_1994_),
    .B(net271),
    .C_N(net268),
    .X(_2051_));
 sky130_fd_sc_hd__nand3b_1 _2327_ (.A_N(_1961_),
    .B(_2050_),
    .C(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hd__nor2_2 _2328_ (.A(net274),
    .B(net173),
    .Y(_2053_));
 sky130_fd_sc_hd__nand2_2 _2329_ (.A(net176),
    .B(_2045_),
    .Y(_2054_));
 sky130_fd_sc_hd__nor2_2 _2330_ (.A(_2021_),
    .B(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__or2_4 _2331_ (.A(_2021_),
    .B(_2054_),
    .X(_2056_));
 sky130_fd_sc_hd__and3_2 _2332_ (.A(net229),
    .B(_1999_),
    .C(_2045_),
    .X(_2057_));
 sky130_fd_sc_hd__or3_4 _2333_ (.A(net201),
    .B(_2000_),
    .C(net184),
    .X(_2058_));
 sky130_fd_sc_hd__a211o_1 _2334_ (.A1(_1947_),
    .A2(_2052_),
    .B1(net133),
    .C1(_2057_),
    .X(_2059_));
 sky130_fd_sc_hd__and4_2 _2335_ (.A(net268),
    .B(_1950_),
    .C(_2042_),
    .D(_2045_),
    .X(_2060_));
 sky130_fd_sc_hd__inv_2 _2336_ (.A(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__or3_2 _2337_ (.A(net134),
    .B(_2059_),
    .C(_2060_),
    .X(_2062_));
 sky130_fd_sc_hd__or2_1 _2338_ (.A(net268),
    .B(_1994_),
    .X(_2063_));
 sky130_fd_sc_hd__or2_4 _2339_ (.A(net273),
    .B(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__nor2_4 _2340_ (.A(_1948_),
    .B(_2064_),
    .Y(_2065_));
 sky130_fd_sc_hd__or2_4 _2341_ (.A(_1948_),
    .B(_2064_),
    .X(_2066_));
 sky130_fd_sc_hd__or3_4 _2342_ (.A(net268),
    .B(_1959_),
    .C(_2043_),
    .X(_2067_));
 sky130_fd_sc_hd__nor2_4 _2343_ (.A(\as1802.instr_cycle[1] ),
    .B(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__and2_4 _2344_ (.A(_1947_),
    .B(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__nand2_4 _2345_ (.A(_1947_),
    .B(_2068_),
    .Y(_2070_));
 sky130_fd_sc_hd__or3_1 _2346_ (.A(net269),
    .B(_1959_),
    .C(_2043_),
    .X(_2071_));
 sky130_fd_sc_hd__or3_4 _2347_ (.A(\as1802.instr_cycle[1] ),
    .B(_1948_),
    .C(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__or3_2 _2348_ (.A(_2062_),
    .B(_2065_),
    .C(_2069_),
    .X(_2073_));
 sky130_fd_sc_hd__nand2_4 _2349_ (.A(\as1802.instr_cycle[1] ),
    .B(_1947_),
    .Y(_2074_));
 sky130_fd_sc_hd__nor2_4 _2350_ (.A(_2067_),
    .B(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__nor4_4 _2351_ (.A(net268),
    .B(_1959_),
    .C(_2043_),
    .D(_2074_),
    .Y(_2076_));
 sky130_fd_sc_hd__or2_4 _2352_ (.A(_2071_),
    .B(_2074_),
    .X(_2077_));
 sky130_fd_sc_hd__or2_2 _2353_ (.A(_2073_),
    .B(_2075_),
    .X(_2078_));
 sky130_fd_sc_hd__or2_4 _2354_ (.A(net271),
    .B(_2019_),
    .X(_2079_));
 sky130_fd_sc_hd__nor2_8 _2355_ (.A(net282),
    .B(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__or2_4 _2356_ (.A(net282),
    .B(_2079_),
    .X(_2081_));
 sky130_fd_sc_hd__a21oi_2 _2357_ (.A1(_1939_),
    .A2(_1940_),
    .B1(net220),
    .Y(_2082_));
 sky130_fd_sc_hd__or3b_4 _2358_ (.A(net222),
    .B(net184),
    .C_N(_2082_),
    .X(_2083_));
 sky130_fd_sc_hd__o21ai_2 _2359_ (.A1(_2016_),
    .A2(net184),
    .B1(_2083_),
    .Y(_2084_));
 sky130_fd_sc_hd__or4_4 _2360_ (.A(_1924_),
    .B(net222),
    .C(_1939_),
    .D(net184),
    .X(_2085_));
 sky130_fd_sc_hd__nor3_4 _2361_ (.A(_1939_),
    .B(_2018_),
    .C(net184),
    .Y(_2086_));
 sky130_fd_sc_hd__or3_4 _2362_ (.A(_1939_),
    .B(_2018_),
    .C(net184),
    .X(_2087_));
 sky130_fd_sc_hd__or2_2 _2363_ (.A(_2084_),
    .B(_2086_),
    .X(_2088_));
 sky130_fd_sc_hd__nor2_2 _2364_ (.A(_2080_),
    .B(_2088_),
    .Y(_2089_));
 sky130_fd_sc_hd__or2_2 _2365_ (.A(_2080_),
    .B(_2088_),
    .X(_2090_));
 sky130_fd_sc_hd__or3_4 _2366_ (.A(net236),
    .B(net231),
    .C(net201),
    .X(_2091_));
 sky130_fd_sc_hd__nor2_8 _2367_ (.A(_1925_),
    .B(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__or2_1 _2368_ (.A(_1925_),
    .B(_2091_),
    .X(_2093_));
 sky130_fd_sc_hd__nor2_2 _2369_ (.A(_2054_),
    .B(net167),
    .Y(_2094_));
 sky130_fd_sc_hd__or2_2 _2370_ (.A(_2054_),
    .B(net167),
    .X(_2095_));
 sky130_fd_sc_hd__and4_4 _2371_ (.A(net201),
    .B(net176),
    .C(_1987_),
    .D(_2045_),
    .X(_2096_));
 sky130_fd_sc_hd__or3_4 _2372_ (.A(net230),
    .B(_1986_),
    .C(_2054_),
    .X(_2097_));
 sky130_fd_sc_hd__nor4_2 _2373_ (.A(net235),
    .B(net237),
    .C(net232),
    .D(net229),
    .Y(_2098_));
 sky130_fd_sc_hd__nand2_4 _2374_ (.A(_1952_),
    .B(_2003_),
    .Y(_2099_));
 sky130_fd_sc_hd__a211o_1 _2375_ (.A1(_1964_),
    .A2(_1976_),
    .B1(_2004_),
    .C1(_2022_),
    .X(_2100_));
 sky130_fd_sc_hd__a211o_4 _2376_ (.A1(_2099_),
    .A2(_2100_),
    .B1(_2024_),
    .C1(net184),
    .X(_2101_));
 sky130_fd_sc_hd__inv_2 _2377_ (.A(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__o21a_1 _2378_ (.A1(_1976_),
    .A2(_2020_),
    .B1(_1964_),
    .X(_2103_));
 sky130_fd_sc_hd__o32a_4 _2379_ (.A1(net173),
    .A2(_2004_),
    .A3(_2103_),
    .B1(_2099_),
    .B2(_2024_),
    .X(_2104_));
 sky130_fd_sc_hd__nor2_8 _2380_ (.A(_2046_),
    .B(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__nor2_1 _2381_ (.A(_2096_),
    .B(_2105_),
    .Y(_2106_));
 sky130_fd_sc_hd__or2_4 _2382_ (.A(_2096_),
    .B(_2105_),
    .X(_2107_));
 sky130_fd_sc_hd__a221o_4 _2383_ (.A1(net236),
    .A2(net83),
    .B1(_2107_),
    .B2(\as1802.X[1] ),
    .C1(net131),
    .X(_2108_));
 sky130_fd_sc_hd__and4_4 _2384_ (.A(net176),
    .B(_1973_),
    .C(_2003_),
    .D(_2045_),
    .X(_2109_));
 sky130_fd_sc_hd__nor2_8 _2385_ (.A(_2105_),
    .B(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__a21oi_4 _2386_ (.A1(\as1802.P[1] ),
    .A2(net81),
    .B1(_2108_),
    .Y(_2111_));
 sky130_fd_sc_hd__a21o_4 _2387_ (.A1(\as1802.P[1] ),
    .A2(net81),
    .B1(_2108_),
    .X(_2112_));
 sky130_fd_sc_hd__a221o_4 _2388_ (.A1(\as1802.P[0] ),
    .A2(net81),
    .B1(net84),
    .B2(net237),
    .C1(_2107_),
    .X(_2113_));
 sky130_fd_sc_hd__nand2_1 _2389_ (.A(net128),
    .B(_2106_),
    .Y(_2114_));
 sky130_fd_sc_hd__o21a_4 _2390_ (.A1(\as1802.X[0] ),
    .A2(_2110_),
    .B1(_2113_),
    .X(_2115_));
 sky130_fd_sc_hd__o21ai_4 _2391_ (.A1(\as1802.X[0] ),
    .A2(_2110_),
    .B1(_2113_),
    .Y(_2116_));
 sky130_fd_sc_hd__nor2_8 _2392_ (.A(_2111_),
    .B(_2116_),
    .Y(_2117_));
 sky130_fd_sc_hd__a221o_2 _2393_ (.A1(\as1802.P[3] ),
    .A2(net81),
    .B1(net83),
    .B2(net225),
    .C1(_2107_),
    .X(_2118_));
 sky130_fd_sc_hd__o21a_2 _2394_ (.A1(\as1802.X[3] ),
    .A2(_2110_),
    .B1(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__o21ai_4 _2395_ (.A1(\as1802.X[3] ),
    .A2(_2110_),
    .B1(_2118_),
    .Y(_2120_));
 sky130_fd_sc_hd__a221o_4 _2396_ (.A1(\as1802.P[2] ),
    .A2(net81),
    .B1(net84),
    .B2(net234),
    .C1(_2107_),
    .X(_2121_));
 sky130_fd_sc_hd__o21a_2 _2397_ (.A1(\as1802.X[2] ),
    .A2(_2110_),
    .B1(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__o21ai_4 _2398_ (.A1(\as1802.X[2] ),
    .A2(_2110_),
    .B1(_2121_),
    .Y(_2123_));
 sky130_fd_sc_hd__nor2_4 _2399_ (.A(_2120_),
    .B(_2123_),
    .Y(_2124_));
 sky130_fd_sc_hd__or4_4 _2400_ (.A(net282),
    .B(_2073_),
    .C(_2088_),
    .D(_2114_),
    .X(_2125_));
 sky130_fd_sc_hd__and3_4 _2401_ (.A(_2117_),
    .B(_2124_),
    .C(net72),
    .X(_2126_));
 sky130_fd_sc_hd__mux4_1 _2402_ (.A0(\as1802.regs[8][0] ),
    .A1(\as1802.regs[9][0] ),
    .A2(\as1802.regs[10][0] ),
    .A3(\as1802.regs[11][0] ),
    .S0(net256),
    .S1(net246),
    .X(_2127_));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(\as1802.regs[14][0] ),
    .A1(\as1802.regs[15][0] ),
    .S(net257),
    .X(_2128_));
 sky130_fd_sc_hd__nand2_1 _2404_ (.A(net245),
    .B(_2128_),
    .Y(_2129_));
 sky130_fd_sc_hd__mux2_1 _2405_ (.A0(\as1802.regs[12][0] ),
    .A1(\as1802.regs[13][0] ),
    .S(net257),
    .X(_2130_));
 sky130_fd_sc_hd__nand2b_1 _2406_ (.A_N(net245),
    .B(_2130_),
    .Y(_2131_));
 sky130_fd_sc_hd__o21ai_1 _2407_ (.A1(net242),
    .A2(_2127_),
    .B1(net239),
    .Y(_2132_));
 sky130_fd_sc_hd__a31o_4 _2408_ (.A1(net242),
    .A2(_2129_),
    .A3(_2131_),
    .B1(_2132_),
    .X(_2133_));
 sky130_fd_sc_hd__mux4_1 _2409_ (.A0(\as1802.regs[4][0] ),
    .A1(\as1802.regs[5][0] ),
    .A2(\as1802.regs[6][0] ),
    .A3(\as1802.regs[7][0] ),
    .S0(net260),
    .S1(net249),
    .X(_2134_));
 sky130_fd_sc_hd__mux4_1 _2410_ (.A0(\as1802.regs[0][0] ),
    .A1(\as1802.regs[1][0] ),
    .A2(\as1802.regs[2][0] ),
    .A3(\as1802.regs[3][0] ),
    .S0(net260),
    .S1(net249),
    .X(_2135_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(_2134_),
    .A1(_2135_),
    .S(net198),
    .X(_2136_));
 sky130_fd_sc_hd__nand2_2 _2412_ (.A(net197),
    .B(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__and2_4 _2413_ (.A(_2133_),
    .B(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__nand2_4 _2414_ (.A(_2133_),
    .B(_2137_),
    .Y(_2139_));
 sky130_fd_sc_hd__nor2_4 _2415_ (.A(net200),
    .B(net156),
    .Y(_2140_));
 sky130_fd_sc_hd__nand2_4 _2416_ (.A(net228),
    .B(net155),
    .Y(_2141_));
 sky130_fd_sc_hd__nor2_1 _2417_ (.A(net228),
    .B(net155),
    .Y(_2142_));
 sky130_fd_sc_hd__nor2_1 _2418_ (.A(_2140_),
    .B(_2142_),
    .Y(_2143_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(net209),
    .A1(net156),
    .S(_2066_),
    .X(_2144_));
 sky130_fd_sc_hd__mux2_1 _2420_ (.A0(_2143_),
    .A1(_2144_),
    .S(_2056_),
    .X(_2145_));
 sky130_fd_sc_hd__xnor2_1 _2421_ (.A(net134),
    .B(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__nor2_1 _2422_ (.A(_2069_),
    .B(_2146_),
    .Y(_2147_));
 sky130_fd_sc_hd__nor2_8 _2423_ (.A(_1948_),
    .B(_2050_),
    .Y(_2148_));
 sky130_fd_sc_hd__or2_2 _2424_ (.A(_1948_),
    .B(_2050_),
    .X(_2149_));
 sky130_fd_sc_hd__nor2_2 _2425_ (.A(_2025_),
    .B(net184),
    .Y(_2150_));
 sky130_fd_sc_hd__a211o_1 _2426_ (.A1(net16),
    .A2(_2069_),
    .B1(_2147_),
    .C1(_2148_),
    .X(_2151_));
 sky130_fd_sc_hd__o211a_1 _2427_ (.A1(_2143_),
    .A2(net126),
    .B1(_2151_),
    .C1(net81),
    .X(_2152_));
 sky130_fd_sc_hd__or4b_2 _2428_ (.A(net270),
    .B(net192),
    .C(net191),
    .D_N(_1945_),
    .X(_2153_));
 sky130_fd_sc_hd__o31a_1 _2429_ (.A1(net270),
    .A2(_1966_),
    .A3(net187),
    .B1(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__or4b_1 _2430_ (.A(net270),
    .B(\as1802.instr_latch[5] ),
    .C(net220),
    .D_N(net223),
    .X(_2155_));
 sky130_fd_sc_hd__nor2_4 _2431_ (.A(net274),
    .B(_1944_),
    .Y(_2156_));
 sky130_fd_sc_hd__or2_2 _2432_ (.A(net270),
    .B(_1944_),
    .X(_2157_));
 sky130_fd_sc_hd__o31a_1 _2433_ (.A1(net270),
    .A2(_1944_),
    .A3(_2098_),
    .B1(_2155_),
    .X(_2158_));
 sky130_fd_sc_hd__o311a_4 _2434_ (.A1(net270),
    .A2(_1966_),
    .A3(net187),
    .B1(_2153_),
    .C1(_2158_),
    .X(_2159_));
 sky130_fd_sc_hd__nand2_8 _2435_ (.A(_2083_),
    .B(_2159_),
    .Y(_2160_));
 sky130_fd_sc_hd__and3_1 _2436_ (.A(\as1802.X[1] ),
    .B(_2083_),
    .C(_2159_),
    .X(_2161_));
 sky130_fd_sc_hd__a21o_1 _2437_ (.A1(net236),
    .A2(_2160_),
    .B1(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__a21oi_2 _2438_ (.A1(net236),
    .A2(_2160_),
    .B1(_2161_),
    .Y(_2163_));
 sky130_fd_sc_hd__a21o_1 _2439_ (.A1(_2083_),
    .A2(_2159_),
    .B1(\as1802.instr_latch[0] ),
    .X(_2164_));
 sky130_fd_sc_hd__nand3b_2 _2440_ (.A_N(\as1802.X[0] ),
    .B(_2083_),
    .C(_2159_),
    .Y(_2165_));
 sky130_fd_sc_hd__nand2_1 _2441_ (.A(net147),
    .B(net139),
    .Y(_2166_));
 sky130_fd_sc_hd__and3_1 _2442_ (.A(\as1802.regs[15][0] ),
    .B(net147),
    .C(net139),
    .X(_2167_));
 sky130_fd_sc_hd__mux2_8 _2443_ (.A0(_1910_),
    .A1(net202),
    .S(_2160_),
    .X(_2168_));
 sky130_fd_sc_hd__mux2_2 _2444_ (.A0(\as1802.X[2] ),
    .A1(net234),
    .S(_2160_),
    .X(_2169_));
 sky130_fd_sc_hd__and3_1 _2445_ (.A(\as1802.regs[13][0] ),
    .B(net147),
    .C(net139),
    .X(_2170_));
 sky130_fd_sc_hd__a211o_1 _2446_ (.A1(\as1802.regs[12][0] ),
    .A2(net97),
    .B1(_2170_),
    .C1(net120),
    .X(_2171_));
 sky130_fd_sc_hd__a211o_1 _2447_ (.A1(\as1802.regs[14][0] ),
    .A2(net97),
    .B1(_2167_),
    .C1(net112),
    .X(_2172_));
 sky130_fd_sc_hd__a21oi_2 _2448_ (.A1(_2171_),
    .A2(_2172_),
    .B1(net93),
    .Y(_2173_));
 sky130_fd_sc_hd__a21o_1 _2449_ (.A1(net148),
    .A2(net140),
    .B1(\as1802.regs[8][0] ),
    .X(_2174_));
 sky130_fd_sc_hd__o211a_1 _2450_ (.A1(\as1802.regs[9][0] ),
    .A2(net96),
    .B1(_2174_),
    .C1(net113),
    .X(_2175_));
 sky130_fd_sc_hd__a21o_1 _2451_ (.A1(net147),
    .A2(net139),
    .B1(\as1802.regs[10][0] ),
    .X(_0359_));
 sky130_fd_sc_hd__o211a_1 _2452_ (.A1(\as1802.regs[11][0] ),
    .A2(net96),
    .B1(_0359_),
    .C1(net120),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_8 _2453_ (.A0(_1909_),
    .A1(net200),
    .S(_2160_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_2 _2454_ (.A0(\as1802.X[3] ),
    .A1(net226),
    .S(_2160_),
    .X(_0362_));
 sky130_fd_sc_hd__o31ai_4 _2455_ (.A1(net89),
    .A2(_2175_),
    .A3(_0360_),
    .B1(net85),
    .Y(_0363_));
 sky130_fd_sc_hd__and3_1 _2456_ (.A(\as1802.regs[3][0] ),
    .B(net151),
    .C(net143),
    .X(_0364_));
 sky130_fd_sc_hd__and3_1 _2457_ (.A(\as1802.regs[1][0] ),
    .B(net151),
    .C(net143),
    .X(_0365_));
 sky130_fd_sc_hd__a211o_1 _2458_ (.A1(\as1802.regs[0][0] ),
    .A2(net101),
    .B1(_0365_),
    .C1(net121),
    .X(_0366_));
 sky130_fd_sc_hd__a211o_1 _2459_ (.A1(\as1802.regs[2][0] ),
    .A2(net104),
    .B1(_0364_),
    .C1(net114),
    .X(_0367_));
 sky130_fd_sc_hd__a21oi_1 _2460_ (.A1(_0366_),
    .A2(_0367_),
    .B1(net90),
    .Y(_0368_));
 sky130_fd_sc_hd__and3_1 _2461_ (.A(\as1802.regs[7][0] ),
    .B(net150),
    .C(net142),
    .X(_0369_));
 sky130_fd_sc_hd__and3_1 _2462_ (.A(\as1802.regs[5][0] ),
    .B(net150),
    .C(net142),
    .X(_0370_));
 sky130_fd_sc_hd__a211o_1 _2463_ (.A1(\as1802.regs[4][0] ),
    .A2(net101),
    .B1(_0370_),
    .C1(net121),
    .X(_0371_));
 sky130_fd_sc_hd__a211o_1 _2464_ (.A1(\as1802.regs[6][0] ),
    .A2(net101),
    .B1(_0369_),
    .C1(net114),
    .X(_0372_));
 sky130_fd_sc_hd__a21oi_1 _2465_ (.A1(_0371_),
    .A2(_0372_),
    .B1(net94),
    .Y(_0373_));
 sky130_fd_sc_hd__o32a_4 _2466_ (.A1(net85),
    .A2(_0368_),
    .A3(_0373_),
    .B1(_0363_),
    .B2(_2173_),
    .X(_0374_));
 sky130_fd_sc_hd__o21a_1 _2467_ (.A1(net219),
    .A2(_2085_),
    .B1(net84),
    .X(_0375_));
 sky130_fd_sc_hd__o32a_1 _2468_ (.A1(_2096_),
    .A2(_2102_),
    .A3(_0375_),
    .B1(_0374_),
    .B2(_2086_),
    .X(_0376_));
 sky130_fd_sc_hd__a211o_2 _2469_ (.A1(_1930_),
    .A2(net131),
    .B1(_2152_),
    .C1(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _2470_ (.A0(\as1802.regs[15][0] ),
    .A1(net68),
    .S(_2126_),
    .X(_0012_));
 sky130_fd_sc_hd__or2_4 _2471_ (.A(net220),
    .B(_1939_),
    .X(_0378_));
 sky130_fd_sc_hd__nor3_4 _2472_ (.A(_1937_),
    .B(_1939_),
    .C(net184),
    .Y(_0379_));
 sky130_fd_sc_hd__or3_4 _2473_ (.A(_1937_),
    .B(_1939_),
    .C(net184),
    .X(_0380_));
 sky130_fd_sc_hd__and3_1 _2474_ (.A(\as1802.regs[11][1] ),
    .B(net147),
    .C(net139),
    .X(_0381_));
 sky130_fd_sc_hd__a211o_1 _2475_ (.A1(\as1802.regs[10][1] ),
    .A2(net96),
    .B1(_0381_),
    .C1(net112),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _2476_ (.A0(\as1802.regs[9][1] ),
    .A1(\as1802.regs[8][1] ),
    .S(net96),
    .X(_0383_));
 sky130_fd_sc_hd__o211a_2 _2477_ (.A1(net120),
    .A2(_0383_),
    .B1(_0382_),
    .C1(net93),
    .X(_0384_));
 sky130_fd_sc_hd__and3_1 _2478_ (.A(\as1802.regs[15][1] ),
    .B(net148),
    .C(net140),
    .X(_0385_));
 sky130_fd_sc_hd__a211o_1 _2479_ (.A1(\as1802.regs[14][1] ),
    .A2(net96),
    .B1(_0385_),
    .C1(net113),
    .X(_0386_));
 sky130_fd_sc_hd__and3_1 _2480_ (.A(\as1802.regs[13][1] ),
    .B(net148),
    .C(net140),
    .X(_0387_));
 sky130_fd_sc_hd__a211o_1 _2481_ (.A1(\as1802.regs[12][1] ),
    .A2(net97),
    .B1(_0387_),
    .C1(net120),
    .X(_0388_));
 sky130_fd_sc_hd__a31o_2 _2482_ (.A1(net89),
    .A2(_0386_),
    .A3(_0388_),
    .B1(net87),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _2483_ (.A0(\as1802.regs[1][1] ),
    .A1(\as1802.regs[0][1] ),
    .S(net102),
    .X(_0390_));
 sky130_fd_sc_hd__and3_1 _2484_ (.A(\as1802.regs[3][1] ),
    .B(net150),
    .C(net142),
    .X(_0391_));
 sky130_fd_sc_hd__a211o_1 _2485_ (.A1(\as1802.regs[2][1] ),
    .A2(net102),
    .B1(_0391_),
    .C1(net115),
    .X(_0392_));
 sky130_fd_sc_hd__o211a_1 _2486_ (.A1(net122),
    .A2(_0390_),
    .B1(_0392_),
    .C1(net94),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _2487_ (.A0(\as1802.regs[5][1] ),
    .A1(\as1802.regs[4][1] ),
    .S(net102),
    .X(_0394_));
 sky130_fd_sc_hd__and3_1 _2488_ (.A(\as1802.regs[7][1] ),
    .B(net151),
    .C(net143),
    .X(_0395_));
 sky130_fd_sc_hd__a211o_1 _2489_ (.A1(\as1802.regs[6][1] ),
    .A2(net102),
    .B1(_0395_),
    .C1(net115),
    .X(_0396_));
 sky130_fd_sc_hd__o211a_1 _2490_ (.A1(net122),
    .A2(_0394_),
    .B1(_0396_),
    .C1(net90),
    .X(_0397_));
 sky130_fd_sc_hd__o32ai_4 _2491_ (.A1(net85),
    .A2(_0393_),
    .A3(_0397_),
    .B1(_0384_),
    .B2(_0389_),
    .Y(_0398_));
 sky130_fd_sc_hd__nor2_1 _2492_ (.A(net82),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2_1 _2493_ (.A(net82),
    .B(_0398_),
    .Y(_0400_));
 sky130_fd_sc_hd__nand2b_2 _2494_ (.A_N(_0399_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__xnor2_1 _2495_ (.A(net165),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__mux2_1 _2496_ (.A0(\as1802.D[1] ),
    .A1(_0402_),
    .S(_2087_),
    .X(_0403_));
 sky130_fd_sc_hd__and2b_1 _2497_ (.A_N(net256),
    .B(\as1802.regs[10][1] ),
    .X(_0404_));
 sky130_fd_sc_hd__a21bo_1 _2498_ (.A1(net256),
    .A2(\as1802.regs[11][1] ),
    .B1_N(net245),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _2499_ (.A0(\as1802.regs[8][1] ),
    .A1(\as1802.regs[9][1] ),
    .S(net256),
    .X(_0406_));
 sky130_fd_sc_hd__o221a_2 _2500_ (.A1(_0404_),
    .A2(_0405_),
    .B1(_0406_),
    .B2(net245),
    .C1(net198),
    .X(_0407_));
 sky130_fd_sc_hd__mux4_1 _2501_ (.A0(\as1802.regs[12][1] ),
    .A1(\as1802.regs[13][1] ),
    .A2(\as1802.regs[14][1] ),
    .A3(\as1802.regs[15][1] ),
    .S0(net256),
    .S1(net246),
    .X(_0408_));
 sky130_fd_sc_hd__a21o_1 _2502_ (.A1(net242),
    .A2(_0408_),
    .B1(net197),
    .X(_0409_));
 sky130_fd_sc_hd__mux4_1 _2503_ (.A0(\as1802.regs[0][1] ),
    .A1(\as1802.regs[1][1] ),
    .A2(\as1802.regs[2][1] ),
    .A3(\as1802.regs[3][1] ),
    .S0(net260),
    .S1(net249),
    .X(_0410_));
 sky130_fd_sc_hd__mux4_1 _2504_ (.A0(\as1802.regs[4][1] ),
    .A1(\as1802.regs[5][1] ),
    .A2(\as1802.regs[6][1] ),
    .A3(\as1802.regs[7][1] ),
    .S0(net261),
    .S1(net250),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _2505_ (.A0(_0410_),
    .A1(_0411_),
    .S(net243),
    .X(_0412_));
 sky130_fd_sc_hd__o22a_4 _2506_ (.A1(_0407_),
    .A2(_0409_),
    .B1(_0412_),
    .B2(net240),
    .X(_0413_));
 sky130_fd_sc_hd__nor2_1 _2507_ (.A(net155),
    .B(net164),
    .Y(_0414_));
 sky130_fd_sc_hd__a21o_1 _2508_ (.A1(net155),
    .A2(_0413_),
    .B1(_2065_),
    .X(_0415_));
 sky130_fd_sc_hd__a2bb2o_1 _2509_ (.A1_N(_0414_),
    .A2_N(_0415_),
    .B1(net208),
    .B2(_2065_),
    .X(_0416_));
 sky130_fd_sc_hd__nand2_1 _2510_ (.A(_2141_),
    .B(_0413_),
    .Y(_0417_));
 sky130_fd_sc_hd__xnor2_1 _2511_ (.A(_2141_),
    .B(net164),
    .Y(_0418_));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(_0416_),
    .A1(_0418_),
    .S(net133),
    .X(_0419_));
 sky130_fd_sc_hd__nand2_1 _2513_ (.A(net134),
    .B(_0413_),
    .Y(_0420_));
 sky130_fd_sc_hd__o211a_1 _2514_ (.A1(net134),
    .A2(_0419_),
    .B1(_0420_),
    .C1(_2070_),
    .X(_0421_));
 sky130_fd_sc_hd__a211o_1 _2515_ (.A1(net208),
    .A2(_2069_),
    .B1(_2148_),
    .C1(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__o211a_1 _2516_ (.A1(net126),
    .A2(_0418_),
    .B1(_0422_),
    .C1(net80),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(_2105_),
    .A1(_2109_),
    .S(_0401_),
    .X(_0424_));
 sky130_fd_sc_hd__a211o_1 _2518_ (.A1(net84),
    .A2(_0403_),
    .B1(_0424_),
    .C1(net131),
    .X(_0425_));
 sky130_fd_sc_hd__xnor2_1 _2519_ (.A(\as1802.regs[2][0] ),
    .B(\as1802.regs[2][1] ),
    .Y(_0426_));
 sky130_fd_sc_hd__o22a_4 _2520_ (.A1(_0423_),
    .A2(_0425_),
    .B1(_0426_),
    .B2(net129),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _2521_ (.A0(\as1802.regs[15][1] ),
    .A1(net66),
    .S(_2126_),
    .X(_0013_));
 sky130_fd_sc_hd__and3_1 _2522_ (.A(\as1802.regs[13][2] ),
    .B(net154),
    .C(net146),
    .X(_0428_));
 sky130_fd_sc_hd__a211o_1 _2523_ (.A1(\as1802.regs[12][2] ),
    .A2(net100),
    .B1(_0428_),
    .C1(net120),
    .X(_0429_));
 sky130_fd_sc_hd__and3_1 _2524_ (.A(\as1802.regs[15][2] ),
    .B(net148),
    .C(net140),
    .X(_0430_));
 sky130_fd_sc_hd__a211o_1 _2525_ (.A1(\as1802.regs[14][2] ),
    .A2(net96),
    .B1(_0430_),
    .C1(net112),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(\as1802.regs[9][2] ),
    .A1(\as1802.regs[8][2] ),
    .S(net101),
    .X(_0432_));
 sky130_fd_sc_hd__and3_1 _2527_ (.A(\as1802.regs[11][2] ),
    .B(net150),
    .C(net142),
    .X(_0433_));
 sky130_fd_sc_hd__a211o_1 _2528_ (.A1(\as1802.regs[10][2] ),
    .A2(net101),
    .B1(_0433_),
    .C1(net114),
    .X(_0434_));
 sky130_fd_sc_hd__o211a_2 _2529_ (.A1(net121),
    .A2(_0432_),
    .B1(_0434_),
    .C1(net94),
    .X(_0435_));
 sky130_fd_sc_hd__a31o_2 _2530_ (.A1(net89),
    .A2(_0429_),
    .A3(_0431_),
    .B1(net87),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(\as1802.regs[1][2] ),
    .A1(\as1802.regs[0][2] ),
    .S(net103),
    .X(_0437_));
 sky130_fd_sc_hd__and3_1 _2532_ (.A(\as1802.regs[3][2] ),
    .B(net151),
    .C(net143),
    .X(_0438_));
 sky130_fd_sc_hd__a211o_1 _2533_ (.A1(\as1802.regs[2][2] ),
    .A2(net103),
    .B1(_0438_),
    .C1(net114),
    .X(_0439_));
 sky130_fd_sc_hd__o211a_1 _2534_ (.A1(net121),
    .A2(_0437_),
    .B1(_0439_),
    .C1(net94),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _2535_ (.A0(\as1802.regs[5][2] ),
    .A1(\as1802.regs[4][2] ),
    .S(net102),
    .X(_0441_));
 sky130_fd_sc_hd__and3_1 _2536_ (.A(\as1802.regs[7][2] ),
    .B(net151),
    .C(net143),
    .X(_0442_));
 sky130_fd_sc_hd__a211o_1 _2537_ (.A1(\as1802.regs[6][2] ),
    .A2(net102),
    .B1(_0442_),
    .C1(net115),
    .X(_0443_));
 sky130_fd_sc_hd__o211a_2 _2538_ (.A1(net121),
    .A2(_0441_),
    .B1(_0443_),
    .C1(net90),
    .X(_0444_));
 sky130_fd_sc_hd__o32ai_4 _2539_ (.A1(net85),
    .A2(_0440_),
    .A3(_0444_),
    .B1(_0435_),
    .B2(_0436_),
    .Y(_0445_));
 sky130_fd_sc_hd__xnor2_1 _2540_ (.A(_0400_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__xnor2_1 _2541_ (.A(_0399_),
    .B(_0445_),
    .Y(_0447_));
 sky130_fd_sc_hd__mux4_1 _2542_ (.A0(\as1802.regs[12][2] ),
    .A1(\as1802.regs[13][2] ),
    .A2(\as1802.regs[14][2] ),
    .A3(\as1802.regs[15][2] ),
    .S0(net257),
    .S1(net246),
    .X(_0448_));
 sky130_fd_sc_hd__nand2_2 _2543_ (.A(net242),
    .B(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__and2b_1 _2544_ (.A_N(net260),
    .B(\as1802.regs[10][2] ),
    .X(_0450_));
 sky130_fd_sc_hd__a21bo_1 _2545_ (.A1(net260),
    .A2(\as1802.regs[11][2] ),
    .B1_N(net249),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_2 _2546_ (.A0(\as1802.regs[8][2] ),
    .A1(\as1802.regs[9][2] ),
    .S(net260),
    .X(_0452_));
 sky130_fd_sc_hd__o221ai_4 _2547_ (.A1(_0450_),
    .A2(_0451_),
    .B1(_0452_),
    .B2(net249),
    .C1(net198),
    .Y(_0453_));
 sky130_fd_sc_hd__mux4_1 _2548_ (.A0(\as1802.regs[0][2] ),
    .A1(\as1802.regs[1][2] ),
    .A2(\as1802.regs[2][2] ),
    .A3(\as1802.regs[3][2] ),
    .S0(net261),
    .S1(net250),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_2 _2549_ (.A(net198),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__mux4_2 _2550_ (.A0(\as1802.regs[4][2] ),
    .A1(\as1802.regs[5][2] ),
    .A2(\as1802.regs[6][2] ),
    .A3(\as1802.regs[7][2] ),
    .S0(net260),
    .S1(net249),
    .X(_0456_));
 sky130_fd_sc_hd__a21oi_4 _2551_ (.A1(net243),
    .A2(_0456_),
    .B1(net239),
    .Y(_0457_));
 sky130_fd_sc_hd__a32oi_4 _2552_ (.A1(net240),
    .A2(_0449_),
    .A3(_0453_),
    .B1(_0455_),
    .B2(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__a32o_4 _2553_ (.A1(net240),
    .A2(_0449_),
    .A3(_0453_),
    .B1(_0455_),
    .B2(_0457_),
    .X(_0459_));
 sky130_fd_sc_hd__xnor2_1 _2554_ (.A(net164),
    .B(_0458_),
    .Y(_0460_));
 sky130_fd_sc_hd__mux2_2 _2555_ (.A0(_0459_),
    .A1(_0460_),
    .S(_0417_),
    .X(_0461_));
 sky130_fd_sc_hd__or3b_2 _2556_ (.A(_0459_),
    .B(net156),
    .C_N(_0413_),
    .X(_0462_));
 sky130_fd_sc_hd__a21o_1 _2557_ (.A1(net155),
    .A2(net164),
    .B1(_0458_),
    .X(_0463_));
 sky130_fd_sc_hd__and3_1 _2558_ (.A(_2066_),
    .B(_0462_),
    .C(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__a211oi_1 _2559_ (.A1(net206),
    .A2(_2065_),
    .B1(_0464_),
    .C1(net133),
    .Y(_0465_));
 sky130_fd_sc_hd__a211o_1 _2560_ (.A1(net133),
    .A2(_0461_),
    .B1(_0465_),
    .C1(net134),
    .X(_0466_));
 sky130_fd_sc_hd__o211a_1 _2561_ (.A1(_2049_),
    .A2(_0460_),
    .B1(_0466_),
    .C1(_2070_),
    .X(_0467_));
 sky130_fd_sc_hd__o21ai_2 _2562_ (.A1(net206),
    .A2(_2070_),
    .B1(net126),
    .Y(_0468_));
 sky130_fd_sc_hd__o22ai_4 _2563_ (.A1(net127),
    .A2(_0461_),
    .B1(_0467_),
    .B2(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__a221o_1 _2564_ (.A1(_2102_),
    .A2(_0447_),
    .B1(_0469_),
    .B2(net81),
    .C1(net131),
    .X(_0470_));
 sky130_fd_sc_hd__o21bai_1 _2565_ (.A1(_2097_),
    .A2(_0446_),
    .B1_N(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__nor2_1 _2566_ (.A(_0380_),
    .B(_0446_),
    .Y(_0472_));
 sky130_fd_sc_hd__a211o_1 _2567_ (.A1(_0380_),
    .A2(_0447_),
    .B1(_0472_),
    .C1(_2086_),
    .X(_0473_));
 sky130_fd_sc_hd__o211a_1 _2568_ (.A1(net215),
    .A2(_2087_),
    .B1(net83),
    .C1(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__o21a_1 _2569_ (.A1(\as1802.regs[2][0] ),
    .A2(\as1802.regs[2][1] ),
    .B1(\as1802.regs[2][2] ),
    .X(_0475_));
 sky130_fd_sc_hd__or3_1 _2570_ (.A(\as1802.regs[2][0] ),
    .B(\as1802.regs[2][1] ),
    .C(\as1802.regs[2][2] ),
    .X(_0476_));
 sky130_fd_sc_hd__or3b_1 _2571_ (.A(net129),
    .B(_0475_),
    .C_N(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__o21a_1 _2572_ (.A1(_0471_),
    .A2(_0474_),
    .B1(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(\as1802.regs[15][2] ),
    .A1(net64),
    .S(_2126_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(\as1802.regs[9][3] ),
    .A1(\as1802.regs[8][3] ),
    .S(net104),
    .X(_0479_));
 sky130_fd_sc_hd__and3_1 _2575_ (.A(\as1802.regs[11][3] ),
    .B(net151),
    .C(net143),
    .X(_0480_));
 sky130_fd_sc_hd__a211o_1 _2576_ (.A1(\as1802.regs[10][3] ),
    .A2(net104),
    .B1(_0480_),
    .C1(net115),
    .X(_0481_));
 sky130_fd_sc_hd__o211a_4 _2577_ (.A1(net119),
    .A2(_0479_),
    .B1(_0481_),
    .C1(net94),
    .X(_0482_));
 sky130_fd_sc_hd__and3_1 _2578_ (.A(\as1802.regs[15][3] ),
    .B(net149),
    .C(net141),
    .X(_0483_));
 sky130_fd_sc_hd__a211o_1 _2579_ (.A1(\as1802.regs[14][3] ),
    .A2(net99),
    .B1(_0483_),
    .C1(net113),
    .X(_0484_));
 sky130_fd_sc_hd__and3_1 _2580_ (.A(\as1802.regs[13][3] ),
    .B(net149),
    .C(net141),
    .X(_0485_));
 sky130_fd_sc_hd__a211o_1 _2581_ (.A1(\as1802.regs[12][3] ),
    .A2(net99),
    .B1(_0485_),
    .C1(net119),
    .X(_0486_));
 sky130_fd_sc_hd__a31o_4 _2582_ (.A1(net89),
    .A2(_0484_),
    .A3(_0486_),
    .B1(net87),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _2583_ (.A0(\as1802.regs[1][3] ),
    .A1(\as1802.regs[0][3] ),
    .S(net104),
    .X(_0488_));
 sky130_fd_sc_hd__and3_1 _2584_ (.A(\as1802.regs[3][3] ),
    .B(net151),
    .C(net143),
    .X(_0489_));
 sky130_fd_sc_hd__a211o_1 _2585_ (.A1(\as1802.regs[2][3] ),
    .A2(net104),
    .B1(_0489_),
    .C1(net115),
    .X(_0490_));
 sky130_fd_sc_hd__o211a_2 _2586_ (.A1(net122),
    .A2(_0488_),
    .B1(_0490_),
    .C1(net94),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(\as1802.regs[5][3] ),
    .A1(\as1802.regs[4][3] ),
    .S(net103),
    .X(_0492_));
 sky130_fd_sc_hd__and3_1 _2588_ (.A(\as1802.regs[7][3] ),
    .B(net150),
    .C(net142),
    .X(_0493_));
 sky130_fd_sc_hd__a211o_1 _2589_ (.A1(\as1802.regs[6][3] ),
    .A2(net103),
    .B1(_0493_),
    .C1(net114),
    .X(_0494_));
 sky130_fd_sc_hd__o211a_2 _2590_ (.A1(net121),
    .A2(_0492_),
    .B1(_0494_),
    .C1(net90),
    .X(_0495_));
 sky130_fd_sc_hd__o32a_4 _2591_ (.A1(net85),
    .A2(_0491_),
    .A3(_0495_),
    .B1(_0482_),
    .B2(_0487_),
    .X(_0496_));
 sky130_fd_sc_hd__o32ai_4 _2592_ (.A1(net86),
    .A2(_0491_),
    .A3(_0495_),
    .B1(_0482_),
    .B2(_0487_),
    .Y(_0497_));
 sky130_fd_sc_hd__and4_2 _2593_ (.A(net82),
    .B(_0398_),
    .C(_0445_),
    .D(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__a31o_1 _2594_ (.A1(net82),
    .A2(_0398_),
    .A3(_0445_),
    .B1(_0497_),
    .X(_0499_));
 sky130_fd_sc_hd__nand2b_1 _2595_ (.A_N(_0498_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__and2b_1 _2596_ (.A_N(net262),
    .B(\as1802.regs[10][3] ),
    .X(_0501_));
 sky130_fd_sc_hd__a21bo_1 _2597_ (.A1(net262),
    .A2(\as1802.regs[11][3] ),
    .B1_N(net251),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _2598_ (.A0(\as1802.regs[8][3] ),
    .A1(\as1802.regs[9][3] ),
    .S(net262),
    .X(_0503_));
 sky130_fd_sc_hd__o221a_1 _2599_ (.A1(_0501_),
    .A2(_0502_),
    .B1(_0503_),
    .B2(net251),
    .C1(net199),
    .X(_0504_));
 sky130_fd_sc_hd__mux4_1 _2600_ (.A0(\as1802.regs[12][3] ),
    .A1(\as1802.regs[13][3] ),
    .A2(\as1802.regs[14][3] ),
    .A3(\as1802.regs[15][3] ),
    .S0(net259),
    .S1(net247),
    .X(_0505_));
 sky130_fd_sc_hd__a21o_1 _2601_ (.A1(net242),
    .A2(_0505_),
    .B1(net197),
    .X(_0506_));
 sky130_fd_sc_hd__mux4_1 _2602_ (.A0(\as1802.regs[0][3] ),
    .A1(\as1802.regs[1][3] ),
    .A2(\as1802.regs[2][3] ),
    .A3(\as1802.regs[3][3] ),
    .S0(net262),
    .S1(net251),
    .X(_0507_));
 sky130_fd_sc_hd__mux4_1 _2603_ (.A0(\as1802.regs[4][3] ),
    .A1(\as1802.regs[5][3] ),
    .A2(\as1802.regs[6][3] ),
    .A3(\as1802.regs[7][3] ),
    .S0(net261),
    .S1(net249),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_2 _2604_ (.A0(_0507_),
    .A1(_0508_),
    .S(net243),
    .X(_0509_));
 sky130_fd_sc_hd__o22a_4 _2605_ (.A1(_0504_),
    .A2(_0506_),
    .B1(_0509_),
    .B2(net240),
    .X(_0510_));
 sky130_fd_sc_hd__and3_1 _2606_ (.A(net164),
    .B(_0458_),
    .C(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__xnor2_1 _2607_ (.A(_0462_),
    .B(_0510_),
    .Y(_0512_));
 sky130_fd_sc_hd__mux2_1 _2608_ (.A0(net33),
    .A1(_0512_),
    .S(_2066_),
    .X(_0513_));
 sky130_fd_sc_hd__a21oi_1 _2609_ (.A1(net164),
    .A2(_0458_),
    .B1(_0510_),
    .Y(_0514_));
 sky130_fd_sc_hd__nor2_1 _2610_ (.A(_0511_),
    .B(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(_0510_),
    .A1(_0515_),
    .S(_2140_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _2612_ (.A0(_0513_),
    .A1(_0516_),
    .S(net133),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _2613_ (.A0(_0515_),
    .A1(_0517_),
    .S(_2049_),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _2614_ (.A0(net33),
    .A1(_0518_),
    .S(_2072_),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _2615_ (.A0(_0516_),
    .A1(_0519_),
    .S(net127),
    .X(_0520_));
 sky130_fd_sc_hd__o31a_1 _2616_ (.A1(net82),
    .A2(_0398_),
    .A3(_0445_),
    .B1(_0497_),
    .X(_0521_));
 sky130_fd_sc_hd__or4_4 _2617_ (.A(net82),
    .B(_0398_),
    .C(_0445_),
    .D(_0497_),
    .X(_0522_));
 sky130_fd_sc_hd__nor2_1 _2618_ (.A(net214),
    .B(_2087_),
    .Y(_0523_));
 sky130_fd_sc_hd__and2b_1 _2619_ (.A_N(_0521_),
    .B(_0522_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _2620_ (.A0(_0500_),
    .A1(_0524_),
    .S(_0380_),
    .X(_0525_));
 sky130_fd_sc_hd__o21ai_1 _2621_ (.A1(_2086_),
    .A2(_0525_),
    .B1(net84),
    .Y(_0526_));
 sky130_fd_sc_hd__or2_1 _2622_ (.A(_2096_),
    .B(_0524_),
    .X(_0527_));
 sky130_fd_sc_hd__o211a_1 _2623_ (.A1(_2097_),
    .A2(_0500_),
    .B1(_0527_),
    .C1(_2107_),
    .X(_0528_));
 sky130_fd_sc_hd__a211o_1 _2624_ (.A1(net81),
    .A2(_0520_),
    .B1(_0528_),
    .C1(net131),
    .X(_0529_));
 sky130_fd_sc_hd__o21bai_2 _2625_ (.A1(_0523_),
    .A2(_0526_),
    .B1_N(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__o31a_1 _2626_ (.A1(\as1802.regs[2][0] ),
    .A2(\as1802.regs[2][1] ),
    .A3(\as1802.regs[2][2] ),
    .B1(\as1802.regs[2][3] ),
    .X(_0531_));
 sky130_fd_sc_hd__or4_4 _2627_ (.A(\as1802.regs[2][0] ),
    .B(\as1802.regs[2][1] ),
    .C(\as1802.regs[2][2] ),
    .D(\as1802.regs[2][3] ),
    .X(_0532_));
 sky130_fd_sc_hd__inv_2 _2628_ (.A(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__o31a_2 _2629_ (.A1(net129),
    .A2(_0531_),
    .A3(_0533_),
    .B1(_0530_),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _2630_ (.A0(\as1802.regs[15][3] ),
    .A1(net62),
    .S(_2126_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _2631_ (.A0(\as1802.regs[11][4] ),
    .A1(\as1802.regs[10][4] ),
    .S(net96),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(\as1802.regs[9][4] ),
    .A1(\as1802.regs[8][4] ),
    .S(net96),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_1 _2633_ (.A0(_0535_),
    .A1(_0536_),
    .S(net112),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(\as1802.regs[15][4] ),
    .A1(\as1802.regs[14][4] ),
    .S(net96),
    .X(_0538_));
 sky130_fd_sc_hd__or2_1 _2635_ (.A(net112),
    .B(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(\as1802.regs[13][4] ),
    .A1(\as1802.regs[12][4] ),
    .S(net96),
    .X(_0540_));
 sky130_fd_sc_hd__o21a_1 _2637_ (.A1(net120),
    .A2(_0540_),
    .B1(net89),
    .X(_0541_));
 sky130_fd_sc_hd__a221o_4 _2638_ (.A1(net93),
    .A2(_0537_),
    .B1(_0539_),
    .B2(_0541_),
    .C1(net87),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_1 _2639_ (.A0(\as1802.regs[3][4] ),
    .A1(\as1802.regs[2][4] ),
    .S(net102),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _2640_ (.A0(\as1802.regs[1][4] ),
    .A1(\as1802.regs[0][4] ),
    .S(net102),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_1 _2641_ (.A0(_0543_),
    .A1(_0544_),
    .S(net114),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _2642_ (.A0(\as1802.regs[5][4] ),
    .A1(\as1802.regs[4][4] ),
    .S(net103),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _2643_ (.A0(\as1802.regs[7][4] ),
    .A1(\as1802.regs[6][4] ),
    .S(net103),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _2644_ (.A0(_0546_),
    .A1(_0547_),
    .S(net122),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(_0545_),
    .A1(_0548_),
    .S(net90),
    .X(_0549_));
 sky130_fd_sc_hd__o21ai_2 _2646_ (.A1(net85),
    .A2(_0549_),
    .B1(_0542_),
    .Y(_0550_));
 sky130_fd_sc_hd__or2_1 _2647_ (.A(_0522_),
    .B(net79),
    .X(_0551_));
 sky130_fd_sc_hd__nand2_1 _2648_ (.A(_0522_),
    .B(net79),
    .Y(_0552_));
 sky130_fd_sc_hd__nand2_1 _2649_ (.A(_0551_),
    .B(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__o21ai_1 _2650_ (.A1(net165),
    .A2(_0553_),
    .B1(_2087_),
    .Y(_0554_));
 sky130_fd_sc_hd__o211a_1 _2651_ (.A1(net213),
    .A2(_2085_),
    .B1(net84),
    .C1(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__nor2_1 _2652_ (.A(_2101_),
    .B(_0553_),
    .Y(_0556_));
 sky130_fd_sc_hd__nand2_1 _2653_ (.A(_0498_),
    .B(net78),
    .Y(_0557_));
 sky130_fd_sc_hd__or2_1 _2654_ (.A(_0498_),
    .B(net78),
    .X(_0558_));
 sky130_fd_sc_hd__nor2_4 _2655_ (.A(_2096_),
    .B(net165),
    .Y(_0559_));
 sky130_fd_sc_hd__a21oi_1 _2656_ (.A1(_0557_),
    .A2(_0558_),
    .B1(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__mux4_2 _2657_ (.A0(\as1802.regs[12][4] ),
    .A1(\as1802.regs[13][4] ),
    .A2(\as1802.regs[14][4] ),
    .A3(\as1802.regs[15][4] ),
    .S0(net256),
    .S1(net246),
    .X(_0561_));
 sky130_fd_sc_hd__nand2_2 _2658_ (.A(net243),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__and2b_1 _2659_ (.A_N(net256),
    .B(\as1802.regs[10][4] ),
    .X(_0563_));
 sky130_fd_sc_hd__a21bo_1 _2660_ (.A1(net256),
    .A2(\as1802.regs[11][4] ),
    .B1_N(net246),
    .X(_0564_));
 sky130_fd_sc_hd__mux2_2 _2661_ (.A0(\as1802.regs[8][4] ),
    .A1(\as1802.regs[9][4] ),
    .S(net256),
    .X(_0565_));
 sky130_fd_sc_hd__o221ai_4 _2662_ (.A1(_0563_),
    .A2(_0564_),
    .B1(_0565_),
    .B2(net246),
    .C1(net198),
    .Y(_0566_));
 sky130_fd_sc_hd__mux4_2 _2663_ (.A0(\as1802.regs[0][4] ),
    .A1(\as1802.regs[1][4] ),
    .A2(\as1802.regs[2][4] ),
    .A3(\as1802.regs[3][4] ),
    .S0(net261),
    .S1(net250),
    .X(_0567_));
 sky130_fd_sc_hd__nand2_2 _2664_ (.A(net199),
    .B(_0567_),
    .Y(_0568_));
 sky130_fd_sc_hd__mux4_2 _2665_ (.A0(\as1802.regs[4][4] ),
    .A1(\as1802.regs[5][4] ),
    .A2(\as1802.regs[6][4] ),
    .A3(\as1802.regs[7][4] ),
    .S0(net261),
    .S1(net250),
    .X(_0569_));
 sky130_fd_sc_hd__a21oi_4 _2666_ (.A1(net243),
    .A2(_0569_),
    .B1(net240),
    .Y(_0570_));
 sky130_fd_sc_hd__a32oi_4 _2667_ (.A1(net240),
    .A2(_0562_),
    .A3(_0566_),
    .B1(_0568_),
    .B2(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__a32o_4 _2668_ (.A1(net240),
    .A2(_0562_),
    .A3(_0566_),
    .B1(_0568_),
    .B2(_0570_),
    .X(_0572_));
 sky130_fd_sc_hd__and4_4 _2669_ (.A(net164),
    .B(_0458_),
    .C(_0510_),
    .D(_0571_),
    .X(_0573_));
 sky130_fd_sc_hd__nor2_1 _2670_ (.A(_0511_),
    .B(_0571_),
    .Y(_0574_));
 sky130_fd_sc_hd__or2_1 _2671_ (.A(_0573_),
    .B(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _2672_ (.A0(_0572_),
    .A1(_0575_),
    .S(_2140_),
    .X(_0576_));
 sky130_fd_sc_hd__a21oi_1 _2673_ (.A1(net155),
    .A2(_0511_),
    .B1(_0571_),
    .Y(_0577_));
 sky130_fd_sc_hd__a21o_1 _2674_ (.A1(net155),
    .A2(_0573_),
    .B1(_0577_),
    .X(_0578_));
 sky130_fd_sc_hd__nor2_1 _2675_ (.A(net34),
    .B(_2066_),
    .Y(_0579_));
 sky130_fd_sc_hd__a211o_1 _2676_ (.A1(_2066_),
    .A2(_0578_),
    .B1(_0579_),
    .C1(net133),
    .X(_0580_));
 sky130_fd_sc_hd__o211a_1 _2677_ (.A1(_2056_),
    .A2(_0576_),
    .B1(_0580_),
    .C1(_2049_),
    .X(_0581_));
 sky130_fd_sc_hd__and2_1 _2678_ (.A(net134),
    .B(_0575_),
    .X(_0582_));
 sky130_fd_sc_hd__o21ai_1 _2679_ (.A1(_0581_),
    .A2(_0582_),
    .B1(_2072_),
    .Y(_0583_));
 sky130_fd_sc_hd__o211a_1 _2680_ (.A1(net34),
    .A2(_2070_),
    .B1(net127),
    .C1(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__nor2_1 _2681_ (.A(net127),
    .B(_0576_),
    .Y(_0585_));
 sky130_fd_sc_hd__or3_1 _2682_ (.A(net132),
    .B(_0584_),
    .C(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__o2bb2a_1 _2683_ (.A1_N(net132),
    .A2_N(_0578_),
    .B1(_2073_),
    .B2(_2075_),
    .X(_0587_));
 sky130_fd_sc_hd__a2111o_1 _2684_ (.A1(_0586_),
    .A2(_0587_),
    .B1(net130),
    .C1(_0556_),
    .D1(_0560_),
    .X(_0588_));
 sky130_fd_sc_hd__or2_1 _2685_ (.A(_0555_),
    .B(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__and2_1 _2686_ (.A(\as1802.regs[2][4] ),
    .B(_0532_),
    .X(_0590_));
 sky130_fd_sc_hd__nor2_1 _2687_ (.A(\as1802.regs[2][4] ),
    .B(_0532_),
    .Y(_0591_));
 sky130_fd_sc_hd__o31a_2 _2688_ (.A1(net129),
    .A2(_0590_),
    .A3(_0591_),
    .B1(_0589_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _2689_ (.A0(\as1802.regs[15][4] ),
    .A1(net60),
    .S(_2126_),
    .X(_0016_));
 sky130_fd_sc_hd__and3_1 _2690_ (.A(\as1802.regs[13][5] ),
    .B(net147),
    .C(net139),
    .X(_0593_));
 sky130_fd_sc_hd__a211o_1 _2691_ (.A1(\as1802.regs[12][5] ),
    .A2(net97),
    .B1(_0593_),
    .C1(net120),
    .X(_0594_));
 sky130_fd_sc_hd__and3_1 _2692_ (.A(\as1802.regs[15][5] ),
    .B(net147),
    .C(net139),
    .X(_0595_));
 sky130_fd_sc_hd__a211o_1 _2693_ (.A1(\as1802.regs[14][5] ),
    .A2(net97),
    .B1(_0595_),
    .C1(net112),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _2694_ (.A0(\as1802.regs[9][5] ),
    .A1(\as1802.regs[8][5] ),
    .S(net97),
    .X(_0597_));
 sky130_fd_sc_hd__and3_1 _2695_ (.A(\as1802.regs[11][5] ),
    .B(net147),
    .C(net139),
    .X(_0598_));
 sky130_fd_sc_hd__a211o_1 _2696_ (.A1(\as1802.regs[10][5] ),
    .A2(net97),
    .B1(_0598_),
    .C1(net112),
    .X(_0599_));
 sky130_fd_sc_hd__o211a_2 _2697_ (.A1(net120),
    .A2(_0597_),
    .B1(_0599_),
    .C1(net93),
    .X(_0600_));
 sky130_fd_sc_hd__a31o_2 _2698_ (.A1(net89),
    .A2(_0594_),
    .A3(_0596_),
    .B1(net87),
    .X(_0601_));
 sky130_fd_sc_hd__mux2_1 _2699_ (.A0(\as1802.regs[1][5] ),
    .A1(\as1802.regs[0][5] ),
    .S(net102),
    .X(_0602_));
 sky130_fd_sc_hd__and3_1 _2700_ (.A(\as1802.regs[3][5] ),
    .B(net150),
    .C(net142),
    .X(_0603_));
 sky130_fd_sc_hd__a211o_1 _2701_ (.A1(\as1802.regs[2][5] ),
    .A2(net102),
    .B1(_0603_),
    .C1(net115),
    .X(_0604_));
 sky130_fd_sc_hd__o211a_1 _2702_ (.A1(net122),
    .A2(_0602_),
    .B1(_0604_),
    .C1(net94),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_1 _2703_ (.A0(\as1802.regs[5][5] ),
    .A1(\as1802.regs[4][5] ),
    .S(net101),
    .X(_0606_));
 sky130_fd_sc_hd__and3_1 _2704_ (.A(\as1802.regs[7][5] ),
    .B(net150),
    .C(net142),
    .X(_0607_));
 sky130_fd_sc_hd__a211o_1 _2705_ (.A1(\as1802.regs[6][5] ),
    .A2(net101),
    .B1(_0607_),
    .C1(net114),
    .X(_0608_));
 sky130_fd_sc_hd__o211a_1 _2706_ (.A1(net121),
    .A2(_0606_),
    .B1(_0608_),
    .C1(net90),
    .X(_0609_));
 sky130_fd_sc_hd__o32ai_4 _2707_ (.A1(net85),
    .A2(_0605_),
    .A3(_0609_),
    .B1(_0600_),
    .B2(_0601_),
    .Y(_0610_));
 sky130_fd_sc_hd__or3_4 _2708_ (.A(_0522_),
    .B(net79),
    .C(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__nand2_1 _2709_ (.A(_0551_),
    .B(_0610_),
    .Y(_0612_));
 sky130_fd_sc_hd__nand2_1 _2710_ (.A(_0611_),
    .B(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__o21a_1 _2711_ (.A1(_0379_),
    .A2(_0613_),
    .B1(_2087_),
    .X(_0614_));
 sky130_fd_sc_hd__nor2_1 _2712_ (.A(net212),
    .B(_2085_),
    .Y(_0615_));
 sky130_fd_sc_hd__and3_1 _2713_ (.A(_0498_),
    .B(net78),
    .C(_0610_),
    .X(_0616_));
 sky130_fd_sc_hd__a21oi_1 _2714_ (.A1(_0498_),
    .A2(net78),
    .B1(_0610_),
    .Y(_0617_));
 sky130_fd_sc_hd__nor2_1 _2715_ (.A(_0616_),
    .B(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__and2b_1 _2716_ (.A_N(net257),
    .B(\as1802.regs[10][5] ),
    .X(_0619_));
 sky130_fd_sc_hd__a21bo_1 _2717_ (.A1(net257),
    .A2(\as1802.regs[11][5] ),
    .B1_N(net245),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _2718_ (.A0(\as1802.regs[8][5] ),
    .A1(\as1802.regs[9][5] ),
    .S(net257),
    .X(_0621_));
 sky130_fd_sc_hd__o221a_1 _2719_ (.A1(_0619_),
    .A2(_0620_),
    .B1(_0621_),
    .B2(net245),
    .C1(net198),
    .X(_0622_));
 sky130_fd_sc_hd__mux4_1 _2720_ (.A0(\as1802.regs[12][5] ),
    .A1(\as1802.regs[13][5] ),
    .A2(\as1802.regs[14][5] ),
    .A3(\as1802.regs[15][5] ),
    .S0(net257),
    .S1(net245),
    .X(_0623_));
 sky130_fd_sc_hd__a21o_1 _2721_ (.A1(net242),
    .A2(_0623_),
    .B1(net197),
    .X(_0624_));
 sky130_fd_sc_hd__mux4_1 _2722_ (.A0(\as1802.regs[0][5] ),
    .A1(\as1802.regs[1][5] ),
    .A2(\as1802.regs[2][5] ),
    .A3(\as1802.regs[3][5] ),
    .S0(net261),
    .S1(net250),
    .X(_0625_));
 sky130_fd_sc_hd__mux4_1 _2723_ (.A0(\as1802.regs[4][5] ),
    .A1(\as1802.regs[5][5] ),
    .A2(\as1802.regs[6][5] ),
    .A3(\as1802.regs[7][5] ),
    .S0(net260),
    .S1(net249),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_2 _2724_ (.A0(_0625_),
    .A1(_0626_),
    .S(net243),
    .X(_0627_));
 sky130_fd_sc_hd__o22a_4 _2725_ (.A1(_0622_),
    .A2(_0624_),
    .B1(_0627_),
    .B2(net239),
    .X(_0628_));
 sky130_fd_sc_hd__nand2_2 _2726_ (.A(_0573_),
    .B(net163),
    .Y(_0629_));
 sky130_fd_sc_hd__nor2_1 _2727_ (.A(net156),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__a21o_1 _2728_ (.A1(_2139_),
    .A2(_0573_),
    .B1(net163),
    .X(_0631_));
 sky130_fd_sc_hd__o21a_1 _2729_ (.A1(net156),
    .A2(_0629_),
    .B1(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__or2_1 _2730_ (.A(net35),
    .B(_2066_),
    .X(_0633_));
 sky130_fd_sc_hd__o211a_1 _2731_ (.A1(_2065_),
    .A2(_0632_),
    .B1(_0633_),
    .C1(_2056_),
    .X(_0634_));
 sky130_fd_sc_hd__or2_1 _2732_ (.A(_0573_),
    .B(net163),
    .X(_0635_));
 sky130_fd_sc_hd__and2_1 _2733_ (.A(_0629_),
    .B(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _2734_ (.A0(_0628_),
    .A1(_0636_),
    .S(_2140_),
    .X(_0637_));
 sky130_fd_sc_hd__a211o_1 _2735_ (.A1(net133),
    .A2(_0637_),
    .B1(_0634_),
    .C1(net134),
    .X(_0638_));
 sky130_fd_sc_hd__o21a_1 _2736_ (.A1(_2049_),
    .A2(_0636_),
    .B1(_2061_),
    .X(_0639_));
 sky130_fd_sc_hd__a21o_1 _2737_ (.A1(_2060_),
    .A2(_0632_),
    .B1(_2069_),
    .X(_0640_));
 sky130_fd_sc_hd__a21o_1 _2738_ (.A1(_0638_),
    .A2(_0639_),
    .B1(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__o211a_1 _2739_ (.A1(net35),
    .A2(_2070_),
    .B1(net127),
    .C1(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__a21o_1 _2740_ (.A1(_2148_),
    .A2(_0637_),
    .B1(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__a21oi_1 _2741_ (.A1(net80),
    .A2(_0643_),
    .B1(net130),
    .Y(_0644_));
 sky130_fd_sc_hd__o221a_1 _2742_ (.A1(_2101_),
    .A2(_0613_),
    .B1(_0618_),
    .B2(_0559_),
    .C1(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__o31a_2 _2743_ (.A1(_2089_),
    .A2(_0614_),
    .A3(_0615_),
    .B1(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__o21ai_2 _2744_ (.A1(\as1802.regs[2][4] ),
    .A2(_0532_),
    .B1(\as1802.regs[2][5] ),
    .Y(_0647_));
 sky130_fd_sc_hd__or3_4 _2745_ (.A(\as1802.regs[2][4] ),
    .B(\as1802.regs[2][5] ),
    .C(_0532_),
    .X(_0648_));
 sky130_fd_sc_hd__a31oi_4 _2746_ (.A1(net131),
    .A2(_0647_),
    .A3(_0648_),
    .B1(_0646_),
    .Y(_0649_));
 sky130_fd_sc_hd__mux2_1 _2747_ (.A0(\as1802.regs[15][5] ),
    .A1(net58),
    .S(_2126_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _2748_ (.A0(\as1802.regs[9][6] ),
    .A1(\as1802.regs[8][6] ),
    .S(net100),
    .X(_0650_));
 sky130_fd_sc_hd__and3_1 _2749_ (.A(\as1802.regs[11][6] ),
    .B(net149),
    .C(net141),
    .X(_0651_));
 sky130_fd_sc_hd__a211o_1 _2750_ (.A1(\as1802.regs[10][6] ),
    .A2(net98),
    .B1(_0651_),
    .C1(net118),
    .X(_0652_));
 sky130_fd_sc_hd__o211a_2 _2751_ (.A1(net119),
    .A2(_0650_),
    .B1(_0652_),
    .C1(net93),
    .X(_0653_));
 sky130_fd_sc_hd__and3_1 _2752_ (.A(\as1802.regs[15][6] ),
    .B(net149),
    .C(net141),
    .X(_0654_));
 sky130_fd_sc_hd__a211o_1 _2753_ (.A1(\as1802.regs[14][6] ),
    .A2(net98),
    .B1(_0654_),
    .C1(net112),
    .X(_0655_));
 sky130_fd_sc_hd__and3_1 _2754_ (.A(\as1802.regs[13][6] ),
    .B(net149),
    .C(net141),
    .X(_0656_));
 sky130_fd_sc_hd__a211o_1 _2755_ (.A1(\as1802.regs[12][6] ),
    .A2(net98),
    .B1(_0656_),
    .C1(net119),
    .X(_0657_));
 sky130_fd_sc_hd__a31o_2 _2756_ (.A1(net90),
    .A2(_0655_),
    .A3(_0657_),
    .B1(net87),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_1 _2757_ (.A0(\as1802.regs[1][6] ),
    .A1(\as1802.regs[0][6] ),
    .S(net104),
    .X(_0659_));
 sky130_fd_sc_hd__and3_1 _2758_ (.A(\as1802.regs[3][6] ),
    .B(net151),
    .C(net143),
    .X(_0660_));
 sky130_fd_sc_hd__a211o_1 _2759_ (.A1(\as1802.regs[2][6] ),
    .A2(net104),
    .B1(_0660_),
    .C1(net115),
    .X(_0661_));
 sky130_fd_sc_hd__o211a_1 _2760_ (.A1(net122),
    .A2(_0659_),
    .B1(_0661_),
    .C1(net93),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_1 _2761_ (.A0(\as1802.regs[5][6] ),
    .A1(\as1802.regs[4][6] ),
    .S(net103),
    .X(_0663_));
 sky130_fd_sc_hd__and3_1 _2762_ (.A(\as1802.regs[7][6] ),
    .B(net150),
    .C(net142),
    .X(_0664_));
 sky130_fd_sc_hd__a211o_1 _2763_ (.A1(\as1802.regs[6][6] ),
    .A2(net103),
    .B1(_0664_),
    .C1(net114),
    .X(_0665_));
 sky130_fd_sc_hd__o211a_1 _2764_ (.A1(net121),
    .A2(_0663_),
    .B1(_0665_),
    .C1(net90),
    .X(_0666_));
 sky130_fd_sc_hd__o32ai_4 _2765_ (.A1(net85),
    .A2(_0662_),
    .A3(_0666_),
    .B1(_0653_),
    .B2(_0658_),
    .Y(_0667_));
 sky130_fd_sc_hd__xnor2_1 _2766_ (.A(_0611_),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__o21ai_1 _2767_ (.A1(_0379_),
    .A2(_0668_),
    .B1(_2087_),
    .Y(_0669_));
 sky130_fd_sc_hd__o211a_1 _2768_ (.A1(\as1802.D[6] ),
    .A2(_2085_),
    .B1(net84),
    .C1(_0669_),
    .X(_0670_));
 sky130_fd_sc_hd__mux4_2 _2769_ (.A0(\as1802.regs[12][6] ),
    .A1(\as1802.regs[13][6] ),
    .A2(\as1802.regs[14][6] ),
    .A3(\as1802.regs[15][6] ),
    .S0(net258),
    .S1(net245),
    .X(_0671_));
 sky130_fd_sc_hd__and2b_1 _2770_ (.A_N(net258),
    .B(\as1802.regs[10][6] ),
    .X(_0672_));
 sky130_fd_sc_hd__a21bo_1 _2771_ (.A1(net258),
    .A2(\as1802.regs[11][6] ),
    .B1_N(net247),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_1 _2772_ (.A0(\as1802.regs[8][6] ),
    .A1(\as1802.regs[9][6] ),
    .S(net259),
    .X(_0674_));
 sky130_fd_sc_hd__o221a_1 _2773_ (.A1(_0672_),
    .A2(_0673_),
    .B1(_0674_),
    .B2(net247),
    .C1(net198),
    .X(_0675_));
 sky130_fd_sc_hd__a211o_4 _2774_ (.A1(net242),
    .A2(_0671_),
    .B1(_0675_),
    .C1(net197),
    .X(_0676_));
 sky130_fd_sc_hd__mux4_1 _2775_ (.A0(\as1802.regs[4][6] ),
    .A1(\as1802.regs[5][6] ),
    .A2(\as1802.regs[6][6] ),
    .A3(\as1802.regs[7][6] ),
    .S0(net261),
    .S1(net250),
    .X(_0677_));
 sky130_fd_sc_hd__mux4_1 _2776_ (.A0(\as1802.regs[0][6] ),
    .A1(\as1802.regs[1][6] ),
    .A2(\as1802.regs[2][6] ),
    .A3(\as1802.regs[3][6] ),
    .S0(net262),
    .S1(net251),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_4 _2777_ (.A0(_0677_),
    .A1(_0678_),
    .S(net199),
    .X(_0679_));
 sky130_fd_sc_hd__o21a_4 _2778_ (.A1(net239),
    .A2(_0679_),
    .B1(_0676_),
    .X(_0680_));
 sky130_fd_sc_hd__o21ai_4 _2779_ (.A1(net239),
    .A2(_0679_),
    .B1(_0676_),
    .Y(_0681_));
 sky130_fd_sc_hd__xnor2_1 _2780_ (.A(_0630_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__or2_1 _2781_ (.A(net205),
    .B(_2066_),
    .X(_0683_));
 sky130_fd_sc_hd__o211a_1 _2782_ (.A1(_2065_),
    .A2(_0682_),
    .B1(_0683_),
    .C1(_2056_),
    .X(_0684_));
 sky130_fd_sc_hd__xnor2_1 _2783_ (.A(_0629_),
    .B(_0680_),
    .Y(_0685_));
 sky130_fd_sc_hd__mux2_1 _2784_ (.A0(_0680_),
    .A1(_0685_),
    .S(_2140_),
    .X(_0686_));
 sky130_fd_sc_hd__a211o_1 _2785_ (.A1(net133),
    .A2(_0686_),
    .B1(_0684_),
    .C1(net134),
    .X(_0687_));
 sky130_fd_sc_hd__o211a_1 _2786_ (.A1(_2049_),
    .A2(_0685_),
    .B1(_0687_),
    .C1(_2061_),
    .X(_0688_));
 sky130_fd_sc_hd__a211o_1 _2787_ (.A1(_2060_),
    .A2(_0682_),
    .B1(_0688_),
    .C1(_2069_),
    .X(_0689_));
 sky130_fd_sc_hd__o21a_1 _2788_ (.A1(net205),
    .A2(_2072_),
    .B1(net127),
    .X(_0690_));
 sky130_fd_sc_hd__a22o_1 _2789_ (.A1(_2148_),
    .A2(_0686_),
    .B1(_0689_),
    .B2(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__xor2_1 _2790_ (.A(_0616_),
    .B(_0667_),
    .X(_0692_));
 sky130_fd_sc_hd__o221a_1 _2791_ (.A1(_2101_),
    .A2(_0668_),
    .B1(_0692_),
    .B2(_0559_),
    .C1(net129),
    .X(_0693_));
 sky130_fd_sc_hd__a21bo_1 _2792_ (.A1(_2078_),
    .A2(_0691_),
    .B1_N(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__nor2_1 _2793_ (.A(_0670_),
    .B(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hd__or2_2 _2794_ (.A(\as1802.regs[2][6] ),
    .B(_0648_),
    .X(_0696_));
 sky130_fd_sc_hd__a21oi_1 _2795_ (.A1(\as1802.regs[2][6] ),
    .A2(_0648_),
    .B1(net129),
    .Y(_0697_));
 sky130_fd_sc_hd__a21oi_2 _2796_ (.A1(_0696_),
    .A2(_0697_),
    .B1(_0695_),
    .Y(_0698_));
 sky130_fd_sc_hd__mux2_1 _2797_ (.A0(\as1802.regs[15][6] ),
    .A1(net56),
    .S(_2126_),
    .X(_0018_));
 sky130_fd_sc_hd__and3_1 _2798_ (.A(\as1802.regs[11][7] ),
    .B(net148),
    .C(net140),
    .X(_0699_));
 sky130_fd_sc_hd__a211o_1 _2799_ (.A1(\as1802.regs[10][7] ),
    .A2(net100),
    .B1(_0699_),
    .C1(net112),
    .X(_0700_));
 sky130_fd_sc_hd__mux2_1 _2800_ (.A0(\as1802.regs[9][7] ),
    .A1(\as1802.regs[8][7] ),
    .S(net100),
    .X(_0701_));
 sky130_fd_sc_hd__o211a_2 _2801_ (.A1(net120),
    .A2(_0701_),
    .B1(_0700_),
    .C1(net93),
    .X(_0702_));
 sky130_fd_sc_hd__and3_1 _2802_ (.A(\as1802.regs[15][7] ),
    .B(net147),
    .C(net139),
    .X(_0703_));
 sky130_fd_sc_hd__a211o_1 _2803_ (.A1(\as1802.regs[14][7] ),
    .A2(net97),
    .B1(_0703_),
    .C1(net112),
    .X(_0704_));
 sky130_fd_sc_hd__and3_1 _2804_ (.A(\as1802.regs[13][7] ),
    .B(net147),
    .C(net139),
    .X(_0705_));
 sky130_fd_sc_hd__a211o_1 _2805_ (.A1(\as1802.regs[12][7] ),
    .A2(net97),
    .B1(_0705_),
    .C1(net120),
    .X(_0706_));
 sky130_fd_sc_hd__a31o_2 _2806_ (.A1(net89),
    .A2(_0704_),
    .A3(_0706_),
    .B1(net87),
    .X(_0707_));
 sky130_fd_sc_hd__and3_1 _2807_ (.A(\as1802.regs[7][7] ),
    .B(net150),
    .C(net142),
    .X(_0708_));
 sky130_fd_sc_hd__a211o_1 _2808_ (.A1(\as1802.regs[6][7] ),
    .A2(net101),
    .B1(_0708_),
    .C1(net114),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _2809_ (.A0(\as1802.regs[5][7] ),
    .A1(\as1802.regs[4][7] ),
    .S(net101),
    .X(_0710_));
 sky130_fd_sc_hd__o211a_2 _2810_ (.A1(net121),
    .A2(_0710_),
    .B1(_0709_),
    .C1(net90),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _2811_ (.A0(\as1802.regs[1][7] ),
    .A1(\as1802.regs[0][7] ),
    .S(net104),
    .X(_0712_));
 sky130_fd_sc_hd__and3_1 _2812_ (.A(\as1802.regs[3][7] ),
    .B(net150),
    .C(net142),
    .X(_0713_));
 sky130_fd_sc_hd__a211o_1 _2813_ (.A1(\as1802.regs[2][7] ),
    .A2(net101),
    .B1(_0713_),
    .C1(net114),
    .X(_0714_));
 sky130_fd_sc_hd__o211a_1 _2814_ (.A1(net121),
    .A2(_0712_),
    .B1(_0714_),
    .C1(net94),
    .X(_0715_));
 sky130_fd_sc_hd__o32ai_4 _2815_ (.A1(net85),
    .A2(_0711_),
    .A3(_0715_),
    .B1(_0702_),
    .B2(_0707_),
    .Y(_0716_));
 sky130_fd_sc_hd__or2_1 _2816_ (.A(_0667_),
    .B(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__or4_4 _2817_ (.A(_0522_),
    .B(net78),
    .C(_0610_),
    .D(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__o21a_1 _2818_ (.A1(_0611_),
    .A2(_0667_),
    .B1(_0716_),
    .X(_0719_));
 sky130_fd_sc_hd__o21bai_2 _2819_ (.A1(_0611_),
    .A2(_0717_),
    .B1_N(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__o21a_1 _2820_ (.A1(net165),
    .A2(_0720_),
    .B1(_2087_),
    .X(_0721_));
 sky130_fd_sc_hd__o21ai_1 _2821_ (.A1(net211),
    .A2(_2085_),
    .B1(net83),
    .Y(_0722_));
 sky130_fd_sc_hd__and2b_1 _2822_ (.A_N(net256),
    .B(\as1802.regs[10][7] ),
    .X(_0723_));
 sky130_fd_sc_hd__a21bo_1 _2823_ (.A1(net263),
    .A2(\as1802.regs[11][7] ),
    .B1_N(net245),
    .X(_0724_));
 sky130_fd_sc_hd__mux2_1 _2824_ (.A0(\as1802.regs[8][7] ),
    .A1(\as1802.regs[9][7] ),
    .S(net257),
    .X(_0725_));
 sky130_fd_sc_hd__o221a_1 _2825_ (.A1(_0723_),
    .A2(_0724_),
    .B1(_0725_),
    .B2(net246),
    .C1(net198),
    .X(_0726_));
 sky130_fd_sc_hd__mux4_1 _2826_ (.A0(\as1802.regs[12][7] ),
    .A1(\as1802.regs[13][7] ),
    .A2(\as1802.regs[14][7] ),
    .A3(\as1802.regs[15][7] ),
    .S0(net257),
    .S1(net245),
    .X(_0727_));
 sky130_fd_sc_hd__a21o_1 _2827_ (.A1(net242),
    .A2(_0727_),
    .B1(net197),
    .X(_0728_));
 sky130_fd_sc_hd__mux4_1 _2828_ (.A0(\as1802.regs[0][7] ),
    .A1(\as1802.regs[1][7] ),
    .A2(\as1802.regs[2][7] ),
    .A3(\as1802.regs[3][7] ),
    .S0(net260),
    .S1(net249),
    .X(_0729_));
 sky130_fd_sc_hd__mux4_1 _2829_ (.A0(\as1802.regs[4][7] ),
    .A1(\as1802.regs[5][7] ),
    .A2(\as1802.regs[6][7] ),
    .A3(\as1802.regs[7][7] ),
    .S0(net260),
    .S1(net249),
    .X(_0730_));
 sky130_fd_sc_hd__mux2_1 _2830_ (.A0(_0729_),
    .A1(_0730_),
    .S(_0002_),
    .X(_0731_));
 sky130_fd_sc_hd__o22a_4 _2831_ (.A1(_0726_),
    .A2(_0728_),
    .B1(_0731_),
    .B2(net239),
    .X(_0732_));
 sky130_fd_sc_hd__a41o_1 _2832_ (.A1(net155),
    .A2(_0573_),
    .A3(net163),
    .A4(_0680_),
    .B1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__and4_1 _2833_ (.A(_0573_),
    .B(net163),
    .C(_0680_),
    .D(_0732_),
    .X(_0734_));
 sky130_fd_sc_hd__nand4_4 _2834_ (.A(_0573_),
    .B(net163),
    .C(_0680_),
    .D(_0732_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_1 _2835_ (.A(net156),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__o21ai_1 _2836_ (.A1(net156),
    .A2(_0735_),
    .B1(_0733_),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _2837_ (.A(_2066_),
    .B(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__o21a_1 _2838_ (.A1(net204),
    .A2(_2066_),
    .B1(_2056_),
    .X(_0739_));
 sky130_fd_sc_hd__a31o_1 _2839_ (.A1(_0573_),
    .A2(net163),
    .A3(_0680_),
    .B1(_0732_),
    .X(_0740_));
 sky130_fd_sc_hd__and2_1 _2840_ (.A(_0735_),
    .B(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _2841_ (.A0(_0732_),
    .A1(_0741_),
    .S(_2140_),
    .X(_0742_));
 sky130_fd_sc_hd__a221o_1 _2842_ (.A1(_0738_),
    .A2(_0739_),
    .B1(_0742_),
    .B2(net133),
    .C1(net134),
    .X(_0743_));
 sky130_fd_sc_hd__o211a_1 _2843_ (.A1(_2049_),
    .A2(_0741_),
    .B1(_0743_),
    .C1(_2061_),
    .X(_0744_));
 sky130_fd_sc_hd__nor2_1 _2844_ (.A(_2061_),
    .B(_0737_),
    .Y(_0745_));
 sky130_fd_sc_hd__o32a_1 _2845_ (.A1(_2069_),
    .A2(_0744_),
    .A3(_0745_),
    .B1(_2072_),
    .B2(net204),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_1 _2846_ (.A0(_0742_),
    .A1(_0746_),
    .S(net127),
    .X(_0747_));
 sky130_fd_sc_hd__a21oi_1 _2847_ (.A1(net81),
    .A2(_0747_),
    .B1(net130),
    .Y(_0748_));
 sky130_fd_sc_hd__and3_1 _2848_ (.A(_0610_),
    .B(_0667_),
    .C(_0716_),
    .X(_0749_));
 sky130_fd_sc_hd__and3_1 _2849_ (.A(_0498_),
    .B(net78),
    .C(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__a21o_1 _2850_ (.A1(_0616_),
    .A2(_0667_),
    .B1(_0716_),
    .X(_0751_));
 sky130_fd_sc_hd__and2b_1 _2851_ (.A_N(_0750_),
    .B(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__o221a_1 _2852_ (.A1(_2101_),
    .A2(_0720_),
    .B1(_0752_),
    .B2(_0559_),
    .C1(_0748_),
    .X(_0753_));
 sky130_fd_sc_hd__o21a_2 _2853_ (.A1(_0721_),
    .A2(_0722_),
    .B1(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__or2_2 _2854_ (.A(\as1802.regs[2][7] ),
    .B(_0696_),
    .X(_0755_));
 sky130_fd_sc_hd__a21oi_2 _2855_ (.A1(\as1802.regs[2][7] ),
    .A2(_0696_),
    .B1(net128),
    .Y(_0756_));
 sky130_fd_sc_hd__a21oi_4 _2856_ (.A1(_0755_),
    .A2(_0756_),
    .B1(_0754_),
    .Y(_0757_));
 sky130_fd_sc_hd__mux2_1 _2857_ (.A0(\as1802.regs[15][7] ),
    .A1(net54),
    .S(_2126_),
    .X(_0019_));
 sky130_fd_sc_hd__nor2_8 _2858_ (.A(_2111_),
    .B(_2115_),
    .Y(_0758_));
 sky130_fd_sc_hd__nor2_4 _2859_ (.A(_2120_),
    .B(_2122_),
    .Y(_0759_));
 sky130_fd_sc_hd__or4_1 _2860_ (.A(net282),
    .B(_2076_),
    .C(_2080_),
    .D(_2084_),
    .X(_0760_));
 sky130_fd_sc_hd__or3_2 _2861_ (.A(_2062_),
    .B(_2114_),
    .C(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__and3_4 _2862_ (.A(_0758_),
    .B(_0759_),
    .C(net70),
    .X(_0762_));
 sky130_fd_sc_hd__and3_1 _2863_ (.A(\as1802.regs[11][8] ),
    .B(net154),
    .C(net146),
    .X(_0763_));
 sky130_fd_sc_hd__a211o_1 _2864_ (.A1(\as1802.regs[10][8] ),
    .A2(net99),
    .B1(_0763_),
    .C1(net113),
    .X(_0764_));
 sky130_fd_sc_hd__mux2_1 _2865_ (.A0(\as1802.regs[9][8] ),
    .A1(\as1802.regs[8][8] ),
    .S(net99),
    .X(_0765_));
 sky130_fd_sc_hd__o211a_2 _2866_ (.A1(net119),
    .A2(_0765_),
    .B1(_0764_),
    .C1(net93),
    .X(_0766_));
 sky130_fd_sc_hd__and3_1 _2867_ (.A(\as1802.regs[15][8] ),
    .B(net152),
    .C(net144),
    .X(_0767_));
 sky130_fd_sc_hd__a211o_1 _2868_ (.A1(\as1802.regs[14][8] ),
    .A2(net99),
    .B1(_0767_),
    .C1(net113),
    .X(_0768_));
 sky130_fd_sc_hd__and3_1 _2869_ (.A(\as1802.regs[13][8] ),
    .B(net152),
    .C(net144),
    .X(_0769_));
 sky130_fd_sc_hd__a211o_1 _2870_ (.A1(\as1802.regs[12][8] ),
    .A2(net98),
    .B1(_0769_),
    .C1(net119),
    .X(_0770_));
 sky130_fd_sc_hd__a31o_2 _2871_ (.A1(net89),
    .A2(_0768_),
    .A3(_0770_),
    .B1(net87),
    .X(_0771_));
 sky130_fd_sc_hd__and3_1 _2872_ (.A(\as1802.regs[3][8] ),
    .B(net152),
    .C(net144),
    .X(_0772_));
 sky130_fd_sc_hd__a211o_1 _2873_ (.A1(\as1802.regs[2][8] ),
    .A2(net99),
    .B1(_0772_),
    .C1(net113),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _2874_ (.A0(\as1802.regs[1][8] ),
    .A1(\as1802.regs[0][8] ),
    .S(net99),
    .X(_0774_));
 sky130_fd_sc_hd__o211a_2 _2875_ (.A1(net125),
    .A2(_0774_),
    .B1(_0773_),
    .C1(net95),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _2876_ (.A0(\as1802.regs[5][8] ),
    .A1(\as1802.regs[4][8] ),
    .S(net106),
    .X(_0776_));
 sky130_fd_sc_hd__and3_1 _2877_ (.A(\as1802.regs[7][8] ),
    .B(net152),
    .C(net144),
    .X(_0777_));
 sky130_fd_sc_hd__a211o_1 _2878_ (.A1(\as1802.regs[6][8] ),
    .A2(net106),
    .B1(_0777_),
    .C1(net116),
    .X(_0778_));
 sky130_fd_sc_hd__o211a_2 _2879_ (.A1(net124),
    .A2(_0776_),
    .B1(_0778_),
    .C1(net91),
    .X(_0779_));
 sky130_fd_sc_hd__o32a_4 _2880_ (.A1(net86),
    .A2(_0775_),
    .A3(_0779_),
    .B1(_0766_),
    .B2(_0771_),
    .X(_0780_));
 sky130_fd_sc_hd__o32ai_4 _2881_ (.A1(net86),
    .A2(_0775_),
    .A3(_0779_),
    .B1(_0766_),
    .B2(_0771_),
    .Y(_0781_));
 sky130_fd_sc_hd__o211a_1 _2882_ (.A1(net219),
    .A2(_2081_),
    .B1(net83),
    .C1(_0380_),
    .X(_0782_));
 sky130_fd_sc_hd__o22a_1 _2883_ (.A1(_0718_),
    .A2(_0781_),
    .B1(_0782_),
    .B2(_2102_),
    .X(_0783_));
 sky130_fd_sc_hd__a21boi_1 _2884_ (.A1(_0718_),
    .A2(_0781_),
    .B1_N(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__and4_4 _2885_ (.A(_0498_),
    .B(net78),
    .C(_0749_),
    .D(_0781_),
    .X(_0785_));
 sky130_fd_sc_hd__nor2_1 _2886_ (.A(_0750_),
    .B(_0781_),
    .Y(_0786_));
 sky130_fd_sc_hd__o21ba_1 _2887_ (.A1(_0785_),
    .A2(_0786_),
    .B1_N(_0559_),
    .X(_0787_));
 sky130_fd_sc_hd__mux4_1 _2888_ (.A0(\as1802.regs[12][8] ),
    .A1(\as1802.regs[13][8] ),
    .A2(\as1802.regs[14][8] ),
    .A3(\as1802.regs[15][8] ),
    .S0(net258),
    .S1(net247),
    .X(_0788_));
 sky130_fd_sc_hd__nand2_1 _2889_ (.A(net243),
    .B(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__mux2_1 _2890_ (.A0(\as1802.regs[10][8] ),
    .A1(\as1802.regs[11][8] ),
    .S(net259),
    .X(_0790_));
 sky130_fd_sc_hd__inv_2 _2891_ (.A(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__mux2_1 _2892_ (.A0(\as1802.regs[8][8] ),
    .A1(\as1802.regs[9][8] ),
    .S(net259),
    .X(_0792_));
 sky130_fd_sc_hd__nor2_1 _2893_ (.A(net247),
    .B(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__a211o_1 _2894_ (.A1(net248),
    .A2(_0791_),
    .B1(_0793_),
    .C1(net243),
    .X(_0794_));
 sky130_fd_sc_hd__mux4_1 _2895_ (.A0(\as1802.regs[0][8] ),
    .A1(\as1802.regs[1][8] ),
    .A2(\as1802.regs[2][8] ),
    .A3(\as1802.regs[3][8] ),
    .S0(net258),
    .S1(net247),
    .X(_0795_));
 sky130_fd_sc_hd__mux4_1 _2896_ (.A0(\as1802.regs[4][8] ),
    .A1(\as1802.regs[5][8] ),
    .A2(\as1802.regs[6][8] ),
    .A3(\as1802.regs[7][8] ),
    .S0(net265),
    .S1(net255),
    .X(_0796_));
 sky130_fd_sc_hd__mux2_1 _2897_ (.A0(_0795_),
    .A1(_0796_),
    .S(net244),
    .X(_0797_));
 sky130_fd_sc_hd__nor2_1 _2898_ (.A(net239),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__a31o_4 _2899_ (.A1(net239),
    .A2(_0789_),
    .A3(_0794_),
    .B1(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__clkinv_2 _2900_ (.A(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__xnor2_2 _2901_ (.A(_0736_),
    .B(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__a21oi_4 _2902_ (.A1(net200),
    .A2(net133),
    .B1(_2048_),
    .Y(_0802_));
 sky130_fd_sc_hd__a21o_2 _2903_ (.A1(net200),
    .A2(_2055_),
    .B1(_2048_),
    .X(_0803_));
 sky130_fd_sc_hd__nand2_1 _2904_ (.A(net134),
    .B(_0734_),
    .Y(_0804_));
 sky130_fd_sc_hd__and3_1 _2905_ (.A(_0799_),
    .B(_0803_),
    .C(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__nor2_1 _2906_ (.A(_0799_),
    .B(_0804_),
    .Y(_0806_));
 sky130_fd_sc_hd__or3_1 _2907_ (.A(_2075_),
    .B(_0805_),
    .C(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__a21oi_1 _2908_ (.A1(_0801_),
    .A2(_0802_),
    .B1(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__a211o_1 _2909_ (.A1(net16),
    .A2(_2075_),
    .B1(_2148_),
    .C1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__nor2_1 _2910_ (.A(net200),
    .B(_0801_),
    .Y(_0810_));
 sky130_fd_sc_hd__nor2_1 _2911_ (.A(net228),
    .B(_0799_),
    .Y(_0811_));
 sky130_fd_sc_hd__o31a_1 _2912_ (.A1(net126),
    .A2(_0810_),
    .A3(_0811_),
    .B1(_0809_),
    .X(_0812_));
 sky130_fd_sc_hd__nand2_1 _2913_ (.A(net132),
    .B(_0801_),
    .Y(_0813_));
 sky130_fd_sc_hd__o211a_1 _2914_ (.A1(net132),
    .A2(_0812_),
    .B1(_0813_),
    .C1(net80),
    .X(_0814_));
 sky130_fd_sc_hd__a2111o_1 _2915_ (.A1(net219),
    .A2(_2080_),
    .B1(net130),
    .C1(_0787_),
    .D1(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__nor2_1 _2916_ (.A(_0784_),
    .B(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__or2_2 _2917_ (.A(\as1802.regs[2][8] ),
    .B(_0755_),
    .X(_0817_));
 sky130_fd_sc_hd__a21oi_1 _2918_ (.A1(\as1802.regs[2][8] ),
    .A2(_0755_),
    .B1(net128),
    .Y(_0818_));
 sky130_fd_sc_hd__a21oi_2 _2919_ (.A1(_0817_),
    .A2(_0818_),
    .B1(_0816_),
    .Y(_0819_));
 sky130_fd_sc_hd__mux2_1 _2920_ (.A0(\as1802.regs[10][8] ),
    .A1(net52),
    .S(_0762_),
    .X(_0020_));
 sky130_fd_sc_hd__and3_1 _2921_ (.A(\as1802.regs[11][9] ),
    .B(net149),
    .C(net141),
    .X(_0820_));
 sky130_fd_sc_hd__a211o_1 _2922_ (.A1(\as1802.regs[10][9] ),
    .A2(net98),
    .B1(_0820_),
    .C1(net113),
    .X(_0821_));
 sky130_fd_sc_hd__mux2_1 _2923_ (.A0(\as1802.regs[9][9] ),
    .A1(\as1802.regs[8][9] ),
    .S(net98),
    .X(_0822_));
 sky130_fd_sc_hd__o211a_1 _2924_ (.A1(net119),
    .A2(_0822_),
    .B1(_0821_),
    .C1(net93),
    .X(_0823_));
 sky130_fd_sc_hd__and3_1 _2925_ (.A(\as1802.regs[15][9] ),
    .B(net149),
    .C(net141),
    .X(_0824_));
 sky130_fd_sc_hd__a211o_1 _2926_ (.A1(\as1802.regs[14][9] ),
    .A2(net98),
    .B1(_0824_),
    .C1(net113),
    .X(_0825_));
 sky130_fd_sc_hd__and3_1 _2927_ (.A(\as1802.regs[13][9] ),
    .B(net149),
    .C(net141),
    .X(_0826_));
 sky130_fd_sc_hd__a211o_1 _2928_ (.A1(\as1802.regs[12][9] ),
    .A2(net98),
    .B1(_0826_),
    .C1(net119),
    .X(_0827_));
 sky130_fd_sc_hd__a31o_1 _2929_ (.A1(net89),
    .A2(_0825_),
    .A3(_0827_),
    .B1(net87),
    .X(_0828_));
 sky130_fd_sc_hd__and3_1 _2930_ (.A(\as1802.regs[3][9] ),
    .B(net152),
    .C(net144),
    .X(_0829_));
 sky130_fd_sc_hd__a211o_1 _2931_ (.A1(\as1802.regs[2][9] ),
    .A2(net99),
    .B1(_0829_),
    .C1(net118),
    .X(_0830_));
 sky130_fd_sc_hd__mux2_1 _2932_ (.A0(\as1802.regs[1][9] ),
    .A1(\as1802.regs[0][9] ),
    .S(net99),
    .X(_0831_));
 sky130_fd_sc_hd__o211a_2 _2933_ (.A1(net119),
    .A2(_0831_),
    .B1(_0830_),
    .C1(net93),
    .X(_0832_));
 sky130_fd_sc_hd__mux2_1 _2934_ (.A0(\as1802.regs[5][9] ),
    .A1(\as1802.regs[4][9] ),
    .S(net98),
    .X(_0833_));
 sky130_fd_sc_hd__and3_1 _2935_ (.A(\as1802.regs[7][9] ),
    .B(net152),
    .C(net144),
    .X(_0834_));
 sky130_fd_sc_hd__a211o_1 _2936_ (.A1(\as1802.regs[6][9] ),
    .A2(net98),
    .B1(_0834_),
    .C1(net113),
    .X(_0835_));
 sky130_fd_sc_hd__o211a_1 _2937_ (.A1(net119),
    .A2(_0833_),
    .B1(_0835_),
    .C1(net89),
    .X(_0836_));
 sky130_fd_sc_hd__o32ai_4 _2938_ (.A1(net85),
    .A2(_0832_),
    .A3(_0836_),
    .B1(_0823_),
    .B2(_0828_),
    .Y(_0837_));
 sky130_fd_sc_hd__o21a_1 _2939_ (.A1(_0718_),
    .A2(_0781_),
    .B1(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__or2_2 _2940_ (.A(_0781_),
    .B(_0837_),
    .X(_0839_));
 sky130_fd_sc_hd__nor2_1 _2941_ (.A(_0718_),
    .B(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__or2_1 _2942_ (.A(_0838_),
    .B(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__o21a_1 _2943_ (.A1(net165),
    .A2(_0841_),
    .B1(_2081_),
    .X(_0842_));
 sky130_fd_sc_hd__o21ai_1 _2944_ (.A1(\as1802.D[1] ),
    .A2(_2081_),
    .B1(net83),
    .Y(_0843_));
 sky130_fd_sc_hd__xor2_1 _2945_ (.A(_0785_),
    .B(_0837_),
    .X(_0844_));
 sky130_fd_sc_hd__mux4_1 _2946_ (.A0(\as1802.regs[12][9] ),
    .A1(\as1802.regs[13][9] ),
    .A2(\as1802.regs[14][9] ),
    .A3(\as1802.regs[15][9] ),
    .S0(net258),
    .S1(net247),
    .X(_0845_));
 sky130_fd_sc_hd__and2_1 _2947_ (.A(net242),
    .B(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__and2b_1 _2948_ (.A_N(net258),
    .B(\as1802.regs[10][9] ),
    .X(_0847_));
 sky130_fd_sc_hd__a21bo_1 _2949_ (.A1(net258),
    .A2(\as1802.regs[11][9] ),
    .B1_N(net247),
    .X(_0848_));
 sky130_fd_sc_hd__mux2_1 _2950_ (.A0(\as1802.regs[8][9] ),
    .A1(\as1802.regs[9][9] ),
    .S(net258),
    .X(_0849_));
 sky130_fd_sc_hd__o221a_1 _2951_ (.A1(_0847_),
    .A2(_0848_),
    .B1(_0849_),
    .B2(net247),
    .C1(net198),
    .X(_0850_));
 sky130_fd_sc_hd__mux4_1 _2952_ (.A0(\as1802.regs[4][9] ),
    .A1(\as1802.regs[5][9] ),
    .A2(\as1802.regs[6][9] ),
    .A3(\as1802.regs[7][9] ),
    .S0(net258),
    .S1(net247),
    .X(_0851_));
 sky130_fd_sc_hd__and2_1 _2953_ (.A(net242),
    .B(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__mux4_2 _2954_ (.A0(\as1802.regs[0][9] ),
    .A1(\as1802.regs[1][9] ),
    .A2(\as1802.regs[2][9] ),
    .A3(\as1802.regs[3][9] ),
    .S0(net259),
    .S1(net248),
    .X(_0853_));
 sky130_fd_sc_hd__a21o_1 _2955_ (.A1(net198),
    .A2(_0853_),
    .B1(net239),
    .X(_0854_));
 sky130_fd_sc_hd__o32a_4 _2956_ (.A1(net197),
    .A2(_0846_),
    .A3(_0850_),
    .B1(_0852_),
    .B2(_0854_),
    .X(_0855_));
 sky130_fd_sc_hd__inv_2 _2957_ (.A(_0855_),
    .Y(_0856_));
 sky130_fd_sc_hd__nand2_1 _2958_ (.A(_0806_),
    .B(_0855_),
    .Y(_0857_));
 sky130_fd_sc_hd__or3_1 _2959_ (.A(_0802_),
    .B(_0806_),
    .C(_0855_),
    .X(_0858_));
 sky130_fd_sc_hd__a31o_1 _2960_ (.A1(_2139_),
    .A2(_0734_),
    .A3(_0800_),
    .B1(_0855_),
    .X(_0859_));
 sky130_fd_sc_hd__or4_4 _2961_ (.A(net156),
    .B(_0735_),
    .C(_0799_),
    .D(_0856_),
    .X(_0860_));
 sky130_fd_sc_hd__and2_1 _2962_ (.A(_0859_),
    .B(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__or2_1 _2963_ (.A(_0803_),
    .B(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__and4b_1 _2964_ (.A_N(_2076_),
    .B(_0857_),
    .C(_0858_),
    .D(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__a211o_1 _2965_ (.A1(net24),
    .A2(_2076_),
    .B1(_2150_),
    .C1(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _2966_ (.A0(_0855_),
    .A1(_0861_),
    .S(net227),
    .X(_0865_));
 sky130_fd_sc_hd__o21a_1 _2967_ (.A1(net126),
    .A2(_0865_),
    .B1(_0864_),
    .X(_0866_));
 sky130_fd_sc_hd__a21oi_1 _2968_ (.A1(net80),
    .A2(_0866_),
    .B1(net130),
    .Y(_0867_));
 sky130_fd_sc_hd__o221a_1 _2969_ (.A1(_2101_),
    .A2(_0841_),
    .B1(_0844_),
    .B2(_0559_),
    .C1(_0867_),
    .X(_0868_));
 sky130_fd_sc_hd__o21a_1 _2970_ (.A1(_0842_),
    .A2(_0843_),
    .B1(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__or2_2 _2971_ (.A(\as1802.regs[2][9] ),
    .B(_0817_),
    .X(_0870_));
 sky130_fd_sc_hd__a21oi_1 _2972_ (.A1(\as1802.regs[2][9] ),
    .A2(_0817_),
    .B1(net128),
    .Y(_0871_));
 sky130_fd_sc_hd__a21oi_1 _2973_ (.A1(_0870_),
    .A2(_0871_),
    .B1(_0869_),
    .Y(_0872_));
 sky130_fd_sc_hd__mux2_1 _2974_ (.A0(\as1802.regs[10][9] ),
    .A1(net50),
    .S(_0762_),
    .X(_0021_));
 sky130_fd_sc_hd__xnor2_1 _2975_ (.A(\as1802.regs[2][10] ),
    .B(_0870_),
    .Y(_0873_));
 sky130_fd_sc_hd__and3_1 _2976_ (.A(\as1802.regs[13][10] ),
    .B(net152),
    .C(net144),
    .X(_0874_));
 sky130_fd_sc_hd__a211o_1 _2977_ (.A1(\as1802.regs[12][10] ),
    .A2(net105),
    .B1(_0874_),
    .C1(net124),
    .X(_0875_));
 sky130_fd_sc_hd__and3_1 _2978_ (.A(\as1802.regs[15][10] ),
    .B(net152),
    .C(net144),
    .X(_0876_));
 sky130_fd_sc_hd__a211o_1 _2979_ (.A1(\as1802.regs[14][10] ),
    .A2(net105),
    .B1(_0876_),
    .C1(net116),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(\as1802.regs[9][10] ),
    .A1(\as1802.regs[8][10] ),
    .S(net105),
    .X(_0878_));
 sky130_fd_sc_hd__and3_1 _2981_ (.A(\as1802.regs[11][10] ),
    .B(net153),
    .C(net145),
    .X(_0879_));
 sky130_fd_sc_hd__a211o_1 _2982_ (.A1(\as1802.regs[10][10] ),
    .A2(net105),
    .B1(_0879_),
    .C1(net116),
    .X(_0880_));
 sky130_fd_sc_hd__o211a_1 _2983_ (.A1(net124),
    .A2(_0878_),
    .B1(_0880_),
    .C1(net95),
    .X(_0881_));
 sky130_fd_sc_hd__a31o_1 _2984_ (.A1(net91),
    .A2(_0875_),
    .A3(_0877_),
    .B1(net87),
    .X(_0882_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(\as1802.regs[1][10] ),
    .A1(\as1802.regs[0][10] ),
    .S(net105),
    .X(_0883_));
 sky130_fd_sc_hd__and3_1 _2986_ (.A(\as1802.regs[3][10] ),
    .B(net152),
    .C(net144),
    .X(_0884_));
 sky130_fd_sc_hd__a211o_1 _2987_ (.A1(\as1802.regs[2][10] ),
    .A2(net105),
    .B1(_0884_),
    .C1(net116),
    .X(_0885_));
 sky130_fd_sc_hd__o211a_1 _2988_ (.A1(net124),
    .A2(_0883_),
    .B1(_0885_),
    .C1(net95),
    .X(_0886_));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(\as1802.regs[5][10] ),
    .A1(\as1802.regs[4][10] ),
    .S(net105),
    .X(_0887_));
 sky130_fd_sc_hd__and3_1 _2990_ (.A(\as1802.regs[7][10] ),
    .B(net152),
    .C(net144),
    .X(_0888_));
 sky130_fd_sc_hd__a211o_1 _2991_ (.A1(\as1802.regs[6][10] ),
    .A2(net105),
    .B1(_0888_),
    .C1(net116),
    .X(_0889_));
 sky130_fd_sc_hd__o211a_1 _2992_ (.A1(net124),
    .A2(_0887_),
    .B1(_0889_),
    .C1(net91),
    .X(_0890_));
 sky130_fd_sc_hd__o32ai_4 _2993_ (.A1(net86),
    .A2(_0886_),
    .A3(_0890_),
    .B1(_0881_),
    .B2(_0882_),
    .Y(_0891_));
 sky130_fd_sc_hd__xnor2_1 _2994_ (.A(_0840_),
    .B(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__nand2_2 _2995_ (.A(_0837_),
    .B(_0891_),
    .Y(_0893_));
 sky130_fd_sc_hd__or3b_2 _2996_ (.A(_0780_),
    .B(_0893_),
    .C_N(_0750_),
    .X(_0894_));
 sky130_fd_sc_hd__a21o_1 _2997_ (.A1(_0785_),
    .A2(_0837_),
    .B1(_0891_),
    .X(_0895_));
 sky130_fd_sc_hd__a21oi_1 _2998_ (.A1(_0894_),
    .A2(_0895_),
    .B1(_0380_),
    .Y(_0896_));
 sky130_fd_sc_hd__a211o_1 _2999_ (.A1(_0380_),
    .A2(_0892_),
    .B1(_0896_),
    .C1(_2080_),
    .X(_0897_));
 sky130_fd_sc_hd__or2_1 _3000_ (.A(\as1802.D[2] ),
    .B(_2081_),
    .X(_0898_));
 sky130_fd_sc_hd__and2b_1 _3001_ (.A_N(net264),
    .B(\as1802.regs[10][10] ),
    .X(_0899_));
 sky130_fd_sc_hd__a21bo_1 _3002_ (.A1(net264),
    .A2(\as1802.regs[11][10] ),
    .B1_N(net252),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _3003_ (.A0(\as1802.regs[8][10] ),
    .A1(\as1802.regs[9][10] ),
    .S(net264),
    .X(_0901_));
 sky130_fd_sc_hd__o221a_1 _3004_ (.A1(_0899_),
    .A2(_0900_),
    .B1(_0901_),
    .B2(net252),
    .C1(net199),
    .X(_0902_));
 sky130_fd_sc_hd__mux4_1 _3005_ (.A0(\as1802.regs[12][10] ),
    .A1(\as1802.regs[13][10] ),
    .A2(\as1802.regs[14][10] ),
    .A3(\as1802.regs[15][10] ),
    .S0(net264),
    .S1(net252),
    .X(_0903_));
 sky130_fd_sc_hd__a21o_1 _3006_ (.A1(net244),
    .A2(_0903_),
    .B1(net197),
    .X(_0904_));
 sky130_fd_sc_hd__mux4_1 _3007_ (.A0(\as1802.regs[0][10] ),
    .A1(\as1802.regs[1][10] ),
    .A2(\as1802.regs[2][10] ),
    .A3(\as1802.regs[3][10] ),
    .S0(net264),
    .S1(net252),
    .X(_0905_));
 sky130_fd_sc_hd__mux4_1 _3008_ (.A0(\as1802.regs[4][10] ),
    .A1(\as1802.regs[5][10] ),
    .A2(\as1802.regs[6][10] ),
    .A3(\as1802.regs[7][10] ),
    .S0(net264),
    .S1(net252),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _3009_ (.A0(_0905_),
    .A1(_0906_),
    .S(net244),
    .X(_0907_));
 sky130_fd_sc_hd__o22a_4 _3010_ (.A1(_0902_),
    .A2(_0904_),
    .B1(_0907_),
    .B2(net241),
    .X(_0908_));
 sky130_fd_sc_hd__clkinv_2 _3011_ (.A(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__nand2_1 _3012_ (.A(_0860_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__or4_4 _3013_ (.A(_0735_),
    .B(_0799_),
    .C(_0856_),
    .D(_0909_),
    .X(_0911_));
 sky130_fd_sc_hd__o21a_1 _3014_ (.A1(net156),
    .A2(_0911_),
    .B1(_0910_),
    .X(_0912_));
 sky130_fd_sc_hd__or2_2 _3015_ (.A(_2049_),
    .B(_0911_),
    .X(_0913_));
 sky130_fd_sc_hd__a21oi_1 _3016_ (.A1(_0857_),
    .A2(_0909_),
    .B1(_0802_),
    .Y(_0914_));
 sky130_fd_sc_hd__a22o_1 _3017_ (.A1(_0802_),
    .A2(_0912_),
    .B1(_0913_),
    .B2(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_1 _3018_ (.A0(net206),
    .A1(_0915_),
    .S(_2077_),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _3019_ (.A0(_0908_),
    .A1(_0912_),
    .S(net228),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _3020_ (.A0(_0916_),
    .A1(_0917_),
    .S(_2148_),
    .X(_0918_));
 sky130_fd_sc_hd__a21oi_1 _3021_ (.A1(_0894_),
    .A2(_0895_),
    .B1(_2097_),
    .Y(_0919_));
 sky130_fd_sc_hd__a211o_1 _3022_ (.A1(_2097_),
    .A2(_0892_),
    .B1(_0919_),
    .C1(_2106_),
    .X(_0920_));
 sky130_fd_sc_hd__or2_1 _3023_ (.A(_2058_),
    .B(_0912_),
    .X(_0921_));
 sky130_fd_sc_hd__o211a_1 _3024_ (.A1(net132),
    .A2(_0918_),
    .B1(_0921_),
    .C1(net80),
    .X(_0922_));
 sky130_fd_sc_hd__a311o_1 _3025_ (.A1(net83),
    .A2(_0897_),
    .A3(_0898_),
    .B1(_0922_),
    .C1(_2107_),
    .X(_0923_));
 sky130_fd_sc_hd__a22o_1 _3026_ (.A1(net130),
    .A2(_0873_),
    .B1(_0920_),
    .B2(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_1 _3027_ (.A0(\as1802.regs[10][10] ),
    .A1(net48),
    .S(_0762_),
    .X(_0022_));
 sky130_fd_sc_hd__and2b_1 _3028_ (.A_N(net266),
    .B(\as1802.regs[10][11] ),
    .X(_0925_));
 sky130_fd_sc_hd__a21bo_1 _3029_ (.A1(net266),
    .A2(\as1802.regs[11][11] ),
    .B1_N(net253),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _3030_ (.A0(\as1802.regs[8][11] ),
    .A1(\as1802.regs[9][11] ),
    .S(net266),
    .X(_0927_));
 sky130_fd_sc_hd__o221a_1 _3031_ (.A1(_0925_),
    .A2(_0926_),
    .B1(_0927_),
    .B2(net253),
    .C1(net199),
    .X(_0928_));
 sky130_fd_sc_hd__mux4_1 _3032_ (.A0(\as1802.regs[12][11] ),
    .A1(\as1802.regs[13][11] ),
    .A2(\as1802.regs[14][11] ),
    .A3(\as1802.regs[15][11] ),
    .S0(net266),
    .S1(net253),
    .X(_0929_));
 sky130_fd_sc_hd__a21o_1 _3033_ (.A1(net244),
    .A2(_0929_),
    .B1(net197),
    .X(_0930_));
 sky130_fd_sc_hd__mux4_1 _3034_ (.A0(\as1802.regs[4][11] ),
    .A1(\as1802.regs[5][11] ),
    .A2(\as1802.regs[6][11] ),
    .A3(\as1802.regs[7][11] ),
    .S0(net266),
    .S1(net253),
    .X(_0931_));
 sky130_fd_sc_hd__mux4_2 _3035_ (.A0(\as1802.regs[0][11] ),
    .A1(\as1802.regs[1][11] ),
    .A2(\as1802.regs[2][11] ),
    .A3(\as1802.regs[3][11] ),
    .S0(net267),
    .S1(net254),
    .X(_0932_));
 sky130_fd_sc_hd__mux2_1 _3036_ (.A0(_0931_),
    .A1(_0932_),
    .S(net199),
    .X(_0933_));
 sky130_fd_sc_hd__o22a_4 _3037_ (.A1(_0928_),
    .A2(_0930_),
    .B1(_0933_),
    .B2(net241),
    .X(_0934_));
 sky130_fd_sc_hd__o21ba_1 _3038_ (.A1(net156),
    .A2(_0911_),
    .B1_N(_0934_),
    .X(_0935_));
 sky130_fd_sc_hd__and3b_1 _3039_ (.A_N(_0860_),
    .B(_0908_),
    .C(_0934_),
    .X(_0936_));
 sky130_fd_sc_hd__or2_2 _3040_ (.A(_0935_),
    .B(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__nor3b_1 _3041_ (.A(_2049_),
    .B(_0911_),
    .C_N(_0934_),
    .Y(_0938_));
 sky130_fd_sc_hd__nor2_1 _3042_ (.A(_0802_),
    .B(_0934_),
    .Y(_0939_));
 sky130_fd_sc_hd__a221o_1 _3043_ (.A1(_0802_),
    .A2(_0937_),
    .B1(_0939_),
    .B2(_0913_),
    .C1(_0938_),
    .X(_0940_));
 sky130_fd_sc_hd__nand2_1 _3044_ (.A(_2077_),
    .B(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__o211a_1 _3045_ (.A1(net33),
    .A2(_2077_),
    .B1(net126),
    .C1(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__nand2_1 _3046_ (.A(net227),
    .B(_0937_),
    .Y(_0943_));
 sky130_fd_sc_hd__o211a_1 _3047_ (.A1(net227),
    .A2(_0934_),
    .B1(_0943_),
    .C1(_2148_),
    .X(_0944_));
 sky130_fd_sc_hd__or3_1 _3048_ (.A(net132),
    .B(_0942_),
    .C(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__nand2_1 _3049_ (.A(net132),
    .B(_0937_),
    .Y(_0946_));
 sky130_fd_sc_hd__a31o_1 _3050_ (.A1(net80),
    .A2(_0945_),
    .A3(_0946_),
    .B1(net83),
    .X(_0947_));
 sky130_fd_sc_hd__mux2_1 _3051_ (.A0(\as1802.regs[9][11] ),
    .A1(\as1802.regs[8][11] ),
    .S(net108),
    .X(_0948_));
 sky130_fd_sc_hd__mux2_1 _3052_ (.A0(\as1802.regs[11][11] ),
    .A1(\as1802.regs[10][11] ),
    .S(net108),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_1 _3053_ (.A0(_0948_),
    .A1(_0949_),
    .S(net123),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _3054_ (.A0(\as1802.regs[15][11] ),
    .A1(\as1802.regs[14][11] ),
    .S(net107),
    .X(_0951_));
 sky130_fd_sc_hd__or2_1 _3055_ (.A(net117),
    .B(_0951_),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_1 _3056_ (.A0(\as1802.regs[13][11] ),
    .A1(\as1802.regs[12][11] ),
    .S(net107),
    .X(_0953_));
 sky130_fd_sc_hd__o21a_1 _3057_ (.A1(net123),
    .A2(_0953_),
    .B1(net91),
    .X(_0954_));
 sky130_fd_sc_hd__a221o_2 _3058_ (.A1(net95),
    .A2(_0950_),
    .B1(_0952_),
    .B2(_0954_),
    .C1(net88),
    .X(_0955_));
 sky130_fd_sc_hd__mux2_1 _3059_ (.A0(\as1802.regs[1][11] ),
    .A1(\as1802.regs[0][11] ),
    .S(net109),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _3060_ (.A0(\as1802.regs[3][11] ),
    .A1(\as1802.regs[2][11] ),
    .S(net109),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _3061_ (.A0(_0956_),
    .A1(_0957_),
    .S(net123),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _3062_ (.A0(\as1802.regs[5][11] ),
    .A1(\as1802.regs[4][11] ),
    .S(net107),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _3063_ (.A0(\as1802.regs[7][11] ),
    .A1(\as1802.regs[6][11] ),
    .S(net108),
    .X(_0960_));
 sky130_fd_sc_hd__mux2_1 _3064_ (.A0(_0959_),
    .A1(_0960_),
    .S(net123),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _3065_ (.A0(_0958_),
    .A1(_0961_),
    .S(net91),
    .X(_0962_));
 sky130_fd_sc_hd__o21a_4 _3066_ (.A1(net86),
    .A2(_0962_),
    .B1(_0955_),
    .X(_0963_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__nor2_4 _3068_ (.A(_0893_),
    .B(_0963_),
    .Y(_0965_));
 sky130_fd_sc_hd__nand2_1 _3069_ (.A(_0785_),
    .B(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__a21boi_1 _3070_ (.A1(_0894_),
    .A2(_0963_),
    .B1_N(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__o31ai_2 _3071_ (.A1(_0718_),
    .A2(_0839_),
    .A3(_0891_),
    .B1(_0964_),
    .Y(_0968_));
 sky130_fd_sc_hd__or3b_2 _3072_ (.A(_0839_),
    .B(_0891_),
    .C_N(_0963_),
    .X(_0969_));
 sky130_fd_sc_hd__or2_2 _3073_ (.A(_0718_),
    .B(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__nand2_1 _3074_ (.A(_0968_),
    .B(_0970_),
    .Y(_0971_));
 sky130_fd_sc_hd__a21oi_1 _3075_ (.A1(_0968_),
    .A2(_0970_),
    .B1(net165),
    .Y(_0972_));
 sky130_fd_sc_hd__a211o_1 _3076_ (.A1(net165),
    .A2(_0967_),
    .B1(_0972_),
    .C1(_2080_),
    .X(_0973_));
 sky130_fd_sc_hd__a21oi_1 _3077_ (.A1(net214),
    .A2(_2080_),
    .B1(_2089_),
    .Y(_0974_));
 sky130_fd_sc_hd__a21bo_1 _3078_ (.A1(_0973_),
    .A2(_0974_),
    .B1_N(_0947_),
    .X(_0975_));
 sky130_fd_sc_hd__o221a_1 _3079_ (.A1(_2097_),
    .A2(_0967_),
    .B1(_0971_),
    .B2(_2101_),
    .C1(net128),
    .X(_0976_));
 sky130_fd_sc_hd__or3_1 _3080_ (.A(\as1802.regs[2][10] ),
    .B(\as1802.regs[2][11] ),
    .C(_0870_),
    .X(_0977_));
 sky130_fd_sc_hd__o21ai_1 _3081_ (.A1(\as1802.regs[2][10] ),
    .A2(_0870_),
    .B1(\as1802.regs[2][11] ),
    .Y(_0978_));
 sky130_fd_sc_hd__and3_1 _3082_ (.A(net130),
    .B(_0977_),
    .C(_0978_),
    .X(_0979_));
 sky130_fd_sc_hd__a21oi_2 _3083_ (.A1(_0975_),
    .A2(_0976_),
    .B1(_0979_),
    .Y(_0980_));
 sky130_fd_sc_hd__mux2_1 _3084_ (.A0(\as1802.regs[10][11] ),
    .A1(net46),
    .S(_0762_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _3085_ (.A0(\as1802.regs[13][12] ),
    .A1(\as1802.regs[12][12] ),
    .S(net106),
    .X(_0981_));
 sky130_fd_sc_hd__or2_1 _3086_ (.A(net124),
    .B(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__mux2_1 _3087_ (.A0(\as1802.regs[15][12] ),
    .A1(\as1802.regs[14][12] ),
    .S(net106),
    .X(_0983_));
 sky130_fd_sc_hd__o211a_2 _3088_ (.A1(net116),
    .A2(_0983_),
    .B1(_0982_),
    .C1(net91),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _3089_ (.A0(\as1802.regs[9][12] ),
    .A1(\as1802.regs[8][12] ),
    .S(net105),
    .X(_0985_));
 sky130_fd_sc_hd__and3_1 _3090_ (.A(\as1802.regs[11][12] ),
    .B(net153),
    .C(net145),
    .X(_0986_));
 sky130_fd_sc_hd__a211o_1 _3091_ (.A1(\as1802.regs[10][12] ),
    .A2(net105),
    .B1(_0986_),
    .C1(net116),
    .X(_0987_));
 sky130_fd_sc_hd__o211a_1 _3092_ (.A1(net124),
    .A2(_0985_),
    .B1(_0987_),
    .C1(net95),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_1 _3093_ (.A0(\as1802.regs[3][12] ),
    .A1(\as1802.regs[2][12] ),
    .S(net110),
    .X(_0989_));
 sky130_fd_sc_hd__mux2_1 _3094_ (.A0(\as1802.regs[1][12] ),
    .A1(\as1802.regs[0][12] ),
    .S(net110),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_1 _3095_ (.A0(_0989_),
    .A1(_0990_),
    .S(net116),
    .X(_0991_));
 sky130_fd_sc_hd__mux2_1 _3096_ (.A0(\as1802.regs[5][12] ),
    .A1(\as1802.regs[4][12] ),
    .S(net106),
    .X(_0992_));
 sky130_fd_sc_hd__and3_1 _3097_ (.A(\as1802.regs[7][12] ),
    .B(net153),
    .C(net145),
    .X(_0993_));
 sky130_fd_sc_hd__a211o_1 _3098_ (.A1(\as1802.regs[6][12] ),
    .A2(net106),
    .B1(_0993_),
    .C1(net116),
    .X(_0994_));
 sky130_fd_sc_hd__o211a_1 _3099_ (.A1(net124),
    .A2(_0992_),
    .B1(_0994_),
    .C1(net91),
    .X(_0995_));
 sky130_fd_sc_hd__a211o_1 _3100_ (.A1(net95),
    .A2(_0991_),
    .B1(_0995_),
    .C1(net86),
    .X(_0996_));
 sky130_fd_sc_hd__o31ai_4 _3101_ (.A1(net88),
    .A2(_0984_),
    .A3(_0988_),
    .B1(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__xnor2_1 _3102_ (.A(_0970_),
    .B(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__o21a_1 _3103_ (.A1(net165),
    .A2(_0998_),
    .B1(_2081_),
    .X(_0999_));
 sky130_fd_sc_hd__o21ai_1 _3104_ (.A1(net213),
    .A2(_2081_),
    .B1(net83),
    .Y(_1000_));
 sky130_fd_sc_hd__xnor2_1 _3105_ (.A(_0966_),
    .B(_0997_),
    .Y(_1001_));
 sky130_fd_sc_hd__and2b_1 _3106_ (.A_N(net264),
    .B(\as1802.regs[10][12] ),
    .X(_1002_));
 sky130_fd_sc_hd__a21bo_1 _3107_ (.A1(net264),
    .A2(\as1802.regs[11][12] ),
    .B1_N(net252),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _3108_ (.A0(\as1802.regs[8][12] ),
    .A1(\as1802.regs[9][12] ),
    .S(net264),
    .X(_1004_));
 sky130_fd_sc_hd__o221a_1 _3109_ (.A1(_1002_),
    .A2(_1003_),
    .B1(_1004_),
    .B2(net252),
    .C1(net199),
    .X(_1005_));
 sky130_fd_sc_hd__mux4_1 _3110_ (.A0(\as1802.regs[12][12] ),
    .A1(\as1802.regs[13][12] ),
    .A2(\as1802.regs[14][12] ),
    .A3(\as1802.regs[15][12] ),
    .S0(net264),
    .S1(net252),
    .X(_1006_));
 sky130_fd_sc_hd__a21o_1 _3111_ (.A1(net244),
    .A2(_1006_),
    .B1(net197),
    .X(_1007_));
 sky130_fd_sc_hd__mux4_1 _3112_ (.A0(\as1802.regs[0][12] ),
    .A1(\as1802.regs[1][12] ),
    .A2(\as1802.regs[2][12] ),
    .A3(\as1802.regs[3][12] ),
    .S0(net265),
    .S1(net255),
    .X(_1008_));
 sky130_fd_sc_hd__mux4_1 _3113_ (.A0(\as1802.regs[4][12] ),
    .A1(\as1802.regs[5][12] ),
    .A2(\as1802.regs[6][12] ),
    .A3(\as1802.regs[7][12] ),
    .S0(net265),
    .S1(net252),
    .X(_1009_));
 sky130_fd_sc_hd__mux2_1 _3114_ (.A0(_1008_),
    .A1(_1009_),
    .S(net244),
    .X(_1010_));
 sky130_fd_sc_hd__o22a_4 _3115_ (.A1(_1005_),
    .A2(_1007_),
    .B1(_1010_),
    .B2(net241),
    .X(_1011_));
 sky130_fd_sc_hd__o21a_1 _3116_ (.A1(_0938_),
    .A2(_1011_),
    .B1(_0803_),
    .X(_1012_));
 sky130_fd_sc_hd__nand2_1 _3117_ (.A(_0934_),
    .B(_1011_),
    .Y(_1013_));
 sky130_fd_sc_hd__or2_1 _3118_ (.A(_0913_),
    .B(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__or3_4 _3119_ (.A(_0860_),
    .B(_0909_),
    .C(_1013_),
    .X(_1015_));
 sky130_fd_sc_hd__o21ai_1 _3120_ (.A1(_0936_),
    .A2(_1011_),
    .B1(_1015_),
    .Y(_1016_));
 sky130_fd_sc_hd__a2bb2o_1 _3121_ (.A1_N(_0803_),
    .A2_N(_1016_),
    .B1(_1014_),
    .B2(_1012_),
    .X(_1017_));
 sky130_fd_sc_hd__a21o_1 _3122_ (.A1(net34),
    .A2(_2075_),
    .B1(_2148_),
    .X(_1018_));
 sky130_fd_sc_hd__a21o_1 _3123_ (.A1(_2077_),
    .A2(_1017_),
    .B1(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__nor2_1 _3124_ (.A(net200),
    .B(_1016_),
    .Y(_1020_));
 sky130_fd_sc_hd__a211o_1 _3125_ (.A1(net200),
    .A2(_1011_),
    .B1(_1020_),
    .C1(net126),
    .X(_1021_));
 sky130_fd_sc_hd__and3_1 _3126_ (.A(net80),
    .B(_1019_),
    .C(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__nor2_1 _3127_ (.A(net130),
    .B(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__o221a_1 _3128_ (.A1(_2101_),
    .A2(_0998_),
    .B1(_1001_),
    .B2(_0559_),
    .C1(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__o21a_1 _3129_ (.A1(_0999_),
    .A2(_1000_),
    .B1(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__or2_2 _3130_ (.A(\as1802.regs[2][12] ),
    .B(_0977_),
    .X(_1026_));
 sky130_fd_sc_hd__a21oi_1 _3131_ (.A1(\as1802.regs[2][12] ),
    .A2(_0977_),
    .B1(net128),
    .Y(_1027_));
 sky130_fd_sc_hd__a21oi_1 _3132_ (.A1(_1026_),
    .A2(_1027_),
    .B1(_1025_),
    .Y(_1028_));
 sky130_fd_sc_hd__mux2_1 _3133_ (.A0(\as1802.regs[10][12] ),
    .A1(net44),
    .S(_0762_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _3134_ (.A0(\as1802.regs[9][13] ),
    .A1(\as1802.regs[8][13] ),
    .S(net106),
    .X(_1029_));
 sky130_fd_sc_hd__and3_1 _3135_ (.A(\as1802.regs[11][13] ),
    .B(net153),
    .C(net145),
    .X(_1030_));
 sky130_fd_sc_hd__a211o_1 _3136_ (.A1(\as1802.regs[10][13] ),
    .A2(net110),
    .B1(_1030_),
    .C1(net117),
    .X(_1031_));
 sky130_fd_sc_hd__o211a_1 _3137_ (.A1(net124),
    .A2(_1029_),
    .B1(_1031_),
    .C1(net95),
    .X(_1032_));
 sky130_fd_sc_hd__mux2_1 _3138_ (.A0(\as1802.regs[15][13] ),
    .A1(\as1802.regs[14][13] ),
    .S(net106),
    .X(_1033_));
 sky130_fd_sc_hd__or2_1 _3139_ (.A(net116),
    .B(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__mux2_1 _3140_ (.A0(\as1802.regs[13][13] ),
    .A1(\as1802.regs[12][13] ),
    .S(net106),
    .X(_1035_));
 sky130_fd_sc_hd__o211a_1 _3141_ (.A1(net124),
    .A2(_1035_),
    .B1(_1034_),
    .C1(net91),
    .X(_1036_));
 sky130_fd_sc_hd__mux2_1 _3142_ (.A0(\as1802.regs[1][13] ),
    .A1(\as1802.regs[0][13] ),
    .S(net109),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _3143_ (.A0(\as1802.regs[3][13] ),
    .A1(\as1802.regs[2][13] ),
    .S(net109),
    .X(_1038_));
 sky130_fd_sc_hd__mux2_1 _3144_ (.A0(_1037_),
    .A1(_1038_),
    .S(net125),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _3145_ (.A0(\as1802.regs[5][13] ),
    .A1(\as1802.regs[4][13] ),
    .S(net109),
    .X(_1040_));
 sky130_fd_sc_hd__and3_1 _3146_ (.A(\as1802.regs[7][13] ),
    .B(net153),
    .C(net145),
    .X(_1041_));
 sky130_fd_sc_hd__a211o_1 _3147_ (.A1(\as1802.regs[6][13] ),
    .A2(net109),
    .B1(_1041_),
    .C1(net117),
    .X(_1042_));
 sky130_fd_sc_hd__o211a_1 _3148_ (.A1(net125),
    .A2(_1040_),
    .B1(_1042_),
    .C1(net92),
    .X(_1043_));
 sky130_fd_sc_hd__a211o_1 _3149_ (.A1(_2168_),
    .A2(_1039_),
    .B1(_1043_),
    .C1(net86),
    .X(_1044_));
 sky130_fd_sc_hd__o31ai_4 _3150_ (.A1(net88),
    .A2(_1032_),
    .A3(_1036_),
    .B1(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__and2_2 _3151_ (.A(_0997_),
    .B(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__nand3_2 _3152_ (.A(_0785_),
    .B(_0965_),
    .C(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__a31o_1 _3153_ (.A1(_0785_),
    .A2(_0965_),
    .A3(_0997_),
    .B1(_1045_),
    .X(_1048_));
 sky130_fd_sc_hd__a21oi_1 _3154_ (.A1(_1047_),
    .A2(_1048_),
    .B1(_0380_),
    .Y(_1049_));
 sky130_fd_sc_hd__o31a_1 _3155_ (.A1(_0718_),
    .A2(_0969_),
    .A3(_0997_),
    .B1(_1045_),
    .X(_1050_));
 sky130_fd_sc_hd__or2_1 _3156_ (.A(_0997_),
    .B(_1045_),
    .X(_1051_));
 sky130_fd_sc_hd__or3_2 _3157_ (.A(_0718_),
    .B(_0969_),
    .C(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__and2b_1 _3158_ (.A_N(_1050_),
    .B(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__a211o_1 _3159_ (.A1(_0380_),
    .A2(_1053_),
    .B1(_1049_),
    .C1(_2080_),
    .X(_1054_));
 sky130_fd_sc_hd__o211a_1 _3160_ (.A1(net212),
    .A2(_2081_),
    .B1(net83),
    .C1(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__and2b_1 _3161_ (.A_N(net265),
    .B(\as1802.regs[10][13] ),
    .X(_1056_));
 sky130_fd_sc_hd__a21bo_1 _3162_ (.A1(net267),
    .A2(\as1802.regs[11][13] ),
    .B1_N(net252),
    .X(_1057_));
 sky130_fd_sc_hd__mux2_1 _3163_ (.A0(\as1802.regs[8][13] ),
    .A1(\as1802.regs[9][13] ),
    .S(net265),
    .X(_1058_));
 sky130_fd_sc_hd__o221a_1 _3164_ (.A1(_1056_),
    .A2(_1057_),
    .B1(_1058_),
    .B2(net255),
    .C1(net199),
    .X(_1059_));
 sky130_fd_sc_hd__mux4_1 _3165_ (.A0(\as1802.regs[12][13] ),
    .A1(\as1802.regs[13][13] ),
    .A2(\as1802.regs[14][13] ),
    .A3(\as1802.regs[15][13] ),
    .S0(net265),
    .S1(net255),
    .X(_1060_));
 sky130_fd_sc_hd__a21o_1 _3166_ (.A1(net244),
    .A2(_1060_),
    .B1(_1932_),
    .X(_1061_));
 sky130_fd_sc_hd__mux4_1 _3167_ (.A0(\as1802.regs[0][13] ),
    .A1(\as1802.regs[1][13] ),
    .A2(\as1802.regs[2][13] ),
    .A3(\as1802.regs[3][13] ),
    .S0(net267),
    .S1(net254),
    .X(_1062_));
 sky130_fd_sc_hd__mux4_1 _3168_ (.A0(\as1802.regs[4][13] ),
    .A1(\as1802.regs[5][13] ),
    .A2(\as1802.regs[6][13] ),
    .A3(\as1802.regs[7][13] ),
    .S0(net267),
    .S1(net254),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_1 _3169_ (.A0(_1062_),
    .A1(_1063_),
    .S(_0002_),
    .X(_1064_));
 sky130_fd_sc_hd__o22a_2 _3170_ (.A1(_1059_),
    .A2(_1061_),
    .B1(_1064_),
    .B2(net241),
    .X(_1065_));
 sky130_fd_sc_hd__inv_2 _3171_ (.A(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__or2_4 _3172_ (.A(_1015_),
    .B(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__xnor2_2 _3173_ (.A(_1015_),
    .B(_1066_),
    .Y(_1068_));
 sky130_fd_sc_hd__and3_1 _3174_ (.A(_0803_),
    .B(_1014_),
    .C(_1066_),
    .X(_1069_));
 sky130_fd_sc_hd__nor2_1 _3175_ (.A(_1014_),
    .B(_1066_),
    .Y(_1070_));
 sky130_fd_sc_hd__or3_1 _3176_ (.A(_0913_),
    .B(_1013_),
    .C(_1066_),
    .X(_1071_));
 sky130_fd_sc_hd__a211oi_1 _3177_ (.A1(_0802_),
    .A2(_1068_),
    .B1(_1069_),
    .C1(_1070_),
    .Y(_1072_));
 sky130_fd_sc_hd__or2_1 _3178_ (.A(net35),
    .B(_2077_),
    .X(_1073_));
 sky130_fd_sc_hd__o211a_1 _3179_ (.A1(_2076_),
    .A2(_1072_),
    .B1(_1073_),
    .C1(net126),
    .X(_1074_));
 sky130_fd_sc_hd__nand2_1 _3180_ (.A(net227),
    .B(_1068_),
    .Y(_1075_));
 sky130_fd_sc_hd__o211a_1 _3181_ (.A1(net227),
    .A2(_1065_),
    .B1(_1075_),
    .C1(_2148_),
    .X(_1076_));
 sky130_fd_sc_hd__or3_1 _3182_ (.A(net132),
    .B(_1074_),
    .C(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__nand2_1 _3183_ (.A(net132),
    .B(_1068_),
    .Y(_1078_));
 sky130_fd_sc_hd__a31o_1 _3184_ (.A1(net80),
    .A2(_1077_),
    .A3(_1078_),
    .B1(net130),
    .X(_1079_));
 sky130_fd_sc_hd__nand3_1 _3185_ (.A(_2096_),
    .B(_1047_),
    .C(_1048_),
    .Y(_1080_));
 sky130_fd_sc_hd__o211a_1 _3186_ (.A1(_2096_),
    .A2(_1053_),
    .B1(_1080_),
    .C1(_2107_),
    .X(_1081_));
 sky130_fd_sc_hd__a21oi_1 _3187_ (.A1(\as1802.regs[2][13] ),
    .A2(_1026_),
    .B1(net128),
    .Y(_1082_));
 sky130_fd_sc_hd__o21ai_1 _3188_ (.A1(\as1802.regs[2][13] ),
    .A2(_1026_),
    .B1(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__o31a_2 _3189_ (.A1(_1055_),
    .A2(_1079_),
    .A3(_1081_),
    .B1(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__mux2_1 _3190_ (.A0(\as1802.regs[10][13] ),
    .A1(net42),
    .S(_0762_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _3191_ (.A0(\as1802.regs[9][14] ),
    .A1(\as1802.regs[8][14] ),
    .S(net108),
    .X(_1085_));
 sky130_fd_sc_hd__and3_1 _3192_ (.A(\as1802.regs[11][14] ),
    .B(net153),
    .C(net145),
    .X(_1086_));
 sky130_fd_sc_hd__a211o_1 _3193_ (.A1(\as1802.regs[10][14] ),
    .A2(net107),
    .B1(_1086_),
    .C1(net117),
    .X(_1087_));
 sky130_fd_sc_hd__o211a_1 _3194_ (.A1(net123),
    .A2(_1085_),
    .B1(_1087_),
    .C1(net95),
    .X(_1088_));
 sky130_fd_sc_hd__mux2_1 _3195_ (.A0(\as1802.regs[15][14] ),
    .A1(\as1802.regs[14][14] ),
    .S(net107),
    .X(_1089_));
 sky130_fd_sc_hd__or2_1 _3196_ (.A(net117),
    .B(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__mux2_1 _3197_ (.A0(\as1802.regs[13][14] ),
    .A1(\as1802.regs[12][14] ),
    .S(net107),
    .X(_1091_));
 sky130_fd_sc_hd__or2_1 _3198_ (.A(net123),
    .B(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__a31o_1 _3199_ (.A1(net91),
    .A2(_1090_),
    .A3(_1092_),
    .B1(net88),
    .X(_1093_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(\as1802.regs[3][14] ),
    .A1(\as1802.regs[2][14] ),
    .S(net110),
    .X(_1094_));
 sky130_fd_sc_hd__mux2_1 _3201_ (.A0(\as1802.regs[1][14] ),
    .A1(\as1802.regs[0][14] ),
    .S(net110),
    .X(_1095_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(_1094_),
    .A1(_1095_),
    .S(net117),
    .X(_1096_));
 sky130_fd_sc_hd__mux2_1 _3203_ (.A0(\as1802.regs[5][14] ),
    .A1(\as1802.regs[4][14] ),
    .S(net108),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_1 _3204_ (.A0(\as1802.regs[7][14] ),
    .A1(\as1802.regs[6][14] ),
    .S(net108),
    .X(_1098_));
 sky130_fd_sc_hd__mux2_1 _3205_ (.A0(_1097_),
    .A1(_1098_),
    .S(net123),
    .X(_1099_));
 sky130_fd_sc_hd__mux2_1 _3206_ (.A0(_1096_),
    .A1(_1099_),
    .S(net92),
    .X(_1100_));
 sky130_fd_sc_hd__o22a_4 _3207_ (.A1(_1088_),
    .A2(_1093_),
    .B1(_1100_),
    .B2(net86),
    .X(_1101_));
 sky130_fd_sc_hd__inv_2 _3208_ (.A(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__or4_1 _3209_ (.A(_0718_),
    .B(_0969_),
    .C(_1051_),
    .D(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__xnor2_1 _3210_ (.A(_1052_),
    .B(_1101_),
    .Y(_1104_));
 sky130_fd_sc_hd__nand2_1 _3211_ (.A(_0380_),
    .B(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__xnor2_1 _3212_ (.A(_1047_),
    .B(_1101_),
    .Y(_1106_));
 sky130_fd_sc_hd__mux4_1 _3213_ (.A0(\as1802.regs[12][14] ),
    .A1(\as1802.regs[13][14] ),
    .A2(\as1802.regs[14][14] ),
    .A3(\as1802.regs[15][14] ),
    .S0(net266),
    .S1(net253),
    .X(_1107_));
 sky130_fd_sc_hd__and2b_1 _3214_ (.A_N(net266),
    .B(\as1802.regs[10][14] ),
    .X(_1108_));
 sky130_fd_sc_hd__a21bo_1 _3215_ (.A1(net266),
    .A2(\as1802.regs[11][14] ),
    .B1_N(net253),
    .X(_1109_));
 sky130_fd_sc_hd__mux2_1 _3216_ (.A0(\as1802.regs[8][14] ),
    .A1(\as1802.regs[9][14] ),
    .S(net266),
    .X(_1110_));
 sky130_fd_sc_hd__o221a_1 _3217_ (.A1(_1108_),
    .A2(_1109_),
    .B1(_1110_),
    .B2(net253),
    .C1(net199),
    .X(_1111_));
 sky130_fd_sc_hd__a211o_2 _3218_ (.A1(net244),
    .A2(_1107_),
    .B1(_1111_),
    .C1(_1932_),
    .X(_1112_));
 sky130_fd_sc_hd__mux4_1 _3219_ (.A0(\as1802.regs[4][14] ),
    .A1(\as1802.regs[5][14] ),
    .A2(\as1802.regs[6][14] ),
    .A3(\as1802.regs[7][14] ),
    .S0(net267),
    .S1(net253),
    .X(_1113_));
 sky130_fd_sc_hd__mux4_1 _3220_ (.A0(\as1802.regs[0][14] ),
    .A1(\as1802.regs[1][14] ),
    .A2(\as1802.regs[2][14] ),
    .A3(\as1802.regs[3][14] ),
    .S0(net267),
    .S1(net254),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_2 _3221_ (.A0(_1113_),
    .A1(_1114_),
    .S(_1931_),
    .X(_1115_));
 sky130_fd_sc_hd__o21ai_4 _3222_ (.A1(net241),
    .A2(_1115_),
    .B1(_1112_),
    .Y(_1116_));
 sky130_fd_sc_hd__xor2_1 _3223_ (.A(_1071_),
    .B(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__nor2_1 _3224_ (.A(net227),
    .B(_1116_),
    .Y(_1118_));
 sky130_fd_sc_hd__a21oi_1 _3225_ (.A1(net165),
    .A2(_1106_),
    .B1(_2080_),
    .Y(_1119_));
 sky130_fd_sc_hd__a221o_1 _3226_ (.A1(_1929_),
    .A2(_2080_),
    .B1(_1105_),
    .B2(_1119_),
    .C1(_2089_),
    .X(_1120_));
 sky130_fd_sc_hd__nor2_1 _3227_ (.A(_2097_),
    .B(_1106_),
    .Y(_1121_));
 sky130_fd_sc_hd__o21ai_1 _3228_ (.A1(_2096_),
    .A2(_1104_),
    .B1(_2107_),
    .Y(_1122_));
 sky130_fd_sc_hd__xor2_4 _3229_ (.A(_1067_),
    .B(_1116_),
    .X(_1123_));
 sky130_fd_sc_hd__nor2_1 _3230_ (.A(_2058_),
    .B(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__mux2_1 _3231_ (.A0(_1117_),
    .A1(_1123_),
    .S(_0802_),
    .X(_1125_));
 sky130_fd_sc_hd__mux2_1 _3232_ (.A0(net205),
    .A1(_1125_),
    .S(_2077_),
    .X(_1126_));
 sky130_fd_sc_hd__a211o_1 _3233_ (.A1(net227),
    .A2(_1123_),
    .B1(_1118_),
    .C1(net126),
    .X(_1127_));
 sky130_fd_sc_hd__o21a_1 _3234_ (.A1(_2148_),
    .A2(_1126_),
    .B1(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__o21ai_1 _3235_ (.A1(net132),
    .A2(_1128_),
    .B1(net80),
    .Y(_1129_));
 sky130_fd_sc_hd__o221a_1 _3236_ (.A1(_1121_),
    .A2(_1122_),
    .B1(_1124_),
    .B2(_1129_),
    .C1(net128),
    .X(_1130_));
 sky130_fd_sc_hd__or3_2 _3237_ (.A(\as1802.regs[2][13] ),
    .B(\as1802.regs[2][14] ),
    .C(_1026_),
    .X(_1131_));
 sky130_fd_sc_hd__o21ai_1 _3238_ (.A1(\as1802.regs[2][13] ),
    .A2(_1026_),
    .B1(\as1802.regs[2][14] ),
    .Y(_1132_));
 sky130_fd_sc_hd__and3_1 _3239_ (.A(net130),
    .B(_1131_),
    .C(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__a21oi_2 _3240_ (.A1(_1120_),
    .A2(_1130_),
    .B1(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__mux2_1 _3241_ (.A0(\as1802.regs[10][14] ),
    .A1(net40),
    .S(_0762_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _3242_ (.A0(\as1802.regs[9][15] ),
    .A1(\as1802.regs[8][15] ),
    .S(net107),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _3243_ (.A0(\as1802.regs[11][15] ),
    .A1(\as1802.regs[10][15] ),
    .S(net107),
    .X(_1136_));
 sky130_fd_sc_hd__mux2_1 _3244_ (.A0(_1135_),
    .A1(_1136_),
    .S(net123),
    .X(_1137_));
 sky130_fd_sc_hd__mux2_1 _3245_ (.A0(\as1802.regs[15][15] ),
    .A1(\as1802.regs[14][15] ),
    .S(net107),
    .X(_1138_));
 sky130_fd_sc_hd__or2_1 _3246_ (.A(net117),
    .B(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__mux2_1 _3247_ (.A0(\as1802.regs[13][15] ),
    .A1(\as1802.regs[12][15] ),
    .S(net107),
    .X(_1140_));
 sky130_fd_sc_hd__o21a_1 _3248_ (.A1(net123),
    .A2(_1140_),
    .B1(net91),
    .X(_1141_));
 sky130_fd_sc_hd__a221o_1 _3249_ (.A1(_2168_),
    .A2(_1137_),
    .B1(_1139_),
    .B2(_1141_),
    .C1(net88),
    .X(_1142_));
 sky130_fd_sc_hd__mux2_1 _3250_ (.A0(\as1802.regs[3][15] ),
    .A1(\as1802.regs[2][15] ),
    .S(net111),
    .X(_1143_));
 sky130_fd_sc_hd__mux2_1 _3251_ (.A0(\as1802.regs[1][15] ),
    .A1(\as1802.regs[0][15] ),
    .S(net111),
    .X(_1144_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(_1143_),
    .A1(_1144_),
    .S(net117),
    .X(_1145_));
 sky130_fd_sc_hd__mux2_1 _3253_ (.A0(\as1802.regs[5][15] ),
    .A1(\as1802.regs[4][15] ),
    .S(net109),
    .X(_1146_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(\as1802.regs[7][15] ),
    .A1(\as1802.regs[6][15] ),
    .S(net109),
    .X(_1147_));
 sky130_fd_sc_hd__mux2_1 _3255_ (.A0(_1146_),
    .A1(_1147_),
    .S(net123),
    .X(_1148_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(_1145_),
    .A1(_1148_),
    .S(net92),
    .X(_1149_));
 sky130_fd_sc_hd__o21a_4 _3257_ (.A1(net86),
    .A2(_1149_),
    .B1(_1142_),
    .X(_1150_));
 sky130_fd_sc_hd__inv_2 _3258_ (.A(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__nor2_1 _3259_ (.A(net211),
    .B(_2081_),
    .Y(_1152_));
 sky130_fd_sc_hd__mux4_1 _3260_ (.A0(\as1802.regs[12][15] ),
    .A1(\as1802.regs[13][15] ),
    .A2(\as1802.regs[14][15] ),
    .A3(\as1802.regs[15][15] ),
    .S0(net266),
    .S1(net253),
    .X(_1153_));
 sky130_fd_sc_hd__nand2_1 _3261_ (.A(net244),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__mux2_1 _3262_ (.A0(\as1802.regs[10][15] ),
    .A1(\as1802.regs[11][15] ),
    .S(net267),
    .X(_1155_));
 sky130_fd_sc_hd__inv_2 _3263_ (.A(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__mux2_1 _3264_ (.A0(\as1802.regs[8][15] ),
    .A1(\as1802.regs[9][15] ),
    .S(net267),
    .X(_1157_));
 sky130_fd_sc_hd__nor2_1 _3265_ (.A(net254),
    .B(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hd__a211o_1 _3266_ (.A1(net253),
    .A2(_1156_),
    .B1(_1158_),
    .C1(net244),
    .X(_1159_));
 sky130_fd_sc_hd__mux4_1 _3267_ (.A0(\as1802.regs[4][15] ),
    .A1(\as1802.regs[5][15] ),
    .A2(\as1802.regs[6][15] ),
    .A3(\as1802.regs[7][15] ),
    .S0(net267),
    .S1(net254),
    .X(_1160_));
 sky130_fd_sc_hd__mux4_2 _3268_ (.A0(\as1802.regs[0][15] ),
    .A1(\as1802.regs[1][15] ),
    .A2(\as1802.regs[2][15] ),
    .A3(\as1802.regs[3][15] ),
    .S0(_0000_),
    .S1(net254),
    .X(_1161_));
 sky130_fd_sc_hd__mux2_1 _3269_ (.A0(_1160_),
    .A1(_1161_),
    .S(_1931_),
    .X(_1162_));
 sky130_fd_sc_hd__nor2_1 _3270_ (.A(net241),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__a31o_4 _3271_ (.A1(net241),
    .A2(_1154_),
    .A3(_1159_),
    .B1(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__inv_2 _3272_ (.A(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__or4_2 _3273_ (.A(_0911_),
    .B(_1013_),
    .C(_1066_),
    .D(_1116_),
    .X(_1166_));
 sky130_fd_sc_hd__xnor2_2 _3274_ (.A(_1164_),
    .B(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__mux2_1 _3275_ (.A0(_1164_),
    .A1(_1167_),
    .S(net155),
    .X(_1168_));
 sky130_fd_sc_hd__or3_1 _3276_ (.A(\as1802.cond_inv ),
    .B(_2056_),
    .C(_1164_),
    .X(_1169_));
 sky130_fd_sc_hd__o221a_1 _3277_ (.A1(_2049_),
    .A2(_1167_),
    .B1(_1168_),
    .B2(_0803_),
    .C1(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__nor2_1 _3278_ (.A(_2076_),
    .B(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__a211o_1 _3279_ (.A1(net37),
    .A2(_2076_),
    .B1(_2150_),
    .C1(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__a21oi_1 _3280_ (.A1(_2141_),
    .A2(_1165_),
    .B1(net126),
    .Y(_1173_));
 sky130_fd_sc_hd__o21ai_1 _3281_ (.A1(_2141_),
    .A2(_1167_),
    .B1(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__nand3_1 _3282_ (.A(net80),
    .B(_1172_),
    .C(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__nand2_1 _3283_ (.A(_1101_),
    .B(_1150_),
    .Y(_1176_));
 sky130_fd_sc_hd__a2bb2o_1 _3284_ (.A1_N(_1052_),
    .A2_N(_1176_),
    .B1(_1151_),
    .B2(_1103_),
    .X(_1177_));
 sky130_fd_sc_hd__a41oi_4 _3285_ (.A1(_0785_),
    .A2(_0965_),
    .A3(_1046_),
    .A4(_1102_),
    .B1(_1150_),
    .Y(_1178_));
 sky130_fd_sc_hd__and2b_1 _3286_ (.A_N(_1101_),
    .B(_1150_),
    .X(_1179_));
 sky130_fd_sc_hd__and4_1 _3287_ (.A(_0785_),
    .B(_0965_),
    .C(_1046_),
    .D(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__or3_1 _3288_ (.A(_0380_),
    .B(_1178_),
    .C(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__o211a_1 _3289_ (.A1(net165),
    .A2(_1177_),
    .B1(_1181_),
    .C1(_2081_),
    .X(_1182_));
 sky130_fd_sc_hd__and2_1 _3290_ (.A(_2097_),
    .B(_1177_),
    .X(_1183_));
 sky130_fd_sc_hd__o31a_1 _3291_ (.A1(_2089_),
    .A2(_1152_),
    .A3(_1182_),
    .B1(_1175_),
    .X(_1184_));
 sky130_fd_sc_hd__o21a_1 _3292_ (.A1(_1178_),
    .A2(_1180_),
    .B1(_2109_),
    .X(_1185_));
 sky130_fd_sc_hd__o31a_2 _3293_ (.A1(_2110_),
    .A2(_1183_),
    .A3(_1185_),
    .B1(net128),
    .X(_1186_));
 sky130_fd_sc_hd__a21oi_1 _3294_ (.A1(\as1802.regs[2][15] ),
    .A2(_1131_),
    .B1(net128),
    .Y(_1187_));
 sky130_fd_sc_hd__o21a_1 _3295_ (.A1(\as1802.regs[2][15] ),
    .A2(_1131_),
    .B1(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__a21oi_4 _3296_ (.A1(_1184_),
    .A2(_1186_),
    .B1(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__mux2_1 _3297_ (.A0(\as1802.regs[10][15] ),
    .A1(net39),
    .S(_0762_),
    .X(_0027_));
 sky130_fd_sc_hd__nor2_8 _3298_ (.A(_2112_),
    .B(_2115_),
    .Y(_1190_));
 sky130_fd_sc_hd__nor2_4 _3299_ (.A(_2119_),
    .B(_2122_),
    .Y(_1191_));
 sky130_fd_sc_hd__and3_4 _3300_ (.A(net71),
    .B(_1190_),
    .C(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__mux2_1 _3301_ (.A0(\as1802.regs[0][8] ),
    .A1(net53),
    .S(_1192_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _3302_ (.A0(\as1802.regs[0][9] ),
    .A1(net51),
    .S(_1192_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _3303_ (.A0(\as1802.regs[0][10] ),
    .A1(net49),
    .S(_1192_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _3304_ (.A0(\as1802.regs[0][11] ),
    .A1(net47),
    .S(_1192_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _3305_ (.A0(\as1802.regs[0][12] ),
    .A1(net45),
    .S(_1192_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _3306_ (.A0(\as1802.regs[0][13] ),
    .A1(net43),
    .S(_1192_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _3307_ (.A0(\as1802.regs[0][14] ),
    .A1(net41),
    .S(_1192_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _3308_ (.A0(\as1802.regs[0][15] ),
    .A1(net38),
    .S(_1192_),
    .X(_0035_));
 sky130_fd_sc_hd__and3_4 _3309_ (.A(_0759_),
    .B(net70),
    .C(_1190_),
    .X(_1193_));
 sky130_fd_sc_hd__mux2_1 _3310_ (.A0(\as1802.regs[8][8] ),
    .A1(net52),
    .S(_1193_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _3311_ (.A0(\as1802.regs[8][9] ),
    .A1(net50),
    .S(_1193_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _3312_ (.A0(\as1802.regs[8][10] ),
    .A1(net48),
    .S(_1193_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _3313_ (.A0(\as1802.regs[8][11] ),
    .A1(net46),
    .S(_1193_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _3314_ (.A0(\as1802.regs[8][12] ),
    .A1(net44),
    .S(_1193_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _3315_ (.A0(\as1802.regs[8][13] ),
    .A1(net42),
    .S(_1193_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _3316_ (.A0(\as1802.regs[8][14] ),
    .A1(net40),
    .S(_1193_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _3317_ (.A0(\as1802.regs[8][15] ),
    .A1(net38),
    .S(_1193_),
    .X(_0043_));
 sky130_fd_sc_hd__nor2_4 _3318_ (.A(_2119_),
    .B(_2123_),
    .Y(_1194_));
 sky130_fd_sc_hd__and3_4 _3319_ (.A(net70),
    .B(_1190_),
    .C(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__mux2_1 _3320_ (.A0(\as1802.regs[4][8] ),
    .A1(net52),
    .S(_1195_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _3321_ (.A0(\as1802.regs[4][9] ),
    .A1(net50),
    .S(_1195_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _3322_ (.A0(\as1802.regs[4][10] ),
    .A1(net48),
    .S(_1195_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _3323_ (.A0(\as1802.regs[4][11] ),
    .A1(net46),
    .S(_1195_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _3324_ (.A0(\as1802.regs[4][12] ),
    .A1(net44),
    .S(_1195_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _3325_ (.A0(\as1802.regs[4][13] ),
    .A1(net42),
    .S(_1195_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _3326_ (.A0(\as1802.regs[4][14] ),
    .A1(net40),
    .S(_1195_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _3327_ (.A0(\as1802.regs[4][15] ),
    .A1(net39),
    .S(_1195_),
    .X(_0051_));
 sky130_fd_sc_hd__nor2_8 _3328_ (.A(_2112_),
    .B(_2116_),
    .Y(_1196_));
 sky130_fd_sc_hd__and3_4 _3329_ (.A(net70),
    .B(_1194_),
    .C(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__mux2_1 _3330_ (.A0(\as1802.regs[5][8] ),
    .A1(net53),
    .S(_1197_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _3331_ (.A0(\as1802.regs[5][9] ),
    .A1(net50),
    .S(_1197_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _3332_ (.A0(\as1802.regs[5][10] ),
    .A1(net48),
    .S(_1197_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _3333_ (.A0(\as1802.regs[5][11] ),
    .A1(net46),
    .S(_1197_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _3334_ (.A0(\as1802.regs[5][12] ),
    .A1(net44),
    .S(_1197_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _3335_ (.A0(\as1802.regs[5][13] ),
    .A1(net42),
    .S(_1197_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _3336_ (.A0(\as1802.regs[5][14] ),
    .A1(net41),
    .S(_1197_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _3337_ (.A0(\as1802.regs[5][15] ),
    .A1(net39),
    .S(_1197_),
    .X(_0059_));
 sky130_fd_sc_hd__and3_4 _3338_ (.A(_2117_),
    .B(net71),
    .C(_1194_),
    .X(_1198_));
 sky130_fd_sc_hd__mux2_1 _3339_ (.A0(\as1802.regs[7][8] ),
    .A1(net53),
    .S(_1198_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _3340_ (.A0(\as1802.regs[7][9] ),
    .A1(net51),
    .S(_1198_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _3341_ (.A0(\as1802.regs[7][10] ),
    .A1(net48),
    .S(_1198_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _3342_ (.A0(\as1802.regs[7][11] ),
    .A1(net47),
    .S(_1198_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _3343_ (.A0(\as1802.regs[7][12] ),
    .A1(net44),
    .S(_1198_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _3344_ (.A0(\as1802.regs[7][13] ),
    .A1(net43),
    .S(_1198_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _3345_ (.A0(\as1802.regs[7][14] ),
    .A1(net41),
    .S(_1198_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _3346_ (.A0(\as1802.regs[7][15] ),
    .A1(net39),
    .S(_1198_),
    .X(_0067_));
 sky130_fd_sc_hd__and3_4 _3347_ (.A(_0758_),
    .B(net70),
    .C(_1194_),
    .X(_1199_));
 sky130_fd_sc_hd__mux2_1 _3348_ (.A0(\as1802.regs[6][8] ),
    .A1(net53),
    .S(_1199_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _3349_ (.A0(\as1802.regs[6][9] ),
    .A1(net50),
    .S(_1199_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _3350_ (.A0(\as1802.regs[6][10] ),
    .A1(net48),
    .S(_1199_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _3351_ (.A0(\as1802.regs[6][11] ),
    .A1(net47),
    .S(_1199_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _3352_ (.A0(\as1802.regs[6][12] ),
    .A1(net45),
    .S(_1199_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _3353_ (.A0(\as1802.regs[6][13] ),
    .A1(net42),
    .S(_1199_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _3354_ (.A0(\as1802.regs[6][14] ),
    .A1(net40),
    .S(_1199_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _3355_ (.A0(\as1802.regs[6][15] ),
    .A1(net39),
    .S(_1199_),
    .X(_0075_));
 sky130_fd_sc_hd__and3_4 _3356_ (.A(_2117_),
    .B(net71),
    .C(_1191_),
    .X(_1200_));
 sky130_fd_sc_hd__mux2_1 _3357_ (.A0(\as1802.regs[3][8] ),
    .A1(net53),
    .S(_1200_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _3358_ (.A0(\as1802.regs[3][9] ),
    .A1(net51),
    .S(_1200_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _3359_ (.A0(\as1802.regs[3][10] ),
    .A1(net49),
    .S(_1200_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _3360_ (.A0(\as1802.regs[3][11] ),
    .A1(net47),
    .S(_1200_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _3361_ (.A0(\as1802.regs[3][12] ),
    .A1(net45),
    .S(_1200_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _3362_ (.A0(\as1802.regs[3][13] ),
    .A1(net43),
    .S(_1200_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _3363_ (.A0(\as1802.regs[3][14] ),
    .A1(net41),
    .S(_1200_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _3364_ (.A0(\as1802.regs[3][15] ),
    .A1(net38),
    .S(_1200_),
    .X(_0083_));
 sky130_fd_sc_hd__and3_4 _3365_ (.A(net72),
    .B(_0759_),
    .C(_1196_),
    .X(_1201_));
 sky130_fd_sc_hd__mux2_1 _3366_ (.A0(\as1802.regs[9][0] ),
    .A1(net68),
    .S(_1201_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _3367_ (.A0(\as1802.regs[9][1] ),
    .A1(net66),
    .S(_1201_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _3368_ (.A0(\as1802.regs[9][2] ),
    .A1(net64),
    .S(_1201_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _3369_ (.A0(\as1802.regs[9][3] ),
    .A1(net62),
    .S(_1201_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _3370_ (.A0(\as1802.regs[9][4] ),
    .A1(net60),
    .S(_1201_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _3371_ (.A0(\as1802.regs[9][5] ),
    .A1(net58),
    .S(_1201_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _3372_ (.A0(\as1802.regs[9][6] ),
    .A1(net56),
    .S(_1201_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _3373_ (.A0(\as1802.regs[9][7] ),
    .A1(net54),
    .S(_1201_),
    .X(_0091_));
 sky130_fd_sc_hd__and3_4 _3374_ (.A(net72),
    .B(_0759_),
    .C(_1190_),
    .X(_1202_));
 sky130_fd_sc_hd__mux2_1 _3375_ (.A0(\as1802.regs[8][0] ),
    .A1(net68),
    .S(_1202_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _3376_ (.A0(\as1802.regs[8][1] ),
    .A1(net66),
    .S(_1202_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _3377_ (.A0(\as1802.regs[8][2] ),
    .A1(net64),
    .S(_1202_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _3378_ (.A0(\as1802.regs[8][3] ),
    .A1(net62),
    .S(_1202_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _3379_ (.A0(\as1802.regs[8][4] ),
    .A1(net60),
    .S(_1202_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _3380_ (.A0(\as1802.regs[8][5] ),
    .A1(net58),
    .S(_1202_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _3381_ (.A0(\as1802.regs[8][6] ),
    .A1(net56),
    .S(_1202_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _3382_ (.A0(\as1802.regs[8][7] ),
    .A1(net54),
    .S(_1202_),
    .X(_0099_));
 sky130_fd_sc_hd__nand2_2 _3383_ (.A(\as1802.will_interrupt ),
    .B(net273),
    .Y(_1203_));
 sky130_fd_sc_hd__nor2_2 _3384_ (.A(net270),
    .B(_1993_),
    .Y(_1204_));
 sky130_fd_sc_hd__nand2_2 _3385_ (.A(net203),
    .B(_1994_),
    .Y(_1205_));
 sky130_fd_sc_hd__o21a_1 _3386_ (.A1(_1942_),
    .A2(net159),
    .B1(_1203_),
    .X(_1206_));
 sky130_fd_sc_hd__or2_4 _3387_ (.A(_1940_),
    .B(_1967_),
    .X(_1207_));
 sky130_fd_sc_hd__and3b_1 _3388_ (.A_N(_1940_),
    .B(net203),
    .C(_1936_),
    .X(_1208_));
 sky130_fd_sc_hd__o31a_1 _3389_ (.A1(net272),
    .A2(net220),
    .A3(_1940_),
    .B1(net195),
    .X(_1209_));
 sky130_fd_sc_hd__nand2_2 _3390_ (.A(_2020_),
    .B(_2053_),
    .Y(_1210_));
 sky130_fd_sc_hd__nor2_1 _3391_ (.A(net272),
    .B(_0378_),
    .Y(_1211_));
 sky130_fd_sc_hd__a31oi_4 _3392_ (.A1(net187),
    .A2(_2036_),
    .A3(_0378_),
    .B1(net271),
    .Y(_1212_));
 sky130_fd_sc_hd__nor2_1 _3393_ (.A(\as1802.IE ),
    .B(_1203_),
    .Y(_1213_));
 sky130_fd_sc_hd__o31a_1 _3394_ (.A1(net272),
    .A2(_1923_),
    .A3(_2018_),
    .B1(_2043_),
    .X(_1214_));
 sky130_fd_sc_hd__or3b_1 _3395_ (.A(_1206_),
    .B(_1213_),
    .C_N(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__nand2_1 _3396_ (.A(_1209_),
    .B(_1210_),
    .Y(_1216_));
 sky130_fd_sc_hd__nor3_2 _3397_ (.A(_1212_),
    .B(_1215_),
    .C(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__or2_1 _3398_ (.A(_1940_),
    .B(_1949_),
    .X(_1218_));
 sky130_fd_sc_hd__and2_2 _3399_ (.A(net203),
    .B(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__o211ai_4 _3400_ (.A1(_1938_),
    .A2(_2018_),
    .B1(_1219_),
    .C1(net190),
    .Y(_1220_));
 sky130_fd_sc_hd__nor2_4 _3401_ (.A(net274),
    .B(_2022_),
    .Y(_1221_));
 sky130_fd_sc_hd__o21ai_4 _3402_ (.A1(net235),
    .A2(_2004_),
    .B1(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__o311a_4 _3403_ (.A1(net274),
    .A2(_1923_),
    .A3(_1949_),
    .B1(_1217_),
    .C1(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__mux2_1 _3404_ (.A0(net237),
    .A1(net209),
    .S(net175),
    .X(_1224_));
 sky130_fd_sc_hd__or3b_1 _3405_ (.A(net275),
    .B(_1224_),
    .C_N(_1223_),
    .X(_1225_));
 sky130_fd_sc_hd__o211a_1 _3406_ (.A1(\as1802.P[0] ),
    .A2(_1223_),
    .B1(_1225_),
    .C1(net276),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_1 _3407_ (.A(net236),
    .B(net171),
    .Y(_1226_));
 sky130_fd_sc_hd__o2bb2a_2 _3408_ (.A1_N(net208),
    .A2_N(_2053_),
    .B1(_1226_),
    .B2(net275),
    .X(_1227_));
 sky130_fd_sc_hd__a21oi_4 _3409_ (.A1(_1223_),
    .A2(_1227_),
    .B1(net281),
    .Y(_1228_));
 sky130_fd_sc_hd__o21a_1 _3410_ (.A1(\as1802.P[1] ),
    .A2(_1223_),
    .B1(_1228_),
    .X(_0101_));
 sky130_fd_sc_hd__a21oi_1 _3411_ (.A1(net202),
    .A2(net170),
    .B1(net275),
    .Y(_1229_));
 sky130_fd_sc_hd__o21a_1 _3412_ (.A1(net206),
    .A2(net170),
    .B1(_1229_),
    .X(_1230_));
 sky130_fd_sc_hd__mux2_1 _3413_ (.A0(\as1802.P[2] ),
    .A1(_1230_),
    .S(_1223_),
    .X(_1231_));
 sky130_fd_sc_hd__and2_1 _3414_ (.A(net277),
    .B(_1231_),
    .X(_0102_));
 sky130_fd_sc_hd__a21oi_1 _3415_ (.A1(net201),
    .A2(net170),
    .B1(net275),
    .Y(_1232_));
 sky130_fd_sc_hd__o21a_1 _3416_ (.A1(net33),
    .A2(net170),
    .B1(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__mux2_1 _3417_ (.A0(\as1802.P[3] ),
    .A1(_1233_),
    .S(_1223_),
    .X(_1234_));
 sky130_fd_sc_hd__and2_1 _3418_ (.A(net277),
    .B(_1234_),
    .X(_0103_));
 sky130_fd_sc_hd__and3_4 _3419_ (.A(_2117_),
    .B(net72),
    .C(_1194_),
    .X(_1235_));
 sky130_fd_sc_hd__mux2_1 _3420_ (.A0(\as1802.regs[7][0] ),
    .A1(net69),
    .S(_1235_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _3421_ (.A0(\as1802.regs[7][1] ),
    .A1(net66),
    .S(_1235_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _3422_ (.A0(\as1802.regs[7][2] ),
    .A1(net65),
    .S(_1235_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _3423_ (.A0(\as1802.regs[7][3] ),
    .A1(net62),
    .S(_1235_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _3424_ (.A0(\as1802.regs[7][4] ),
    .A1(net60),
    .S(_1235_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _3425_ (.A0(\as1802.regs[7][5] ),
    .A1(net58),
    .S(_1235_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _3426_ (.A0(\as1802.regs[7][6] ),
    .A1(net56),
    .S(_1235_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _3427_ (.A0(\as1802.regs[7][7] ),
    .A1(net54),
    .S(_1235_),
    .X(_0111_));
 sky130_fd_sc_hd__and3_4 _3428_ (.A(net72),
    .B(_0758_),
    .C(_1194_),
    .X(_1236_));
 sky130_fd_sc_hd__mux2_1 _3429_ (.A0(\as1802.regs[6][0] ),
    .A1(net69),
    .S(_1236_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _3430_ (.A0(\as1802.regs[6][1] ),
    .A1(net66),
    .S(_1236_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _3431_ (.A0(\as1802.regs[6][2] ),
    .A1(net65),
    .S(_1236_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _3432_ (.A0(\as1802.regs[6][3] ),
    .A1(net62),
    .S(_1236_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _3433_ (.A0(\as1802.regs[6][4] ),
    .A1(net61),
    .S(_1236_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _3434_ (.A0(\as1802.regs[6][5] ),
    .A1(net58),
    .S(_1236_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _3435_ (.A0(\as1802.regs[6][6] ),
    .A1(net56),
    .S(_1236_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _3436_ (.A0(\as1802.regs[6][7] ),
    .A1(net54),
    .S(_1236_),
    .X(_0119_));
 sky130_fd_sc_hd__and3_4 _3437_ (.A(net73),
    .B(_1194_),
    .C(_1196_),
    .X(_1237_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(\as1802.regs[5][0] ),
    .A1(net69),
    .S(_1237_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _3439_ (.A0(\as1802.regs[5][1] ),
    .A1(net67),
    .S(_1237_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _3440_ (.A0(\as1802.regs[5][2] ),
    .A1(net65),
    .S(_1237_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _3441_ (.A0(\as1802.regs[5][3] ),
    .A1(net63),
    .S(_1237_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _3442_ (.A0(\as1802.regs[5][4] ),
    .A1(net61),
    .S(_1237_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _3443_ (.A0(\as1802.regs[5][5] ),
    .A1(net59),
    .S(_1237_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _3444_ (.A0(\as1802.regs[5][6] ),
    .A1(net57),
    .S(_1237_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _3445_ (.A0(\as1802.regs[5][7] ),
    .A1(net55),
    .S(_1237_),
    .X(_0127_));
 sky130_fd_sc_hd__and3_4 _3446_ (.A(net73),
    .B(_1190_),
    .C(_1194_),
    .X(_1238_));
 sky130_fd_sc_hd__mux2_1 _3447_ (.A0(\as1802.regs[4][0] ),
    .A1(net69),
    .S(_1238_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(\as1802.regs[4][1] ),
    .A1(net67),
    .S(_1238_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(\as1802.regs[4][2] ),
    .A1(net65),
    .S(_1238_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _3450_ (.A0(\as1802.regs[4][3] ),
    .A1(net63),
    .S(_1238_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _3451_ (.A0(\as1802.regs[4][4] ),
    .A1(net61),
    .S(_1238_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _3452_ (.A0(\as1802.regs[4][5] ),
    .A1(net59),
    .S(_1238_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _3453_ (.A0(\as1802.regs[4][6] ),
    .A1(net57),
    .S(_1238_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _3454_ (.A0(\as1802.regs[4][7] ),
    .A1(net55),
    .S(_1238_),
    .X(_0135_));
 sky130_fd_sc_hd__and3_4 _3455_ (.A(_2117_),
    .B(net73),
    .C(_1191_),
    .X(_1239_));
 sky130_fd_sc_hd__mux2_1 _3456_ (.A0(\as1802.regs[3][0] ),
    .A1(net68),
    .S(_1239_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _3457_ (.A0(\as1802.regs[3][1] ),
    .A1(net67),
    .S(_1239_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _3458_ (.A0(\as1802.regs[3][2] ),
    .A1(net64),
    .S(_1239_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _3459_ (.A0(\as1802.regs[3][3] ),
    .A1(net63),
    .S(_1239_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _3460_ (.A0(\as1802.regs[3][4] ),
    .A1(net61),
    .S(_1239_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _3461_ (.A0(\as1802.regs[3][5] ),
    .A1(net59),
    .S(_1239_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _3462_ (.A0(\as1802.regs[3][6] ),
    .A1(net57),
    .S(_1239_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _3463_ (.A0(\as1802.regs[3][7] ),
    .A1(net55),
    .S(_1239_),
    .X(_0143_));
 sky130_fd_sc_hd__and3_4 _3464_ (.A(net73),
    .B(_0758_),
    .C(_1191_),
    .X(_1240_));
 sky130_fd_sc_hd__mux2_1 _3465_ (.A0(\as1802.regs[2][0] ),
    .A1(net68),
    .S(_1240_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _3466_ (.A0(\as1802.regs[2][1] ),
    .A1(net67),
    .S(_1240_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _3467_ (.A0(\as1802.regs[2][2] ),
    .A1(net64),
    .S(_1240_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _3468_ (.A0(\as1802.regs[2][3] ),
    .A1(net63),
    .S(_1240_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _3469_ (.A0(\as1802.regs[2][4] ),
    .A1(net60),
    .S(_1240_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _3470_ (.A0(\as1802.regs[2][5] ),
    .A1(net59),
    .S(_1240_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _3471_ (.A0(\as1802.regs[2][6] ),
    .A1(net57),
    .S(_1240_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _3472_ (.A0(\as1802.regs[2][7] ),
    .A1(net55),
    .S(_1240_),
    .X(_0151_));
 sky130_fd_sc_hd__and3_4 _3473_ (.A(net73),
    .B(_1191_),
    .C(_1196_),
    .X(_1241_));
 sky130_fd_sc_hd__mux2_1 _3474_ (.A0(\as1802.regs[1][0] ),
    .A1(net69),
    .S(_1241_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _3475_ (.A0(\as1802.regs[1][1] ),
    .A1(net67),
    .S(_1241_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _3476_ (.A0(\as1802.regs[1][2] ),
    .A1(net65),
    .S(_1241_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _3477_ (.A0(\as1802.regs[1][3] ),
    .A1(net63),
    .S(_1241_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _3478_ (.A0(\as1802.regs[1][4] ),
    .A1(net61),
    .S(_1241_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _3479_ (.A0(\as1802.regs[1][5] ),
    .A1(net59),
    .S(_1241_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _3480_ (.A0(\as1802.regs[1][6] ),
    .A1(net57),
    .S(_1241_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _3481_ (.A0(\as1802.regs[1][7] ),
    .A1(net55),
    .S(_1241_),
    .X(_0159_));
 sky130_fd_sc_hd__and3_4 _3482_ (.A(_2117_),
    .B(_2124_),
    .C(net70),
    .X(_1242_));
 sky130_fd_sc_hd__mux2_1 _3483_ (.A0(\as1802.regs[15][8] ),
    .A1(net52),
    .S(_1242_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _3484_ (.A0(\as1802.regs[15][9] ),
    .A1(net50),
    .S(_1242_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _3485_ (.A0(\as1802.regs[15][10] ),
    .A1(net49),
    .S(_1242_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(\as1802.regs[15][11] ),
    .A1(net46),
    .S(_1242_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _3487_ (.A0(\as1802.regs[15][12] ),
    .A1(net44),
    .S(_1242_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _3488_ (.A0(\as1802.regs[15][13] ),
    .A1(net42),
    .S(_1242_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _3489_ (.A0(\as1802.regs[15][14] ),
    .A1(net40),
    .S(_1242_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _3490_ (.A0(\as1802.regs[15][15] ),
    .A1(net38),
    .S(_1242_),
    .X(_0167_));
 sky130_fd_sc_hd__and3_4 _3491_ (.A(_2124_),
    .B(net72),
    .C(_0758_),
    .X(_1243_));
 sky130_fd_sc_hd__mux2_1 _3492_ (.A0(\as1802.regs[14][0] ),
    .A1(net68),
    .S(_1243_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _3493_ (.A0(\as1802.regs[14][1] ),
    .A1(net66),
    .S(_1243_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _3494_ (.A0(\as1802.regs[14][2] ),
    .A1(net64),
    .S(_1243_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _3495_ (.A0(\as1802.regs[14][3] ),
    .A1(net62),
    .S(_1243_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _3496_ (.A0(\as1802.regs[14][4] ),
    .A1(net60),
    .S(_1243_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _3497_ (.A0(\as1802.regs[14][5] ),
    .A1(net58),
    .S(_1243_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _3498_ (.A0(\as1802.regs[14][6] ),
    .A1(net56),
    .S(_1243_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _3499_ (.A0(\as1802.regs[14][7] ),
    .A1(net54),
    .S(_1243_),
    .X(_0175_));
 sky130_fd_sc_hd__and3_4 _3500_ (.A(_2124_),
    .B(net72),
    .C(_1196_),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_1 _3501_ (.A0(\as1802.regs[13][0] ),
    .A1(net68),
    .S(_1244_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _3502_ (.A0(\as1802.regs[13][1] ),
    .A1(net66),
    .S(_1244_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _3503_ (.A0(\as1802.regs[13][2] ),
    .A1(net64),
    .S(_1244_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _3504_ (.A0(\as1802.regs[13][3] ),
    .A1(net62),
    .S(_1244_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _3505_ (.A0(\as1802.regs[13][4] ),
    .A1(net60),
    .S(_1244_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _3506_ (.A0(\as1802.regs[13][5] ),
    .A1(net58),
    .S(_1244_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _3507_ (.A0(\as1802.regs[13][6] ),
    .A1(net56),
    .S(_1244_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _3508_ (.A0(\as1802.regs[13][7] ),
    .A1(net54),
    .S(_1244_),
    .X(_0183_));
 sky130_fd_sc_hd__and3_4 _3509_ (.A(_2124_),
    .B(net70),
    .C(_1190_),
    .X(_1245_));
 sky130_fd_sc_hd__mux2_1 _3510_ (.A0(\as1802.regs[12][8] ),
    .A1(net52),
    .S(_1245_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _3511_ (.A0(\as1802.regs[12][9] ),
    .A1(net50),
    .S(_1245_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _3512_ (.A0(\as1802.regs[12][10] ),
    .A1(net48),
    .S(_1245_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _3513_ (.A0(\as1802.regs[12][11] ),
    .A1(net46),
    .S(_1245_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _3514_ (.A0(\as1802.regs[12][12] ),
    .A1(net44),
    .S(_1245_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _3515_ (.A0(\as1802.regs[12][13] ),
    .A1(net42),
    .S(_1245_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _3516_ (.A0(\as1802.regs[12][14] ),
    .A1(net40),
    .S(_1245_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _3517_ (.A0(\as1802.regs[12][15] ),
    .A1(net38),
    .S(_1245_),
    .X(_0191_));
 sky130_fd_sc_hd__and3_4 _3518_ (.A(_2117_),
    .B(net72),
    .C(_0759_),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_1 _3519_ (.A0(\as1802.regs[11][0] ),
    .A1(net68),
    .S(_1246_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _3520_ (.A0(\as1802.regs[11][1] ),
    .A1(net66),
    .S(_1246_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _3521_ (.A0(\as1802.regs[11][2] ),
    .A1(net64),
    .S(_1246_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _3522_ (.A0(\as1802.regs[11][3] ),
    .A1(net62),
    .S(_1246_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _3523_ (.A0(\as1802.regs[11][4] ),
    .A1(net60),
    .S(_1246_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _3524_ (.A0(\as1802.regs[11][5] ),
    .A1(net58),
    .S(_1246_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _3525_ (.A0(\as1802.regs[11][6] ),
    .A1(net56),
    .S(_1246_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _3526_ (.A0(\as1802.regs[11][7] ),
    .A1(net54),
    .S(_1246_),
    .X(_0199_));
 sky130_fd_sc_hd__and3_4 _3527_ (.A(net72),
    .B(_0758_),
    .C(_0759_),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _3528_ (.A0(\as1802.regs[10][0] ),
    .A1(net68),
    .S(_1247_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _3529_ (.A0(\as1802.regs[10][1] ),
    .A1(net66),
    .S(_1247_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _3530_ (.A0(\as1802.regs[10][2] ),
    .A1(net64),
    .S(_1247_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _3531_ (.A0(\as1802.regs[10][3] ),
    .A1(net62),
    .S(_1247_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _3532_ (.A0(\as1802.regs[10][4] ),
    .A1(net60),
    .S(_1247_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _3533_ (.A0(\as1802.regs[10][5] ),
    .A1(net58),
    .S(_1247_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_1 _3534_ (.A0(\as1802.regs[10][6] ),
    .A1(net56),
    .S(_1247_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _3535_ (.A0(\as1802.regs[10][7] ),
    .A1(net54),
    .S(_1247_),
    .X(_0207_));
 sky130_fd_sc_hd__and3_4 _3536_ (.A(net73),
    .B(_1190_),
    .C(_1191_),
    .X(_1248_));
 sky130_fd_sc_hd__mux2_1 _3537_ (.A0(\as1802.regs[0][0] ),
    .A1(net69),
    .S(_1248_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _3538_ (.A0(\as1802.regs[0][1] ),
    .A1(net67),
    .S(_1248_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _3539_ (.A0(\as1802.regs[0][2] ),
    .A1(net65),
    .S(_1248_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _3540_ (.A0(\as1802.regs[0][3] ),
    .A1(net63),
    .S(_1248_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _3541_ (.A0(\as1802.regs[0][4] ),
    .A1(net61),
    .S(_1248_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _3542_ (.A0(\as1802.regs[0][5] ),
    .A1(net59),
    .S(_1248_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _3543_ (.A0(\as1802.regs[0][6] ),
    .A1(net57),
    .S(_1248_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _3544_ (.A0(\as1802.regs[0][7] ),
    .A1(net55),
    .S(_1248_),
    .X(_0215_));
 sky130_fd_sc_hd__and3_4 _3545_ (.A(_2124_),
    .B(_0758_),
    .C(net70),
    .X(_1249_));
 sky130_fd_sc_hd__mux2_1 _3546_ (.A0(\as1802.regs[14][8] ),
    .A1(net52),
    .S(_1249_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _3547_ (.A0(\as1802.regs[14][9] ),
    .A1(net50),
    .S(_1249_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _3548_ (.A0(\as1802.regs[14][10] ),
    .A1(net49),
    .S(_1249_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _3549_ (.A0(\as1802.regs[14][11] ),
    .A1(net46),
    .S(_1249_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _3550_ (.A0(\as1802.regs[14][12] ),
    .A1(net44),
    .S(_1249_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _3551_ (.A0(\as1802.regs[14][13] ),
    .A1(net42),
    .S(_1249_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _3552_ (.A0(\as1802.regs[14][14] ),
    .A1(net40),
    .S(_1249_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _3553_ (.A0(\as1802.regs[14][15] ),
    .A1(net38),
    .S(_1249_),
    .X(_0223_));
 sky130_fd_sc_hd__and3_4 _3554_ (.A(_2124_),
    .B(net70),
    .C(_1196_),
    .X(_1250_));
 sky130_fd_sc_hd__mux2_1 _3555_ (.A0(\as1802.regs[13][8] ),
    .A1(net52),
    .S(_1250_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _3556_ (.A0(\as1802.regs[13][9] ),
    .A1(net51),
    .S(_1250_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _3557_ (.A0(\as1802.regs[13][10] ),
    .A1(net48),
    .S(_1250_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _3558_ (.A0(\as1802.regs[13][11] ),
    .A1(net46),
    .S(_1250_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _3559_ (.A0(\as1802.regs[13][12] ),
    .A1(net44),
    .S(_1250_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _3560_ (.A0(\as1802.regs[13][13] ),
    .A1(net42),
    .S(_1250_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_1 _3561_ (.A0(\as1802.regs[13][14] ),
    .A1(net40),
    .S(_1250_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _3562_ (.A0(\as1802.regs[13][15] ),
    .A1(net38),
    .S(_1250_),
    .X(_0231_));
 sky130_fd_sc_hd__and3_4 _3563_ (.A(_2124_),
    .B(net72),
    .C(_1190_),
    .X(_1251_));
 sky130_fd_sc_hd__mux2_1 _3564_ (.A0(\as1802.regs[12][0] ),
    .A1(net68),
    .S(_1251_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(\as1802.regs[12][1] ),
    .A1(net66),
    .S(_1251_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _3566_ (.A0(\as1802.regs[12][2] ),
    .A1(net64),
    .S(_1251_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _3567_ (.A0(\as1802.regs[12][3] ),
    .A1(net62),
    .S(_1251_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _3568_ (.A0(\as1802.regs[12][4] ),
    .A1(net60),
    .S(_1251_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _3569_ (.A0(\as1802.regs[12][5] ),
    .A1(net58),
    .S(_1251_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _3570_ (.A0(\as1802.regs[12][6] ),
    .A1(net56),
    .S(_1251_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _3571_ (.A0(\as1802.regs[12][7] ),
    .A1(net54),
    .S(_1251_),
    .X(_0239_));
 sky130_fd_sc_hd__and3_4 _3572_ (.A(_2117_),
    .B(_0759_),
    .C(net71),
    .X(_1252_));
 sky130_fd_sc_hd__mux2_1 _3573_ (.A0(\as1802.regs[11][8] ),
    .A1(net52),
    .S(_1252_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _3574_ (.A0(\as1802.regs[11][9] ),
    .A1(net50),
    .S(_1252_),
    .X(_0241_));
 sky130_fd_sc_hd__mux2_1 _3575_ (.A0(\as1802.regs[11][10] ),
    .A1(net48),
    .S(_1252_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _3576_ (.A0(\as1802.regs[11][11] ),
    .A1(net46),
    .S(_1252_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _3577_ (.A0(\as1802.regs[11][12] ),
    .A1(net44),
    .S(_1252_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _3578_ (.A0(\as1802.regs[11][13] ),
    .A1(net43),
    .S(_1252_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _3579_ (.A0(\as1802.regs[11][14] ),
    .A1(net40),
    .S(_1252_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _3580_ (.A0(\as1802.regs[11][15] ),
    .A1(net39),
    .S(_1252_),
    .X(_0247_));
 sky130_fd_sc_hd__and4_1 _3581_ (.A(_1912_),
    .B(net268),
    .C(_1950_),
    .D(_1958_),
    .X(_1253_));
 sky130_fd_sc_hd__a2bb2o_1 _3582_ (.A1_N(_1991_),
    .A2_N(_2051_),
    .B1(_1253_),
    .B2(_2011_),
    .X(_1254_));
 sky130_fd_sc_hd__o21ai_4 _3583_ (.A1(net230),
    .A2(_1986_),
    .B1(_2091_),
    .Y(_1255_));
 sky130_fd_sc_hd__nor2_2 _3584_ (.A(net233),
    .B(_1964_),
    .Y(_1256_));
 sky130_fd_sc_hd__nand2_4 _3585_ (.A(net202),
    .B(_1963_),
    .Y(_1257_));
 sky130_fd_sc_hd__o21ai_2 _3586_ (.A1(net229),
    .A2(_1257_),
    .B1(_1221_),
    .Y(_1258_));
 sky130_fd_sc_hd__nor2_1 _3587_ (.A(_1255_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__o21ba_1 _3588_ (.A1(_1959_),
    .A2(_2014_),
    .B1_N(_2043_),
    .X(_1260_));
 sky130_fd_sc_hd__o31a_1 _3589_ (.A1(_1254_),
    .A2(_1259_),
    .A3(_1260_),
    .B1(net195),
    .X(_1261_));
 sky130_fd_sc_hd__xnor2_1 _3590_ (.A(\as1802.last_hi_addr[6] ),
    .B(\as1802.addr_buff[14] ),
    .Y(_1262_));
 sky130_fd_sc_hd__xnor2_1 _3591_ (.A(\as1802.last_hi_addr[4] ),
    .B(\as1802.addr_buff[12] ),
    .Y(_1263_));
 sky130_fd_sc_hd__xnor2_1 _3592_ (.A(\as1802.last_hi_addr[1] ),
    .B(\as1802.addr_buff[9] ),
    .Y(_1264_));
 sky130_fd_sc_hd__o221a_1 _3593_ (.A1(\as1802.last_hi_addr[7] ),
    .A2(_1915_),
    .B1(_1916_),
    .B2(\as1802.addr_buff[13] ),
    .C1(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__xnor2_1 _3594_ (.A(\as1802.last_hi_addr[3] ),
    .B(\as1802.addr_buff[11] ),
    .Y(_1266_));
 sky130_fd_sc_hd__o221a_1 _3595_ (.A1(\as1802.last_hi_addr[5] ),
    .A2(_1917_),
    .B1(_1918_),
    .B2(\as1802.addr_buff[8] ),
    .C1(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__o221a_1 _3596_ (.A1(_1914_),
    .A2(\as1802.addr_buff[15] ),
    .B1(\as1802.last_hi_addr[0] ),
    .B2(_1919_),
    .C1(_1263_),
    .X(_1268_));
 sky130_fd_sc_hd__xnor2_1 _3597_ (.A(\as1802.last_hi_addr[2] ),
    .B(\as1802.addr_buff[10] ),
    .Y(_1269_));
 sky130_fd_sc_hd__and3_1 _3598_ (.A(_1262_),
    .B(_1268_),
    .C(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__a31o_4 _3599_ (.A1(_1265_),
    .A2(_1267_),
    .A3(_1270_),
    .B1(net238),
    .X(_1271_));
 sky130_fd_sc_hd__a21oi_1 _3600_ (.A1(_1920_),
    .A2(_1271_),
    .B1(_1921_),
    .Y(_1272_));
 sky130_fd_sc_hd__or3b_1 _3601_ (.A(net203),
    .B(_2038_),
    .C_N(_1960_),
    .X(_1273_));
 sky130_fd_sc_hd__nor2_1 _3602_ (.A(net193),
    .B(_1203_),
    .Y(_1274_));
 sky130_fd_sc_hd__a21o_1 _3603_ (.A1(\as1802.mem_cycle[0] ),
    .A2(\as1802.mem_write ),
    .B1(net280),
    .X(_1275_));
 sky130_fd_sc_hd__nor3b_1 _3604_ (.A(_1275_),
    .B(_1274_),
    .C_N(_1273_),
    .Y(_1276_));
 sky130_fd_sc_hd__or3b_1 _3605_ (.A(net193),
    .B(_1943_),
    .C_N(_1208_),
    .X(_1277_));
 sky130_fd_sc_hd__nor2_1 _3606_ (.A(net272),
    .B(_2099_),
    .Y(_1278_));
 sky130_fd_sc_hd__nand2_1 _3607_ (.A(_1943_),
    .B(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__nor2_1 _3608_ (.A(net193),
    .B(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__o311a_1 _3609_ (.A1(_1946_),
    .A2(_2026_),
    .A3(_1220_),
    .B1(_1276_),
    .C1(_1277_),
    .X(_1281_));
 sky130_fd_sc_hd__o31ai_2 _3610_ (.A1(_1924_),
    .A2(_1939_),
    .A3(_2044_),
    .B1(_2079_),
    .Y(_1282_));
 sky130_fd_sc_hd__a31o_1 _3611_ (.A1(_2063_),
    .A2(_0378_),
    .A3(_1218_),
    .B1(_2044_),
    .X(_1283_));
 sky130_fd_sc_hd__and4bb_1 _3612_ (.A_N(_1280_),
    .B_N(_1282_),
    .C(_1283_),
    .D(_2154_),
    .X(_1284_));
 sky130_fd_sc_hd__and4bb_1 _3613_ (.A_N(_1261_),
    .B_N(_1272_),
    .C(_1281_),
    .D(_1284_),
    .X(_0248_));
 sky130_fd_sc_hd__nand2_1 _3614_ (.A(net238),
    .B(_1921_),
    .Y(_1285_));
 sky130_fd_sc_hd__nor2_4 _3615_ (.A(\as1802.mem_cycle[2] ),
    .B(_1921_),
    .Y(_1286_));
 sky130_fd_sc_hd__nand2_8 _3616_ (.A(_1920_),
    .B(\as1802.mem_cycle[0] ),
    .Y(_1287_));
 sky130_fd_sc_hd__or2_1 _3617_ (.A(net238),
    .B(_1921_),
    .X(_1288_));
 sky130_fd_sc_hd__nor2_8 _3618_ (.A(net238),
    .B(_1287_),
    .Y(_1289_));
 sky130_fd_sc_hd__or2_1 _3619_ (.A(_1271_),
    .B(_1287_),
    .X(_1290_));
 sky130_fd_sc_hd__a21oi_1 _3620_ (.A1(_1285_),
    .A2(_1290_),
    .B1(net280),
    .Y(_0249_));
 sky130_fd_sc_hd__a211oi_1 _3621_ (.A1(_1920_),
    .A2(_1921_),
    .B1(net280),
    .C1(_1272_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand2_1 _3622_ (.A(\as1802.instr_latch[4] ),
    .B(net223),
    .Y(_1291_));
 sky130_fd_sc_hd__and4_1 _3623_ (.A(_1912_),
    .B(net224),
    .C(net220),
    .D(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__or4_1 _3624_ (.A(net280),
    .B(net192),
    .C(_1208_),
    .D(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__o221a_1 _3625_ (.A1(_1958_),
    .A2(_2043_),
    .B1(_1219_),
    .B2(_1961_),
    .C1(_1279_),
    .X(_1294_));
 sky130_fd_sc_hd__o21ai_1 _3626_ (.A1(_2026_),
    .A2(_1220_),
    .B1(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__or3b_1 _3627_ (.A(_1293_),
    .B(_1295_),
    .C_N(_2064_),
    .X(_1296_));
 sky130_fd_sc_hd__nor2_1 _3628_ (.A(_1254_),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__nor2_4 _3629_ (.A(net201),
    .B(_1989_),
    .Y(_1298_));
 sky130_fd_sc_hd__or4b_4 _3630_ (.A(_2068_),
    .B(_1212_),
    .C(_1259_),
    .D_N(_1297_),
    .X(_1299_));
 sky130_fd_sc_hd__o21ba_4 _3631_ (.A1(_2022_),
    .A2(_2092_),
    .B1_N(_2029_),
    .X(_1300_));
 sky130_fd_sc_hd__a31o_2 _3632_ (.A1(net175),
    .A2(_2021_),
    .A3(net167),
    .B1(_2029_),
    .X(_1301_));
 sky130_fd_sc_hd__or2_2 _3633_ (.A(_1943_),
    .B(_2029_),
    .X(_1302_));
 sky130_fd_sc_hd__nand2_8 _3634_ (.A(net176),
    .B(_2020_),
    .Y(_1303_));
 sky130_fd_sc_hd__o21ai_1 _3635_ (.A1(net230),
    .A2(net82),
    .B1(_2141_),
    .Y(_1304_));
 sky130_fd_sc_hd__mux2_1 _3636_ (.A0(net155),
    .A1(_1304_),
    .S(net189),
    .X(_1305_));
 sky130_fd_sc_hd__o22a_1 _3637_ (.A1(net135),
    .A2(_1304_),
    .B1(_1305_),
    .B2(net175),
    .X(_1306_));
 sky130_fd_sc_hd__o31a_1 _3638_ (.A1(\as1802.regs[2][0] ),
    .A2(_2022_),
    .A3(net167),
    .B1(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__o2bb2a_1 _3639_ (.A1_N(net82),
    .A2_N(net138),
    .B1(net136),
    .B2(_1307_),
    .X(_1308_));
 sky130_fd_sc_hd__nor2_1 _3640_ (.A(net159),
    .B(_1308_),
    .Y(_1309_));
 sky130_fd_sc_hd__a221o_1 _3641_ (.A1(net183),
    .A2(net82),
    .B1(net159),
    .B2(_2138_),
    .C1(net77),
    .X(_1310_));
 sky130_fd_sc_hd__a2bb2o_1 _3642_ (.A1_N(_1309_),
    .A2_N(_1310_),
    .B1(\as1802.addr_buff[0] ),
    .B2(net75),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _3643_ (.A(net226),
    .B(net164),
    .Y(_1311_));
 sky130_fd_sc_hd__o21ai_1 _3644_ (.A1(net226),
    .A2(_0398_),
    .B1(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__mux2_1 _3645_ (.A0(net164),
    .A1(_1312_),
    .S(net190),
    .X(_1313_));
 sky130_fd_sc_hd__o22a_1 _3646_ (.A1(net135),
    .A2(_1312_),
    .B1(_1313_),
    .B2(net175),
    .X(_1314_));
 sky130_fd_sc_hd__o31a_1 _3647_ (.A1(\as1802.regs[2][1] ),
    .A2(net171),
    .A3(net167),
    .B1(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__o2bb2a_1 _3648_ (.A1_N(_0398_),
    .A2_N(net138),
    .B1(net136),
    .B2(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__o21ba_1 _3649_ (.A1(net164),
    .A2(net162),
    .B1_N(net76),
    .X(_1317_));
 sky130_fd_sc_hd__o2bb2a_2 _3650_ (.A1_N(net183),
    .A2_N(_0398_),
    .B1(net159),
    .B2(_1316_),
    .X(_1318_));
 sky130_fd_sc_hd__a22o_1 _3651_ (.A1(\as1802.addr_buff[1] ),
    .A2(net76),
    .B1(_1317_),
    .B2(_1318_),
    .X(_0252_));
 sky130_fd_sc_hd__nand2_1 _3652_ (.A(net225),
    .B(_0458_),
    .Y(_1319_));
 sky130_fd_sc_hd__nor2_1 _3653_ (.A(net189),
    .B(_0459_),
    .Y(_1320_));
 sky130_fd_sc_hd__or3_1 _3654_ (.A(\as1802.regs[2][2] ),
    .B(net169),
    .C(net166),
    .X(_1321_));
 sky130_fd_sc_hd__o21ai_1 _3655_ (.A1(net225),
    .A2(_0445_),
    .B1(_1319_),
    .Y(_1322_));
 sky130_fd_sc_hd__a211o_1 _3656_ (.A1(net189),
    .A2(_1322_),
    .B1(_1320_),
    .C1(net174),
    .X(_1323_));
 sky130_fd_sc_hd__o211a_1 _3657_ (.A1(net135),
    .A2(_1322_),
    .B1(_1323_),
    .C1(_1321_),
    .X(_1324_));
 sky130_fd_sc_hd__a2bb2o_1 _3658_ (.A1_N(net136),
    .A2_N(_1324_),
    .B1(_0445_),
    .B2(net138),
    .X(_1325_));
 sky130_fd_sc_hd__a221o_1 _3659_ (.A1(net183),
    .A2(_0445_),
    .B1(_0459_),
    .B2(net159),
    .C1(net77),
    .X(_1326_));
 sky130_fd_sc_hd__a21oi_2 _3660_ (.A1(net161),
    .A2(_1325_),
    .B1(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__a21o_1 _3661_ (.A1(\as1802.addr_buff[2] ),
    .A2(net75),
    .B1(_1327_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _3662_ (.A0(_0496_),
    .A1(_0510_),
    .S(net226),
    .X(_1328_));
 sky130_fd_sc_hd__mux2_1 _3663_ (.A0(_0510_),
    .A1(_1328_),
    .S(net190),
    .X(_1329_));
 sky130_fd_sc_hd__o22a_1 _3664_ (.A1(net135),
    .A2(_1328_),
    .B1(_1329_),
    .B2(net175),
    .X(_1330_));
 sky130_fd_sc_hd__o31a_2 _3665_ (.A1(\as1802.regs[2][3] ),
    .A2(net169),
    .A3(net167),
    .B1(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__o22a_1 _3666_ (.A1(_0496_),
    .A2(_1300_),
    .B1(net136),
    .B2(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__o22a_1 _3667_ (.A1(_1944_),
    .A2(_0496_),
    .B1(_1332_),
    .B2(_1993_),
    .X(_1333_));
 sky130_fd_sc_hd__o22a_1 _3668_ (.A1(_0510_),
    .A2(net162),
    .B1(_1333_),
    .B2(net274),
    .X(_1334_));
 sky130_fd_sc_hd__mux2_1 _3669_ (.A0(_1334_),
    .A1(\as1802.addr_buff[3] ),
    .S(net76),
    .X(_0254_));
 sky130_fd_sc_hd__nand2_1 _3670_ (.A(net225),
    .B(_0571_),
    .Y(_1335_));
 sky130_fd_sc_hd__nor2_1 _3671_ (.A(net189),
    .B(_0572_),
    .Y(_1336_));
 sky130_fd_sc_hd__or3_1 _3672_ (.A(\as1802.regs[2][4] ),
    .B(net169),
    .C(net167),
    .X(_1337_));
 sky130_fd_sc_hd__o21ai_1 _3673_ (.A1(net225),
    .A2(net78),
    .B1(_1335_),
    .Y(_1338_));
 sky130_fd_sc_hd__a211o_1 _3674_ (.A1(net190),
    .A2(_1338_),
    .B1(_1336_),
    .C1(net174),
    .X(_1339_));
 sky130_fd_sc_hd__o211a_1 _3675_ (.A1(net135),
    .A2(_1338_),
    .B1(_1339_),
    .C1(_1337_),
    .X(_1340_));
 sky130_fd_sc_hd__a2bb2o_2 _3676_ (.A1_N(net136),
    .A2_N(_1340_),
    .B1(net78),
    .B2(net138),
    .X(_1341_));
 sky130_fd_sc_hd__a221o_2 _3677_ (.A1(net183),
    .A2(net78),
    .B1(_0572_),
    .B2(net159),
    .C1(net77),
    .X(_1342_));
 sky130_fd_sc_hd__a21oi_4 _3678_ (.A1(net161),
    .A2(_1341_),
    .B1(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__a21o_1 _3679_ (.A1(\as1802.addr_buff[4] ),
    .A2(net76),
    .B1(_1343_),
    .X(_0255_));
 sky130_fd_sc_hd__nand2_1 _3680_ (.A(net226),
    .B(net163),
    .Y(_1344_));
 sky130_fd_sc_hd__o21ai_1 _3681_ (.A1(net226),
    .A2(_0610_),
    .B1(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__mux2_1 _3682_ (.A0(net163),
    .A1(_1345_),
    .S(net189),
    .X(_1346_));
 sky130_fd_sc_hd__o22a_1 _3683_ (.A1(net135),
    .A2(_1345_),
    .B1(_1346_),
    .B2(net174),
    .X(_1347_));
 sky130_fd_sc_hd__o31a_1 _3684_ (.A1(\as1802.regs[2][5] ),
    .A2(net169),
    .A3(net166),
    .B1(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__a2bb2o_1 _3685_ (.A1_N(net136),
    .A2_N(_1348_),
    .B1(_0610_),
    .B2(net138),
    .X(_1349_));
 sky130_fd_sc_hd__o21bai_1 _3686_ (.A1(net163),
    .A2(net161),
    .B1_N(net77),
    .Y(_1350_));
 sky130_fd_sc_hd__a221o_2 _3687_ (.A1(net183),
    .A2(_0610_),
    .B1(net161),
    .B2(_1349_),
    .C1(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__a21bo_1 _3688_ (.A1(\as1802.addr_buff[5] ),
    .A2(net74),
    .B1_N(_1351_),
    .X(_0256_));
 sky130_fd_sc_hd__nand2_1 _3689_ (.A(net226),
    .B(_0680_),
    .Y(_1352_));
 sky130_fd_sc_hd__nor2_1 _3690_ (.A(net189),
    .B(_0681_),
    .Y(_1353_));
 sky130_fd_sc_hd__or3_1 _3691_ (.A(\as1802.regs[2][6] ),
    .B(net169),
    .C(net166),
    .X(_1354_));
 sky130_fd_sc_hd__o21ai_1 _3692_ (.A1(net225),
    .A2(_0667_),
    .B1(_1352_),
    .Y(_1355_));
 sky130_fd_sc_hd__a211o_1 _3693_ (.A1(net189),
    .A2(_1355_),
    .B1(_1353_),
    .C1(net174),
    .X(_1356_));
 sky130_fd_sc_hd__o211a_1 _3694_ (.A1(net135),
    .A2(_1355_),
    .B1(_1356_),
    .C1(_1354_),
    .X(_1357_));
 sky130_fd_sc_hd__a2bb2o_2 _3695_ (.A1_N(net136),
    .A2_N(_1357_),
    .B1(_0667_),
    .B2(net138),
    .X(_1358_));
 sky130_fd_sc_hd__a221o_2 _3696_ (.A1(net183),
    .A2(_0667_),
    .B1(_0681_),
    .B2(net159),
    .C1(net77),
    .X(_1359_));
 sky130_fd_sc_hd__a21oi_4 _3697_ (.A1(net161),
    .A2(_1358_),
    .B1(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hd__a21o_1 _3698_ (.A1(\as1802.addr_buff[6] ),
    .A2(net76),
    .B1(_1360_),
    .X(_0257_));
 sky130_fd_sc_hd__nand2_1 _3699_ (.A(net225),
    .B(_0732_),
    .Y(_1361_));
 sky130_fd_sc_hd__o21ai_1 _3700_ (.A1(net225),
    .A2(_0716_),
    .B1(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__mux2_1 _3701_ (.A0(_0732_),
    .A1(_1362_),
    .S(net189),
    .X(_1363_));
 sky130_fd_sc_hd__o22a_1 _3702_ (.A1(net135),
    .A2(_1362_),
    .B1(_1363_),
    .B2(net174),
    .X(_1364_));
 sky130_fd_sc_hd__o31a_1 _3703_ (.A1(\as1802.regs[2][7] ),
    .A2(net169),
    .A3(net166),
    .B1(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__a2bb2o_1 _3704_ (.A1_N(net136),
    .A2_N(_1365_),
    .B1(_0716_),
    .B2(net138),
    .X(_1366_));
 sky130_fd_sc_hd__o21bai_1 _3705_ (.A1(_0732_),
    .A2(net161),
    .B1_N(net77),
    .Y(_1367_));
 sky130_fd_sc_hd__a221o_4 _3706_ (.A1(net183),
    .A2(_0716_),
    .B1(net161),
    .B2(_1366_),
    .C1(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__a21bo_1 _3707_ (.A1(\as1802.addr_buff[7] ),
    .A2(net74),
    .B1_N(_1368_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _3708_ (.A0(_0780_),
    .A1(_0800_),
    .S(net228),
    .X(_1369_));
 sky130_fd_sc_hd__mux2_1 _3709_ (.A0(_0800_),
    .A1(_1369_),
    .S(net190),
    .X(_1370_));
 sky130_fd_sc_hd__o22a_1 _3710_ (.A1(\as1802.regs[2][8] ),
    .A2(net166),
    .B1(_1369_),
    .B2(_2021_),
    .X(_1371_));
 sky130_fd_sc_hd__mux2_1 _3711_ (.A0(_1370_),
    .A1(_1371_),
    .S(net174),
    .X(_1372_));
 sky130_fd_sc_hd__o22a_1 _3712_ (.A1(_0780_),
    .A2(_1300_),
    .B1(net137),
    .B2(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__nor2_1 _3713_ (.A(net160),
    .B(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__a221o_2 _3714_ (.A1(net183),
    .A2(_0781_),
    .B1(_0799_),
    .B2(net159),
    .C1(net77),
    .X(_1375_));
 sky130_fd_sc_hd__a2bb2o_1 _3715_ (.A1_N(_1374_),
    .A2_N(_1375_),
    .B1(\as1802.addr_buff[8] ),
    .B2(net74),
    .X(_0259_));
 sky130_fd_sc_hd__nand2_1 _3716_ (.A(net225),
    .B(_0855_),
    .Y(_1376_));
 sky130_fd_sc_hd__o21ai_1 _3717_ (.A1(net225),
    .A2(_0837_),
    .B1(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__mux2_1 _3718_ (.A0(_0855_),
    .A1(_1377_),
    .S(net189),
    .X(_1378_));
 sky130_fd_sc_hd__o22a_1 _3719_ (.A1(\as1802.regs[2][9] ),
    .A2(net166),
    .B1(_1377_),
    .B2(_2021_),
    .X(_1379_));
 sky130_fd_sc_hd__mux2_1 _3720_ (.A0(_1378_),
    .A1(_1379_),
    .S(net174),
    .X(_1380_));
 sky130_fd_sc_hd__a2bb2o_1 _3721_ (.A1_N(net136),
    .A2_N(_1380_),
    .B1(_0837_),
    .B2(net138),
    .X(_1381_));
 sky130_fd_sc_hd__a221o_1 _3722_ (.A1(net183),
    .A2(_0837_),
    .B1(_0856_),
    .B2(net159),
    .C1(net77),
    .X(_1382_));
 sky130_fd_sc_hd__a21oi_2 _3723_ (.A1(net161),
    .A2(_1381_),
    .B1(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__a21o_1 _3724_ (.A1(\as1802.addr_buff[9] ),
    .A2(net74),
    .B1(_1383_),
    .X(_0260_));
 sky130_fd_sc_hd__nand2_1 _3725_ (.A(net228),
    .B(_0908_),
    .Y(_1384_));
 sky130_fd_sc_hd__o21ai_1 _3726_ (.A1(net228),
    .A2(_0891_),
    .B1(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__mux2_1 _3727_ (.A0(_0908_),
    .A1(_1385_),
    .S(net189),
    .X(_1386_));
 sky130_fd_sc_hd__o22a_1 _3728_ (.A1(net135),
    .A2(_1385_),
    .B1(_1386_),
    .B2(net174),
    .X(_1387_));
 sky130_fd_sc_hd__o31a_1 _3729_ (.A1(\as1802.regs[2][10] ),
    .A2(net169),
    .A3(net166),
    .B1(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__a2bb2o_1 _3730_ (.A1_N(net136),
    .A2_N(_1388_),
    .B1(_0891_),
    .B2(net138),
    .X(_1389_));
 sky130_fd_sc_hd__a221o_1 _3731_ (.A1(net183),
    .A2(_0891_),
    .B1(_0909_),
    .B2(net159),
    .C1(net77),
    .X(_1390_));
 sky130_fd_sc_hd__a21oi_2 _3732_ (.A1(net162),
    .A2(_1389_),
    .B1(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__a21o_1 _3733_ (.A1(\as1802.addr_buff[10] ),
    .A2(net74),
    .B1(_1391_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _3734_ (.A0(_0934_),
    .A1(_0963_),
    .S(net200),
    .X(_1392_));
 sky130_fd_sc_hd__mux2_1 _3735_ (.A0(_0934_),
    .A1(_1392_),
    .S(net190),
    .X(_1393_));
 sky130_fd_sc_hd__o22a_1 _3736_ (.A1(_1303_),
    .A2(_1392_),
    .B1(_1393_),
    .B2(net174),
    .X(_1394_));
 sky130_fd_sc_hd__o31a_1 _3737_ (.A1(\as1802.regs[2][11] ),
    .A2(net169),
    .A3(net166),
    .B1(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__o22a_1 _3738_ (.A1(_0963_),
    .A2(_1300_),
    .B1(net137),
    .B2(_1395_),
    .X(_1396_));
 sky130_fd_sc_hd__or2_1 _3739_ (.A(_0934_),
    .B(net161),
    .X(_1397_));
 sky130_fd_sc_hd__o221a_1 _3740_ (.A1(_2157_),
    .A2(_0963_),
    .B1(net160),
    .B2(_1396_),
    .C1(_1397_),
    .X(_1398_));
 sky130_fd_sc_hd__mux2_1 _3741_ (.A0(_1398_),
    .A1(\as1802.addr_buff[11] ),
    .S(net74),
    .X(_0262_));
 sky130_fd_sc_hd__nand2_1 _3742_ (.A(net228),
    .B(_1011_),
    .Y(_1399_));
 sky130_fd_sc_hd__o21ai_1 _3743_ (.A1(net228),
    .A2(_0997_),
    .B1(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hd__mux2_1 _3744_ (.A0(_1011_),
    .A1(_1400_),
    .S(net190),
    .X(_1401_));
 sky130_fd_sc_hd__o22a_1 _3745_ (.A1(_1303_),
    .A2(_1400_),
    .B1(_1401_),
    .B2(net174),
    .X(_1402_));
 sky130_fd_sc_hd__o31a_1 _3746_ (.A1(\as1802.regs[2][12] ),
    .A2(net169),
    .A3(net166),
    .B1(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__a2bb2o_1 _3747_ (.A1_N(net137),
    .A2_N(_1403_),
    .B1(_0997_),
    .B2(net138),
    .X(_1404_));
 sky130_fd_sc_hd__a2bb2o_1 _3748_ (.A1_N(_1011_),
    .A2_N(net162),
    .B1(_2156_),
    .B2(_0997_),
    .X(_1405_));
 sky130_fd_sc_hd__a211o_1 _3749_ (.A1(net162),
    .A2(_1404_),
    .B1(_1405_),
    .C1(net77),
    .X(_1406_));
 sky130_fd_sc_hd__a21bo_1 _3750_ (.A1(\as1802.addr_buff[12] ),
    .A2(net74),
    .B1_N(_1406_),
    .X(_0263_));
 sky130_fd_sc_hd__nand2_1 _3751_ (.A(net227),
    .B(_1065_),
    .Y(_1407_));
 sky130_fd_sc_hd__o21ai_1 _3752_ (.A1(net227),
    .A2(_1045_),
    .B1(_1407_),
    .Y(_1408_));
 sky130_fd_sc_hd__mux2_1 _3753_ (.A0(_1065_),
    .A1(_1408_),
    .S(_1951_),
    .X(_1409_));
 sky130_fd_sc_hd__o22a_1 _3754_ (.A1(net135),
    .A2(_1408_),
    .B1(_1409_),
    .B2(net177),
    .X(_1410_));
 sky130_fd_sc_hd__o31a_1 _3755_ (.A1(\as1802.regs[2][13] ),
    .A2(_1969_),
    .A3(net166),
    .B1(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__a2bb2o_1 _3756_ (.A1_N(net137),
    .A2_N(_1411_),
    .B1(_1045_),
    .B2(_1301_),
    .X(_1412_));
 sky130_fd_sc_hd__a221o_1 _3757_ (.A1(_2156_),
    .A2(_1045_),
    .B1(_1066_),
    .B2(net160),
    .C1(net75),
    .X(_1413_));
 sky130_fd_sc_hd__a21oi_1 _3758_ (.A1(net161),
    .A2(_1412_),
    .B1(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__a21o_1 _3759_ (.A1(\as1802.addr_buff[13] ),
    .A2(net74),
    .B1(_1414_),
    .X(_0264_));
 sky130_fd_sc_hd__nor2_1 _3760_ (.A(net200),
    .B(_1116_),
    .Y(_1415_));
 sky130_fd_sc_hd__nor2_1 _3761_ (.A(_1951_),
    .B(_1116_),
    .Y(_1416_));
 sky130_fd_sc_hd__or3_1 _3762_ (.A(\as1802.regs[2][14] ),
    .B(net169),
    .C(net168),
    .X(_1417_));
 sky130_fd_sc_hd__a21o_1 _3763_ (.A1(net200),
    .A2(_1101_),
    .B1(_1415_),
    .X(_1418_));
 sky130_fd_sc_hd__a211o_1 _3764_ (.A1(_1951_),
    .A2(_1418_),
    .B1(_1416_),
    .C1(net177),
    .X(_1419_));
 sky130_fd_sc_hd__o211a_1 _3765_ (.A1(_1303_),
    .A2(_1418_),
    .B1(_1419_),
    .C1(_1417_),
    .X(_1420_));
 sky130_fd_sc_hd__o22a_1 _3766_ (.A1(_1101_),
    .A2(_1300_),
    .B1(net137),
    .B2(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__a21oi_1 _3767_ (.A1(_1116_),
    .A2(net160),
    .B1(net75),
    .Y(_1422_));
 sky130_fd_sc_hd__o221a_1 _3768_ (.A1(_2157_),
    .A2(_1101_),
    .B1(net160),
    .B2(_1421_),
    .C1(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__a21o_1 _3769_ (.A1(\as1802.addr_buff[14] ),
    .A2(net74),
    .B1(_1423_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _3770_ (.A0(_1150_),
    .A1(_1165_),
    .S(net227),
    .X(_1424_));
 sky130_fd_sc_hd__mux2_1 _3771_ (.A0(_1165_),
    .A1(_1424_),
    .S(net190),
    .X(_1425_));
 sky130_fd_sc_hd__o22a_1 _3772_ (.A1(\as1802.regs[2][15] ),
    .A2(net168),
    .B1(_1424_),
    .B2(_2021_),
    .X(_1426_));
 sky130_fd_sc_hd__mux2_1 _3773_ (.A0(_1425_),
    .A1(_1426_),
    .S(net177),
    .X(_1427_));
 sky130_fd_sc_hd__o22a_1 _3774_ (.A1(_1150_),
    .A2(_1300_),
    .B1(net137),
    .B2(_1427_),
    .X(_1428_));
 sky130_fd_sc_hd__a21oi_1 _3775_ (.A1(_1164_),
    .A2(net160),
    .B1(net75),
    .Y(_1429_));
 sky130_fd_sc_hd__o221a_1 _3776_ (.A1(_2157_),
    .A2(_1150_),
    .B1(net160),
    .B2(_1428_),
    .C1(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__a21o_1 _3777_ (.A1(\as1802.addr_buff[15] ),
    .A2(net74),
    .B1(_1430_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _3778_ (.A0(\as1802.addr_buff[8] ),
    .A1(\as1802.addr_buff[0] ),
    .S(_1271_),
    .X(_1431_));
 sky130_fd_sc_hd__or2_1 _3779_ (.A(net17),
    .B(_1286_),
    .X(_1432_));
 sky130_fd_sc_hd__o211a_1 _3780_ (.A1(_1287_),
    .A2(_1431_),
    .B1(_1432_),
    .C1(net278),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _3781_ (.A0(\as1802.addr_buff[9] ),
    .A1(\as1802.addr_buff[1] ),
    .S(_1271_),
    .X(_1433_));
 sky130_fd_sc_hd__or2_1 _3782_ (.A(net18),
    .B(_1286_),
    .X(_1434_));
 sky130_fd_sc_hd__o211a_1 _3783_ (.A1(_1287_),
    .A2(_1433_),
    .B1(_1434_),
    .C1(net278),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _3784_ (.A0(\as1802.addr_buff[10] ),
    .A1(\as1802.addr_buff[2] ),
    .S(_1271_),
    .X(_1435_));
 sky130_fd_sc_hd__or2_1 _3785_ (.A(net19),
    .B(_1286_),
    .X(_1436_));
 sky130_fd_sc_hd__o211a_1 _3786_ (.A1(_1287_),
    .A2(_1435_),
    .B1(_1436_),
    .C1(net278),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _3787_ (.A0(\as1802.addr_buff[11] ),
    .A1(\as1802.addr_buff[3] ),
    .S(_1271_),
    .X(_1437_));
 sky130_fd_sc_hd__or2_1 _3788_ (.A(net20),
    .B(_1286_),
    .X(_1438_));
 sky130_fd_sc_hd__o211a_1 _3789_ (.A1(_1287_),
    .A2(_1437_),
    .B1(_1438_),
    .C1(net278),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _3790_ (.A0(\as1802.addr_buff[12] ),
    .A1(\as1802.addr_buff[4] ),
    .S(_1271_),
    .X(_1439_));
 sky130_fd_sc_hd__or2_1 _3791_ (.A(net21),
    .B(_1286_),
    .X(_1440_));
 sky130_fd_sc_hd__o211a_1 _3792_ (.A1(_1287_),
    .A2(_1439_),
    .B1(_1440_),
    .C1(net278),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _3793_ (.A0(\as1802.addr_buff[13] ),
    .A1(\as1802.addr_buff[5] ),
    .S(_1271_),
    .X(_1441_));
 sky130_fd_sc_hd__or2_1 _3794_ (.A(net22),
    .B(_1286_),
    .X(_1442_));
 sky130_fd_sc_hd__o211a_1 _3795_ (.A1(_1287_),
    .A2(_1441_),
    .B1(_1442_),
    .C1(net278),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _3796_ (.A0(\as1802.addr_buff[14] ),
    .A1(\as1802.addr_buff[6] ),
    .S(_1271_),
    .X(_1443_));
 sky130_fd_sc_hd__or2_1 _3797_ (.A(net23),
    .B(_1286_),
    .X(_1444_));
 sky130_fd_sc_hd__o211a_1 _3798_ (.A1(_1287_),
    .A2(_1443_),
    .B1(_1444_),
    .C1(net279),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _3799_ (.A0(\as1802.addr_buff[15] ),
    .A1(\as1802.addr_buff[7] ),
    .S(_1271_),
    .X(_1445_));
 sky130_fd_sc_hd__or2_1 _3800_ (.A(net25),
    .B(_1286_),
    .X(_1446_));
 sky130_fd_sc_hd__o211a_1 _3801_ (.A1(_1287_),
    .A2(_1445_),
    .B1(_1446_),
    .C1(net278),
    .X(_0274_));
 sky130_fd_sc_hd__or2_1 _3802_ (.A(_1920_),
    .B(_1288_),
    .X(_1447_));
 sky130_fd_sc_hd__or3b_4 _3803_ (.A(\as1802.mem_write ),
    .B(_1447_),
    .C_N(net269),
    .X(_1448_));
 sky130_fd_sc_hd__nor2_8 _3804_ (.A(net280),
    .B(_1448_),
    .Y(_1449_));
 sky130_fd_sc_hd__mux2_1 _3805_ (.A0(net237),
    .A1(net1),
    .S(_1449_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _3806_ (.A0(net236),
    .A1(net5),
    .S(_1449_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _3807_ (.A0(net234),
    .A1(net6),
    .S(_1449_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _3808_ (.A0(net226),
    .A1(net7),
    .S(_1449_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _3809_ (.A0(\as1802.instr_latch[4] ),
    .A1(net8),
    .S(_1449_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _3810_ (.A0(net224),
    .A1(net9),
    .S(_1449_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _3811_ (.A0(net222),
    .A1(net10),
    .S(_1449_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _3812_ (.A0(net221),
    .A1(net11),
    .S(_1449_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _3813_ (.A0(_1918_),
    .A1(_1919_),
    .S(_1289_),
    .X(_1450_));
 sky130_fd_sc_hd__nand2_1 _3814_ (.A(net278),
    .B(_1450_),
    .Y(_0283_));
 sky130_fd_sc_hd__mux2_1 _3815_ (.A0(\as1802.last_hi_addr[1] ),
    .A1(\as1802.addr_buff[9] ),
    .S(_1289_),
    .X(_1451_));
 sky130_fd_sc_hd__or2_1 _3816_ (.A(net282),
    .B(_1451_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _3817_ (.A0(\as1802.last_hi_addr[2] ),
    .A1(\as1802.addr_buff[10] ),
    .S(_1289_),
    .X(_1452_));
 sky130_fd_sc_hd__or2_1 _3818_ (.A(net282),
    .B(_1452_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _3819_ (.A0(\as1802.last_hi_addr[3] ),
    .A1(\as1802.addr_buff[11] ),
    .S(_1289_),
    .X(_1453_));
 sky130_fd_sc_hd__or2_1 _3820_ (.A(net282),
    .B(_1453_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _3821_ (.A0(\as1802.last_hi_addr[4] ),
    .A1(\as1802.addr_buff[12] ),
    .S(_1289_),
    .X(_1454_));
 sky130_fd_sc_hd__or2_1 _3822_ (.A(net282),
    .B(_1454_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _3823_ (.A0(_1916_),
    .A1(_1917_),
    .S(_1289_),
    .X(_1455_));
 sky130_fd_sc_hd__nand2_1 _3824_ (.A(net278),
    .B(_1455_),
    .Y(_0288_));
 sky130_fd_sc_hd__mux2_1 _3825_ (.A0(\as1802.last_hi_addr[6] ),
    .A1(\as1802.addr_buff[14] ),
    .S(_1289_),
    .X(_1456_));
 sky130_fd_sc_hd__or2_1 _3826_ (.A(net282),
    .B(_1456_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _3827_ (.A0(_1914_),
    .A1(_1915_),
    .S(_1289_),
    .X(_1457_));
 sky130_fd_sc_hd__nand2_1 _3828_ (.A(net278),
    .B(_1457_),
    .Y(_0290_));
 sky130_fd_sc_hd__a41o_1 _3829_ (.A1(net273),
    .A2(\as1802.IE ),
    .A3(net12),
    .A4(net195),
    .B1(\as1802.will_interrupt ),
    .X(_1458_));
 sky130_fd_sc_hd__o211a_1 _3830_ (.A1(net193),
    .A2(_1203_),
    .B1(_1458_),
    .C1(net279),
    .X(_0291_));
 sky130_fd_sc_hd__a211o_1 _3831_ (.A1(net222),
    .A2(_1942_),
    .B1(_1993_),
    .C1(_2082_),
    .X(_1459_));
 sky130_fd_sc_hd__or3_2 _3832_ (.A(net272),
    .B(net176),
    .C(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__or4b_2 _3833_ (.A(_1206_),
    .B(_1211_),
    .C(_1216_),
    .D_N(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__and2b_1 _3834_ (.A_N(_1461_),
    .B(_1222_),
    .X(_1462_));
 sky130_fd_sc_hd__mux2_1 _3835_ (.A0(\as1802.IE ),
    .A1(_1278_),
    .S(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__or2_1 _3836_ (.A(net280),
    .B(_1463_),
    .X(_0292_));
 sky130_fd_sc_hd__nand2_1 _3837_ (.A(\as1802.IE ),
    .B(_1274_),
    .Y(_1464_));
 sky130_fd_sc_hd__o211a_1 _3838_ (.A1(\as1802.idle ),
    .A2(_1280_),
    .B1(_1464_),
    .C1(net279),
    .X(_0293_));
 sky130_fd_sc_hd__o21a_1 _3839_ (.A1(_1920_),
    .A2(net238),
    .B1(net15),
    .X(_1465_));
 sky130_fd_sc_hd__a211o_1 _3840_ (.A1(_1921_),
    .A2(\as1802.mem_write ),
    .B1(_1920_),
    .C1(net238),
    .X(_1466_));
 sky130_fd_sc_hd__or3b_1 _3841_ (.A(net281),
    .B(_1465_),
    .C_N(_1466_),
    .X(_0294_));
 sky130_fd_sc_hd__a21oi_1 _3842_ (.A1(net27),
    .A2(_1288_),
    .B1(net280),
    .Y(_1467_));
 sky130_fd_sc_hd__nand2_1 _3843_ (.A(_1447_),
    .B(_1467_),
    .Y(_0295_));
 sky130_fd_sc_hd__o21ai_1 _3844_ (.A1(\as1802.mem_cycle[2] ),
    .A2(_1285_),
    .B1(net29),
    .Y(_1468_));
 sky130_fd_sc_hd__a21oi_1 _3845_ (.A1(_1290_),
    .A2(_1468_),
    .B1(net281),
    .Y(_0296_));
 sky130_fd_sc_hd__and3_1 _3846_ (.A(net235),
    .B(_1926_),
    .C(net229),
    .X(_1469_));
 sky130_fd_sc_hd__or3b_1 _3847_ (.A(net173),
    .B(_2044_),
    .C_N(_1469_),
    .X(_1470_));
 sky130_fd_sc_hd__mux2_1 _3848_ (.A0(_1925_),
    .A1(_1913_),
    .S(_1470_),
    .X(_1471_));
 sky130_fd_sc_hd__nor2_1 _3849_ (.A(net281),
    .B(_1471_),
    .Y(_0297_));
 sky130_fd_sc_hd__o21a_1 _3850_ (.A1(net271),
    .A2(net158),
    .B1(_2067_),
    .X(_1472_));
 sky130_fd_sc_hd__and4b_1 _3851_ (.A_N(_1212_),
    .B(_1258_),
    .C(_1297_),
    .D(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__o32a_1 _3852_ (.A1(_1950_),
    .A2(net176),
    .A3(_1989_),
    .B1(_1941_),
    .B2(net220),
    .X(_1474_));
 sky130_fd_sc_hd__a21oi_1 _3853_ (.A1(_2022_),
    .A2(_1474_),
    .B1(net160),
    .Y(_1475_));
 sky130_fd_sc_hd__mux2_1 _3854_ (.A0(\as1802.lda ),
    .A1(_1475_),
    .S(_1473_),
    .X(_0298_));
 sky130_fd_sc_hd__nand2b_4 _3855_ (.A_N(net204),
    .B(net210),
    .Y(_1476_));
 sky130_fd_sc_hd__and2b_2 _3856_ (.A_N(net210),
    .B(net204),
    .X(_1477_));
 sky130_fd_sc_hd__nand2b_2 _3857_ (.A_N(net210),
    .B(net204),
    .Y(_1478_));
 sky130_fd_sc_hd__and2_2 _3858_ (.A(_1929_),
    .B(net205),
    .X(_1479_));
 sky130_fd_sc_hd__nand2_1 _3859_ (.A(_1929_),
    .B(net205),
    .Y(_1480_));
 sky130_fd_sc_hd__nor2_4 _3860_ (.A(_1929_),
    .B(net205),
    .Y(_1481_));
 sky130_fd_sc_hd__nand2b_4 _3861_ (.A_N(net212),
    .B(net35),
    .Y(_1482_));
 sky130_fd_sc_hd__nand2b_4 _3862_ (.A_N(net35),
    .B(net212),
    .Y(_1483_));
 sky130_fd_sc_hd__and2_2 _3863_ (.A(_1482_),
    .B(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__nand2_2 _3864_ (.A(_1482_),
    .B(_1483_),
    .Y(_1485_));
 sky130_fd_sc_hd__and2b_4 _3865_ (.A_N(net213),
    .B(net34),
    .X(_1486_));
 sky130_fd_sc_hd__and2b_4 _3866_ (.A_N(net34),
    .B(net213),
    .X(_1487_));
 sky130_fd_sc_hd__nor2_8 _3867_ (.A(_1486_),
    .B(_1487_),
    .Y(_1488_));
 sky130_fd_sc_hd__or2_4 _3868_ (.A(_1486_),
    .B(_1487_),
    .X(_1489_));
 sky130_fd_sc_hd__and2b_4 _3869_ (.A_N(net214),
    .B(net33),
    .X(_1490_));
 sky130_fd_sc_hd__nand2_4 _3870_ (.A(_1488_),
    .B(_1490_),
    .Y(_1491_));
 sky130_fd_sc_hd__and2b_4 _3871_ (.A_N(net33),
    .B(net214),
    .X(_1492_));
 sky130_fd_sc_hd__nor2_2 _3872_ (.A(_1490_),
    .B(_1492_),
    .Y(_1493_));
 sky130_fd_sc_hd__or2_4 _3873_ (.A(_1490_),
    .B(_1492_),
    .X(_1494_));
 sky130_fd_sc_hd__nand2b_4 _3874_ (.A_N(net215),
    .B(net206),
    .Y(_1495_));
 sky130_fd_sc_hd__nand2b_4 _3875_ (.A_N(net206),
    .B(net215),
    .Y(_1496_));
 sky130_fd_sc_hd__and2_1 _3876_ (.A(_1495_),
    .B(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__nand2_1 _3877_ (.A(_1495_),
    .B(_1496_),
    .Y(_1498_));
 sky130_fd_sc_hd__nand2b_2 _3878_ (.A_N(net216),
    .B(net207),
    .Y(_1499_));
 sky130_fd_sc_hd__and2b_1 _3879_ (.A_N(net209),
    .B(net218),
    .X(_1500_));
 sky130_fd_sc_hd__nand2b_4 _3880_ (.A_N(net207),
    .B(net216),
    .Y(_1501_));
 sky130_fd_sc_hd__and2_2 _3881_ (.A(_1499_),
    .B(_1501_),
    .X(_1502_));
 sky130_fd_sc_hd__xor2_4 _3882_ (.A(net216),
    .B(net207),
    .X(_1503_));
 sky130_fd_sc_hd__or2_2 _3883_ (.A(_1500_),
    .B(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__a21o_1 _3884_ (.A1(_1499_),
    .A2(_1504_),
    .B1(net180),
    .X(_1505_));
 sky130_fd_sc_hd__inv_2 _3885_ (.A(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__a21o_1 _3886_ (.A1(_1495_),
    .A2(_1505_),
    .B1(_1494_),
    .X(_1507_));
 sky130_fd_sc_hd__o21ai_2 _3887_ (.A1(_1489_),
    .A2(_1507_),
    .B1(_1491_),
    .Y(_1508_));
 sky130_fd_sc_hd__o21ai_2 _3888_ (.A1(_1486_),
    .A2(_1508_),
    .B1(net182),
    .Y(_1509_));
 sky130_fd_sc_hd__and2_1 _3889_ (.A(_1482_),
    .B(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__a21oi_2 _3890_ (.A1(_1480_),
    .A2(_1510_),
    .B1(_1481_),
    .Y(_1511_));
 sky130_fd_sc_hd__a21o_1 _3891_ (.A1(_1476_),
    .A2(_1511_),
    .B1(_1477_),
    .X(_1512_));
 sky130_fd_sc_hd__and2b_1 _3892_ (.A_N(net218),
    .B(net209),
    .X(_1513_));
 sky130_fd_sc_hd__or2_2 _3893_ (.A(_1503_),
    .B(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__or3_1 _3894_ (.A(_1485_),
    .B(_1500_),
    .C(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__and2_4 _3895_ (.A(_1476_),
    .B(_1478_),
    .X(_1516_));
 sky130_fd_sc_hd__nand2_2 _3896_ (.A(_1476_),
    .B(_1478_),
    .Y(_1517_));
 sky130_fd_sc_hd__nor2_4 _3897_ (.A(_1479_),
    .B(_1481_),
    .Y(_1518_));
 sky130_fd_sc_hd__or2_4 _3898_ (.A(_1479_),
    .B(_1481_),
    .X(_1519_));
 sky130_fd_sc_hd__or4_2 _3899_ (.A(_1489_),
    .B(net181),
    .C(net180),
    .D(_1515_),
    .X(_1520_));
 sky130_fd_sc_hd__o31a_1 _3900_ (.A1(_1517_),
    .A2(_1519_),
    .A3(_1520_),
    .B1(_1512_),
    .X(_1521_));
 sky130_fd_sc_hd__a2bb2o_1 _3901_ (.A1_N(_1980_),
    .A2_N(_1521_),
    .B1(_1512_),
    .B2(_1981_),
    .X(_1522_));
 sky130_fd_sc_hd__nand2_2 _3902_ (.A(_1481_),
    .B(_1516_),
    .Y(_1523_));
 sky130_fd_sc_hd__or2_2 _3903_ (.A(_1481_),
    .B(_1516_),
    .X(_1524_));
 sky130_fd_sc_hd__nor2_4 _3904_ (.A(_1483_),
    .B(_1519_),
    .Y(_1525_));
 sky130_fd_sc_hd__and2_2 _3905_ (.A(_1483_),
    .B(_1519_),
    .X(_1526_));
 sky130_fd_sc_hd__nand2_2 _3906_ (.A(net182),
    .B(_1487_),
    .Y(_1527_));
 sky130_fd_sc_hd__or2_1 _3907_ (.A(net182),
    .B(_1487_),
    .X(_1528_));
 sky130_fd_sc_hd__nand2_1 _3908_ (.A(_1527_),
    .B(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__nand2_4 _3909_ (.A(_1488_),
    .B(_1492_),
    .Y(_1530_));
 sky130_fd_sc_hd__or2_2 _3910_ (.A(_1488_),
    .B(_1492_),
    .X(_1531_));
 sky130_fd_sc_hd__nor2_2 _3911_ (.A(net181),
    .B(_1496_),
    .Y(_1532_));
 sky130_fd_sc_hd__or2_1 _3912_ (.A(net181),
    .B(_1496_),
    .X(_1533_));
 sky130_fd_sc_hd__nand2_1 _3913_ (.A(net181),
    .B(_1496_),
    .Y(_1534_));
 sky130_fd_sc_hd__nor2_1 _3914_ (.A(net207),
    .B(net179),
    .Y(_1535_));
 sky130_fd_sc_hd__and2_1 _3915_ (.A(net207),
    .B(net179),
    .X(_1536_));
 sky130_fd_sc_hd__nor2_1 _3916_ (.A(_1535_),
    .B(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__nand2_2 _3917_ (.A(net217),
    .B(net207),
    .Y(_1538_));
 sky130_fd_sc_hd__o21bai_2 _3918_ (.A1(_1911_),
    .A2(_1513_),
    .B1_N(_1500_),
    .Y(_1539_));
 sky130_fd_sc_hd__o21ai_1 _3919_ (.A1(net216),
    .A2(net207),
    .B1(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__nand2_1 _3920_ (.A(_1538_),
    .B(_1540_),
    .Y(_1541_));
 sky130_fd_sc_hd__and2_1 _3921_ (.A(_1537_),
    .B(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__o211a_2 _3922_ (.A1(_1535_),
    .A2(_1542_),
    .B1(_1533_),
    .C1(_1534_),
    .X(_1543_));
 sky130_fd_sc_hd__o211ai_4 _3923_ (.A1(_1532_),
    .A2(_1543_),
    .B1(_1530_),
    .C1(_1531_),
    .Y(_1544_));
 sky130_fd_sc_hd__a21o_2 _3924_ (.A1(_1530_),
    .A2(_1544_),
    .B1(_1529_),
    .X(_1545_));
 sky130_fd_sc_hd__a211oi_4 _3925_ (.A1(_1527_),
    .A2(_1545_),
    .B1(_1525_),
    .C1(_1526_),
    .Y(_1546_));
 sky130_fd_sc_hd__o211a_1 _3926_ (.A1(_1525_),
    .A2(_1546_),
    .B1(_1523_),
    .C1(_1524_),
    .X(_1547_));
 sky130_fd_sc_hd__nor2_4 _3927_ (.A(net230),
    .B(_1980_),
    .Y(_1548_));
 sky130_fd_sc_hd__o211ai_1 _3928_ (.A1(_1476_),
    .A2(_1547_),
    .B1(_1548_),
    .C1(_1523_),
    .Y(_1549_));
 sky130_fd_sc_hd__a21oi_1 _3929_ (.A1(_1476_),
    .A2(_1547_),
    .B1(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__nor2_2 _3930_ (.A(net229),
    .B(_1983_),
    .Y(_1551_));
 sky130_fd_sc_hd__nor2_2 _3931_ (.A(_1964_),
    .B(_2005_),
    .Y(_1552_));
 sky130_fd_sc_hd__a22o_1 _3932_ (.A1(net219),
    .A2(net157),
    .B1(net178),
    .B2(net210),
    .X(_1553_));
 sky130_fd_sc_hd__nand2_2 _3933_ (.A(\as1802.D[6] ),
    .B(net205),
    .Y(_1554_));
 sky130_fd_sc_hd__nand2_2 _3934_ (.A(net212),
    .B(net35),
    .Y(_1555_));
 sky130_fd_sc_hd__nand2_2 _3935_ (.A(net213),
    .B(net34),
    .Y(_1556_));
 sky130_fd_sc_hd__nand2_2 _3936_ (.A(net214),
    .B(net33),
    .Y(_1557_));
 sky130_fd_sc_hd__and2_1 _3937_ (.A(net215),
    .B(net206),
    .X(_1558_));
 sky130_fd_sc_hd__nand2_2 _3938_ (.A(net215),
    .B(net206),
    .Y(_1559_));
 sky130_fd_sc_hd__nand2_2 _3939_ (.A(net218),
    .B(net209),
    .Y(_1560_));
 sky130_fd_sc_hd__or2_2 _3940_ (.A(_1502_),
    .B(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__or2_1 _3941_ (.A(net218),
    .B(net209),
    .X(_1562_));
 sky130_fd_sc_hd__a21bo_1 _3942_ (.A1(\as1802.DF ),
    .A2(_1562_),
    .B1_N(_1560_),
    .X(_1563_));
 sky130_fd_sc_hd__a21bo_1 _3943_ (.A1(_1503_),
    .A2(_1563_),
    .B1_N(_1538_),
    .X(_1564_));
 sky130_fd_sc_hd__nand2_1 _3944_ (.A(net179),
    .B(_1564_),
    .Y(_1565_));
 sky130_fd_sc_hd__a21o_1 _3945_ (.A1(_1559_),
    .A2(_1565_),
    .B1(_1493_),
    .X(_1566_));
 sky130_fd_sc_hd__a21o_1 _3946_ (.A1(_1557_),
    .A2(_1566_),
    .B1(_1488_),
    .X(_1567_));
 sky130_fd_sc_hd__a21o_1 _3947_ (.A1(_1556_),
    .A2(_1567_),
    .B1(net182),
    .X(_1568_));
 sky130_fd_sc_hd__a21o_1 _3948_ (.A1(_1555_),
    .A2(_1568_),
    .B1(_1518_),
    .X(_1569_));
 sky130_fd_sc_hd__a21oi_2 _3949_ (.A1(_1554_),
    .A2(_1569_),
    .B1(_1516_),
    .Y(_1570_));
 sky130_fd_sc_hd__a21o_1 _3950_ (.A1(net211),
    .A2(net204),
    .B1(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__nor2_1 _3951_ (.A(_1480_),
    .B(_1517_),
    .Y(_1572_));
 sky130_fd_sc_hd__nor2_1 _3952_ (.A(_1479_),
    .B(_1516_),
    .Y(_1573_));
 sky130_fd_sc_hd__or2_1 _3953_ (.A(_1572_),
    .B(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__nor2_1 _3954_ (.A(_1482_),
    .B(_1519_),
    .Y(_1575_));
 sky130_fd_sc_hd__or2_1 _3955_ (.A(_1482_),
    .B(_1519_),
    .X(_1576_));
 sky130_fd_sc_hd__and2_2 _3956_ (.A(_1482_),
    .B(_1519_),
    .X(_1577_));
 sky130_fd_sc_hd__nand2_2 _3957_ (.A(_1484_),
    .B(_1486_),
    .Y(_1578_));
 sky130_fd_sc_hd__inv_2 _3958_ (.A(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__nor2_1 _3959_ (.A(_1484_),
    .B(_1486_),
    .Y(_1580_));
 sky130_fd_sc_hd__or2_4 _3960_ (.A(_1488_),
    .B(_1490_),
    .X(_1581_));
 sky130_fd_sc_hd__inv_2 _3961_ (.A(_1581_),
    .Y(_1582_));
 sky130_fd_sc_hd__nor2_8 _3962_ (.A(net181),
    .B(_1495_),
    .Y(_1583_));
 sky130_fd_sc_hd__and2_2 _3963_ (.A(net181),
    .B(_1495_),
    .X(_1584_));
 sky130_fd_sc_hd__nand2_1 _3964_ (.A(_1494_),
    .B(_1495_),
    .Y(_1585_));
 sky130_fd_sc_hd__or2_2 _3965_ (.A(net216),
    .B(net179),
    .X(_1586_));
 sky130_fd_sc_hd__xnor2_2 _3966_ (.A(\as1802.DF ),
    .B(net219),
    .Y(_1587_));
 sky130_fd_sc_hd__nand2_2 _3967_ (.A(net209),
    .B(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__o21ai_4 _3968_ (.A1(_1911_),
    .A2(net218),
    .B1(_1588_),
    .Y(_1589_));
 sky130_fd_sc_hd__xor2_1 _3969_ (.A(net216),
    .B(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__and2_1 _3970_ (.A(net207),
    .B(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__a21o_1 _3971_ (.A1(net216),
    .A2(_1589_),
    .B1(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__nand2_1 _3972_ (.A(net216),
    .B(net179),
    .Y(_1593_));
 sky130_fd_sc_hd__and2_1 _3973_ (.A(_1586_),
    .B(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__nand2_2 _3974_ (.A(_1592_),
    .B(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__a211oi_4 _3975_ (.A1(_1586_),
    .A2(_1595_),
    .B1(_1583_),
    .C1(_1584_),
    .Y(_1596_));
 sky130_fd_sc_hd__o211ai_4 _3976_ (.A1(_1583_),
    .A2(_1596_),
    .B1(_1491_),
    .C1(_1581_),
    .Y(_1597_));
 sky130_fd_sc_hd__a211o_1 _3977_ (.A1(_1491_),
    .A2(_1597_),
    .B1(_1580_),
    .C1(_1579_),
    .X(_1598_));
 sky130_fd_sc_hd__a211o_1 _3978_ (.A1(_1578_),
    .A2(_1598_),
    .B1(_1575_),
    .C1(_1577_),
    .X(_1599_));
 sky130_fd_sc_hd__a21o_1 _3979_ (.A1(_1576_),
    .A2(_1599_),
    .B1(_1574_),
    .X(_1600_));
 sky130_fd_sc_hd__nor2_1 _3980_ (.A(_1477_),
    .B(_1572_),
    .Y(_1601_));
 sky130_fd_sc_hd__o21a_2 _3981_ (.A1(net230),
    .A2(_1976_),
    .B1(net231),
    .X(_1602_));
 sky130_fd_sc_hd__o21ai_4 _3982_ (.A1(net230),
    .A2(_1976_),
    .B1(net231),
    .Y(_1603_));
 sky130_fd_sc_hd__mux2_1 _3983_ (.A0(_1477_),
    .A1(_1601_),
    .S(_1600_),
    .X(_1604_));
 sky130_fd_sc_hd__a22o_1 _3984_ (.A1(net230),
    .A2(_1522_),
    .B1(_1571_),
    .B2(_1954_),
    .X(_1605_));
 sky130_fd_sc_hd__or4_1 _3985_ (.A(_1550_),
    .B(_1553_),
    .C(_1603_),
    .D(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__o211a_1 _3986_ (.A1(_1602_),
    .A2(_1604_),
    .B1(_1606_),
    .C1(net175),
    .X(_1607_));
 sky130_fd_sc_hd__nand2_1 _3987_ (.A(_2022_),
    .B(_2026_),
    .Y(_1608_));
 sky130_fd_sc_hd__and3_1 _3988_ (.A(\as1802.instr_latch[5] ),
    .B(_2018_),
    .C(_1291_),
    .X(_1609_));
 sky130_fd_sc_hd__or4b_1 _3989_ (.A(net192),
    .B(net137),
    .C(_1609_),
    .D_N(_2025_),
    .X(_1610_));
 sky130_fd_sc_hd__or4_1 _3990_ (.A(_1999_),
    .B(_1220_),
    .C(_1459_),
    .D(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__nand2_1 _3991_ (.A(net173),
    .B(_2018_),
    .Y(_1612_));
 sky130_fd_sc_hd__a221o_1 _3992_ (.A1(_1926_),
    .A2(_1608_),
    .B1(_1612_),
    .B2(_2022_),
    .C1(_1611_),
    .X(_1613_));
 sky130_fd_sc_hd__or4_1 _3993_ (.A(net202),
    .B(_1952_),
    .C(_1522_),
    .D(_1553_),
    .X(_1614_));
 sky130_fd_sc_hd__a21oi_2 _3994_ (.A1(_1538_),
    .A2(_1561_),
    .B1(_1497_),
    .Y(_1615_));
 sky130_fd_sc_hd__o21ai_2 _3995_ (.A1(_1558_),
    .A2(_1615_),
    .B1(net181),
    .Y(_1616_));
 sky130_fd_sc_hd__a21o_1 _3996_ (.A1(_1557_),
    .A2(_1616_),
    .B1(_1488_),
    .X(_1617_));
 sky130_fd_sc_hd__a21o_1 _3997_ (.A1(_1556_),
    .A2(_1617_),
    .B1(net182),
    .X(_1618_));
 sky130_fd_sc_hd__a21o_1 _3998_ (.A1(_1555_),
    .A2(_1618_),
    .B1(_1518_),
    .X(_1619_));
 sky130_fd_sc_hd__a21oi_2 _3999_ (.A1(_1554_),
    .A2(_1619_),
    .B1(_1516_),
    .Y(_1620_));
 sky130_fd_sc_hd__a221o_1 _4000_ (.A1(net210),
    .A2(net204),
    .B1(_1953_),
    .B2(net232),
    .C1(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__a311oi_1 _4001_ (.A1(net173),
    .A2(_1614_),
    .A3(_1621_),
    .B1(_1607_),
    .C1(_1613_),
    .Y(_1622_));
 sky130_fd_sc_hd__a211oi_1 _4002_ (.A1(_1911_),
    .A2(_1613_),
    .B1(_1622_),
    .C1(net281),
    .Y(_0299_));
 sky130_fd_sc_hd__or3b_1 _4003_ (.A(_1949_),
    .B(net274),
    .C_N(\as1802.instr_latch[4] ),
    .X(_1623_));
 sky130_fd_sc_hd__o211a_4 _4004_ (.A1(_2092_),
    .A2(_1222_),
    .B1(_1623_),
    .C1(_1217_),
    .X(_1624_));
 sky130_fd_sc_hd__mux2_1 _4005_ (.A0(\as1802.P[0] ),
    .A1(net34),
    .S(net167),
    .X(_1625_));
 sky130_fd_sc_hd__mux2_1 _4006_ (.A0(net237),
    .A1(_1625_),
    .S(net175),
    .X(_1626_));
 sky130_fd_sc_hd__a21bo_1 _4007_ (.A1(net203),
    .A2(_1626_),
    .B1_N(_1624_),
    .X(_1627_));
 sky130_fd_sc_hd__o211a_1 _4008_ (.A1(\as1802.X[0] ),
    .A2(_1624_),
    .B1(_1627_),
    .C1(net277),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _4009_ (.A0(\as1802.P[1] ),
    .A1(net35),
    .S(net167),
    .X(_1628_));
 sky130_fd_sc_hd__nand2_1 _4010_ (.A(net175),
    .B(_1628_),
    .Y(_1629_));
 sky130_fd_sc_hd__nand4_1 _4011_ (.A(net203),
    .B(_1226_),
    .C(_1624_),
    .D(_1629_),
    .Y(_1630_));
 sky130_fd_sc_hd__o211a_1 _4012_ (.A1(\as1802.X[1] ),
    .A2(_1624_),
    .B1(_1630_),
    .C1(net277),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _4013_ (.A0(\as1802.P[2] ),
    .A1(net205),
    .S(net167),
    .X(_1631_));
 sky130_fd_sc_hd__o21a_1 _4014_ (.A1(net170),
    .A2(_1631_),
    .B1(_1229_),
    .X(_1632_));
 sky130_fd_sc_hd__mux2_1 _4015_ (.A0(\as1802.X[2] ),
    .A1(_1632_),
    .S(_1624_),
    .X(_1633_));
 sky130_fd_sc_hd__and2_1 _4016_ (.A(net277),
    .B(_1633_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_2 _4017_ (.A0(\as1802.P[3] ),
    .A1(net204),
    .S(net168),
    .X(_1634_));
 sky130_fd_sc_hd__o21a_1 _4018_ (.A1(net170),
    .A2(_1634_),
    .B1(_1232_),
    .X(_1635_));
 sky130_fd_sc_hd__mux2_1 _4019_ (.A0(\as1802.X[3] ),
    .A1(_1635_),
    .S(_1624_),
    .X(_1636_));
 sky130_fd_sc_hd__and2_1 _4020_ (.A(net277),
    .B(_1636_),
    .X(_0303_));
 sky130_fd_sc_hd__a211o_4 _4021_ (.A1(net168),
    .A2(_1221_),
    .B1(_1461_),
    .C1(_1213_),
    .X(_1637_));
 sky130_fd_sc_hd__mux2_1 _4022_ (.A0(\as1802.P[0] ),
    .A1(\as1802.T[0] ),
    .S(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__and2_1 _4023_ (.A(net276),
    .B(_1638_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _4024_ (.A0(\as1802.P[1] ),
    .A1(\as1802.T[1] ),
    .S(_1637_),
    .X(_1639_));
 sky130_fd_sc_hd__and2_1 _4025_ (.A(net276),
    .B(_1639_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _4026_ (.A0(\as1802.P[2] ),
    .A1(\as1802.T[2] ),
    .S(_1637_),
    .X(_1640_));
 sky130_fd_sc_hd__and2_1 _4027_ (.A(net276),
    .B(_1640_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _4028_ (.A0(\as1802.P[3] ),
    .A1(\as1802.T[3] ),
    .S(_1637_),
    .X(_1641_));
 sky130_fd_sc_hd__and2_1 _4029_ (.A(net276),
    .B(_1641_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _4030_ (.A0(\as1802.X[0] ),
    .A1(\as1802.T[4] ),
    .S(_1637_),
    .X(_1642_));
 sky130_fd_sc_hd__and2_1 _4031_ (.A(net276),
    .B(_1642_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _4032_ (.A0(\as1802.X[1] ),
    .A1(\as1802.T[5] ),
    .S(_1637_),
    .X(_1643_));
 sky130_fd_sc_hd__and2_1 _4033_ (.A(net276),
    .B(_1643_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _4034_ (.A0(\as1802.X[2] ),
    .A1(\as1802.T[6] ),
    .S(_1637_),
    .X(_1644_));
 sky130_fd_sc_hd__and2_1 _4035_ (.A(net276),
    .B(_1644_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _4036_ (.A0(\as1802.X[3] ),
    .A1(\as1802.T[7] ),
    .S(_1637_),
    .X(_1645_));
 sky130_fd_sc_hd__and2_1 _4037_ (.A(net276),
    .B(_1645_),
    .X(_0311_));
 sky130_fd_sc_hd__a21oi_1 _4038_ (.A1(net201),
    .A2(_1944_),
    .B1(_1988_),
    .Y(_1646_));
 sky130_fd_sc_hd__o32a_1 _4039_ (.A1(_2023_),
    .A2(_2098_),
    .A3(_1646_),
    .B1(_2022_),
    .B2(net232),
    .X(_1647_));
 sky130_fd_sc_hd__or2_1 _4040_ (.A(net272),
    .B(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__a31o_1 _4041_ (.A1(_2043_),
    .A2(_1210_),
    .A3(_1648_),
    .B1(net193),
    .X(_1649_));
 sky130_fd_sc_hd__or3_2 _4042_ (.A(net269),
    .B(\as1802.mem_write ),
    .C(_1447_),
    .X(_1650_));
 sky130_fd_sc_hd__a2bb2o_1 _4043_ (.A1_N(net238),
    .A2_N(_1275_),
    .B1(net279),
    .B2(_1920_),
    .X(_1651_));
 sky130_fd_sc_hd__o21a_1 _4044_ (.A1(\as1802.mem_cycle[1] ),
    .A2(\as1802.mem_cycle[0] ),
    .B1(\as1802.mem_cycle[2] ),
    .X(_1652_));
 sky130_fd_sc_hd__o211a_1 _4045_ (.A1(net196),
    .A2(_1652_),
    .B1(_1651_),
    .C1(_1277_),
    .X(_1653_));
 sky130_fd_sc_hd__nand2_1 _4046_ (.A(_1936_),
    .B(_1940_),
    .Y(_1654_));
 sky130_fd_sc_hd__a31o_1 _4047_ (.A1(net203),
    .A2(_2016_),
    .A3(_1654_),
    .B1(net193),
    .X(_1655_));
 sky130_fd_sc_hd__o211a_1 _4048_ (.A1(_2044_),
    .A2(_1218_),
    .B1(_1448_),
    .C1(_1655_),
    .X(_1656_));
 sky130_fd_sc_hd__o22a_1 _4049_ (.A1(net273),
    .A2(net158),
    .B1(_1220_),
    .B2(_2000_),
    .X(_1657_));
 sky130_fd_sc_hd__or3_1 _4050_ (.A(net272),
    .B(_2023_),
    .C(_2099_),
    .X(_1658_));
 sky130_fd_sc_hd__o32a_1 _4051_ (.A1(net192),
    .A2(_1943_),
    .A3(_1658_),
    .B1(_2050_),
    .B2(_1966_),
    .X(_1659_));
 sky130_fd_sc_hd__o211a_1 _4052_ (.A1(\as1802.lda ),
    .A2(_1650_),
    .B1(_1656_),
    .C1(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__o211a_1 _4053_ (.A1(_1946_),
    .A2(_1657_),
    .B1(_1660_),
    .C1(_1653_),
    .X(_1661_));
 sky130_fd_sc_hd__and3b_4 _4054_ (.A_N(_1282_),
    .B(_1649_),
    .C(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__a32o_1 _4055_ (.A1(net218),
    .A2(net209),
    .A3(_1256_),
    .B1(net157),
    .B2(net217),
    .X(_1663_));
 sky130_fd_sc_hd__nor2_4 _4056_ (.A(net236),
    .B(net233),
    .Y(_1664_));
 sky130_fd_sc_hd__or2_4 _4057_ (.A(net236),
    .B(net234),
    .X(_1665_));
 sky130_fd_sc_hd__o211a_1 _4058_ (.A1(_1560_),
    .A2(_1664_),
    .B1(_1562_),
    .C1(_1964_),
    .X(_1666_));
 sky130_fd_sc_hd__or3_1 _4059_ (.A(_2035_),
    .B(_1663_),
    .C(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__o211a_1 _4060_ (.A1(net191),
    .A2(_0780_),
    .B1(_1667_),
    .C1(net185),
    .X(_1668_));
 sky130_fd_sc_hd__nor2_1 _4061_ (.A(net185),
    .B(net82),
    .Y(_1669_));
 sky130_fd_sc_hd__and2_4 _4062_ (.A(net195),
    .B(_2023_),
    .X(_1670_));
 sky130_fd_sc_hd__xnor2_1 _4063_ (.A(net209),
    .B(_1587_),
    .Y(_1671_));
 sky130_fd_sc_hd__a21oi_1 _4064_ (.A1(_1925_),
    .A2(net233),
    .B1(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__a221o_1 _4065_ (.A1(net217),
    .A2(_1551_),
    .B1(_1671_),
    .B2(net188),
    .C1(net172),
    .X(_1673_));
 sky130_fd_sc_hd__a211o_1 _4066_ (.A1(\as1802.DF ),
    .A2(_1552_),
    .B1(_1672_),
    .C1(_1673_),
    .X(_1674_));
 sky130_fd_sc_hd__o311a_1 _4067_ (.A1(net175),
    .A2(_1668_),
    .A3(_1669_),
    .B1(_1670_),
    .C1(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__a21bo_1 _4068_ (.A1(net1),
    .A2(net194),
    .B1_N(_1662_),
    .X(_1676_));
 sky130_fd_sc_hd__o22a_1 _4069_ (.A1(net218),
    .A2(_1662_),
    .B1(_1675_),
    .B2(_1676_),
    .X(_0312_));
 sky130_fd_sc_hd__a22o_1 _4070_ (.A1(net215),
    .A2(net157),
    .B1(net178),
    .B2(net218),
    .X(_1677_));
 sky130_fd_sc_hd__o21a_1 _4071_ (.A1(net217),
    .A2(net208),
    .B1(_1664_),
    .X(_1678_));
 sky130_fd_sc_hd__nand2_1 _4072_ (.A(_1500_),
    .B(_1503_),
    .Y(_1679_));
 sky130_fd_sc_hd__nand2_1 _4073_ (.A(_1502_),
    .B(_1560_),
    .Y(_1680_));
 sky130_fd_sc_hd__nand2_1 _4074_ (.A(_1503_),
    .B(_1513_),
    .Y(_1681_));
 sky130_fd_sc_hd__a31o_1 _4075_ (.A1(net188),
    .A2(_1561_),
    .A3(_1680_),
    .B1(_1677_),
    .X(_1682_));
 sky130_fd_sc_hd__a31o_1 _4076_ (.A1(_1979_),
    .A2(_1514_),
    .A3(_1681_),
    .B1(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__a311oi_2 _4077_ (.A1(_1981_),
    .A2(_1504_),
    .A3(_1679_),
    .B1(_1683_),
    .C1(_1678_),
    .Y(_1684_));
 sky130_fd_sc_hd__o221a_1 _4078_ (.A1(_1986_),
    .A2(_1502_),
    .B1(_1538_),
    .B2(_1257_),
    .C1(_1684_),
    .X(_1685_));
 sky130_fd_sc_hd__mux2_1 _4079_ (.A0(_0837_),
    .A1(_1685_),
    .S(net191),
    .X(_1686_));
 sky130_fd_sc_hd__mux2_1 _4080_ (.A0(_0398_),
    .A1(_1686_),
    .S(net185),
    .X(_1687_));
 sky130_fd_sc_hd__nand2_1 _4081_ (.A(net170),
    .B(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__nor2_1 _4082_ (.A(net207),
    .B(_1590_),
    .Y(_1689_));
 sky130_fd_sc_hd__or2_1 _4083_ (.A(_1591_),
    .B(_1689_),
    .X(_1690_));
 sky130_fd_sc_hd__nor2_1 _4084_ (.A(_1602_),
    .B(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__nor2_2 _4085_ (.A(_1976_),
    .B(_2005_),
    .Y(_1692_));
 sky130_fd_sc_hd__or2_2 _4086_ (.A(_1976_),
    .B(_2005_),
    .X(_1693_));
 sky130_fd_sc_hd__nand2_1 _4087_ (.A(_1502_),
    .B(_1539_),
    .Y(_1694_));
 sky130_fd_sc_hd__or2_1 _4088_ (.A(_1502_),
    .B(_1539_),
    .X(_1695_));
 sky130_fd_sc_hd__and2_1 _4089_ (.A(_1694_),
    .B(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__nor2_2 _4090_ (.A(_1974_),
    .B(_2005_),
    .Y(_1697_));
 sky130_fd_sc_hd__or2_2 _4091_ (.A(_1974_),
    .B(_2005_),
    .X(_1698_));
 sky130_fd_sc_hd__xnor2_1 _4092_ (.A(_1502_),
    .B(_1563_),
    .Y(_1699_));
 sky130_fd_sc_hd__mux2_1 _4093_ (.A0(_1548_),
    .A1(_1697_),
    .S(_1696_),
    .X(_1700_));
 sky130_fd_sc_hd__a221o_1 _4094_ (.A1(_1690_),
    .A2(_1692_),
    .B1(_1699_),
    .B2(net188),
    .C1(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__or4_1 _4095_ (.A(net172),
    .B(_1677_),
    .C(_1691_),
    .D(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__a32o_1 _4096_ (.A1(_1670_),
    .A2(_1688_),
    .A3(_1702_),
    .B1(net194),
    .B2(net5),
    .X(_1703_));
 sky130_fd_sc_hd__mux2_1 _4097_ (.A0(net216),
    .A1(_1703_),
    .S(_1662_),
    .X(_0313_));
 sky130_fd_sc_hd__a21o_1 _4098_ (.A1(_1501_),
    .A2(_1514_),
    .B1(net180),
    .X(_1704_));
 sky130_fd_sc_hd__a31o_1 _4099_ (.A1(net180),
    .A2(_1501_),
    .A3(_1514_),
    .B1(_1980_),
    .X(_1705_));
 sky130_fd_sc_hd__and2b_1 _4100_ (.A_N(_1705_),
    .B(_1704_),
    .X(_1706_));
 sky130_fd_sc_hd__a22o_1 _4101_ (.A1(net214),
    .A2(net157),
    .B1(net178),
    .B2(net216),
    .X(_1707_));
 sky130_fd_sc_hd__o221a_1 _4102_ (.A1(_1986_),
    .A2(_1497_),
    .B1(_1559_),
    .B2(_1257_),
    .C1(_1665_),
    .X(_1708_));
 sky130_fd_sc_hd__and3_1 _4103_ (.A(_1497_),
    .B(_1538_),
    .C(_1561_),
    .X(_1709_));
 sky130_fd_sc_hd__nand2_1 _4104_ (.A(_1981_),
    .B(_1505_),
    .Y(_1710_));
 sky130_fd_sc_hd__a31o_1 _4105_ (.A1(net180),
    .A2(_1499_),
    .A3(_1504_),
    .B1(_1710_),
    .X(_1711_));
 sky130_fd_sc_hd__o31a_1 _4106_ (.A1(_1955_),
    .A2(_1615_),
    .A3(_1709_),
    .B1(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__or4bb_1 _4107_ (.A(_1706_),
    .B(_1707_),
    .C_N(_1708_),
    .D_N(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__o31a_1 _4108_ (.A1(net215),
    .A2(net206),
    .A3(_1665_),
    .B1(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__o21ai_1 _4109_ (.A1(_2035_),
    .A2(_1714_),
    .B1(net185),
    .Y(_1715_));
 sky130_fd_sc_hd__a21o_1 _4110_ (.A1(_2035_),
    .A2(_0891_),
    .B1(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__o211ai_4 _4111_ (.A1(net185),
    .A2(_0445_),
    .B1(_1716_),
    .C1(net171),
    .Y(_1717_));
 sky130_fd_sc_hd__or2_1 _4112_ (.A(_1592_),
    .B(_1594_),
    .X(_1718_));
 sky130_fd_sc_hd__or2_1 _4113_ (.A(net179),
    .B(_1564_),
    .X(_1719_));
 sky130_fd_sc_hd__and3_1 _4114_ (.A(net188),
    .B(_1565_),
    .C(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__a21o_1 _4115_ (.A1(_1501_),
    .A2(_1694_),
    .B1(net179),
    .X(_1721_));
 sky130_fd_sc_hd__and3_1 _4116_ (.A(net179),
    .B(_1501_),
    .C(_1694_),
    .X(_1722_));
 sky130_fd_sc_hd__or3b_1 _4117_ (.A(_1722_),
    .B(_1698_),
    .C_N(_1721_),
    .X(_1723_));
 sky130_fd_sc_hd__o21ai_1 _4118_ (.A1(_1537_),
    .A2(_1541_),
    .B1(_1548_),
    .Y(_1724_));
 sky130_fd_sc_hd__nand2_1 _4119_ (.A(_1501_),
    .B(_1589_),
    .Y(_1725_));
 sky130_fd_sc_hd__a21oi_2 _4120_ (.A1(_1499_),
    .A2(_1725_),
    .B1(net179),
    .Y(_1726_));
 sky130_fd_sc_hd__a311o_1 _4121_ (.A1(net179),
    .A2(_1499_),
    .A3(_1725_),
    .B1(_1726_),
    .C1(_1693_),
    .X(_1727_));
 sky130_fd_sc_hd__o211a_1 _4122_ (.A1(_1542_),
    .A2(_1724_),
    .B1(_1727_),
    .C1(_1723_),
    .X(_1728_));
 sky130_fd_sc_hd__or4b_1 _4123_ (.A(net172),
    .B(_1707_),
    .C(_1720_),
    .D_N(_1728_),
    .X(_1729_));
 sky130_fd_sc_hd__a31o_1 _4124_ (.A1(_1595_),
    .A2(_1603_),
    .A3(_1718_),
    .B1(_1729_),
    .X(_1730_));
 sky130_fd_sc_hd__a32o_1 _4125_ (.A1(_1670_),
    .A2(_1717_),
    .A3(_1730_),
    .B1(net194),
    .B2(net6),
    .X(_1731_));
 sky130_fd_sc_hd__mux2_1 _4126_ (.A0(net215),
    .A1(_1731_),
    .S(_1662_),
    .X(_0314_));
 sky130_fd_sc_hd__or3_1 _4127_ (.A(net181),
    .B(_1558_),
    .C(_1615_),
    .X(_1732_));
 sky130_fd_sc_hd__and3_1 _4128_ (.A(net188),
    .B(_1616_),
    .C(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__o211a_1 _4129_ (.A1(_1506_),
    .A2(_1585_),
    .B1(_1507_),
    .C1(_1981_),
    .X(_1734_));
 sky130_fd_sc_hd__a2bb2o_1 _4130_ (.A1_N(_1257_),
    .A2_N(_1557_),
    .B1(net181),
    .B2(_1987_),
    .X(_1735_));
 sky130_fd_sc_hd__a221o_1 _4131_ (.A1(net213),
    .A2(net157),
    .B1(net178),
    .B2(\as1802.D[2] ),
    .C1(_1664_),
    .X(_1736_));
 sky130_fd_sc_hd__nand2_1 _4132_ (.A(_1496_),
    .B(_1704_),
    .Y(_1737_));
 sky130_fd_sc_hd__a31o_1 _4133_ (.A1(net181),
    .A2(_1496_),
    .A3(_1704_),
    .B1(_1980_),
    .X(_1738_));
 sky130_fd_sc_hd__a21o_1 _4134_ (.A1(_1493_),
    .A2(_1737_),
    .B1(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__or4b_1 _4135_ (.A(_1734_),
    .B(_1735_),
    .C(_1736_),
    .D_N(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__o32a_1 _4136_ (.A1(net214),
    .A2(net33),
    .A3(_1665_),
    .B1(_1733_),
    .B2(_1740_),
    .X(_1741_));
 sky130_fd_sc_hd__o21a_1 _4137_ (.A1(_2035_),
    .A2(_1741_),
    .B1(net185),
    .X(_1742_));
 sky130_fd_sc_hd__o21ai_2 _4138_ (.A1(net191),
    .A2(_0963_),
    .B1(_1742_),
    .Y(_1743_));
 sky130_fd_sc_hd__a21o_1 _4139_ (.A1(_1493_),
    .A2(_1726_),
    .B1(_1583_),
    .X(_1744_));
 sky130_fd_sc_hd__nor2_1 _4140_ (.A(_1585_),
    .B(_1726_),
    .Y(_1745_));
 sky130_fd_sc_hd__a21oi_2 _4141_ (.A1(_1496_),
    .A2(_1721_),
    .B1(_1494_),
    .Y(_1746_));
 sky130_fd_sc_hd__a31o_1 _4142_ (.A1(_1494_),
    .A2(_1496_),
    .A3(_1721_),
    .B1(_1698_),
    .X(_1747_));
 sky130_fd_sc_hd__a221o_1 _4143_ (.A1(net213),
    .A2(net157),
    .B1(net178),
    .B2(\as1802.D[2] ),
    .C1(_1603_),
    .X(_1748_));
 sky130_fd_sc_hd__o21ba_1 _4144_ (.A1(_1746_),
    .A2(_1747_),
    .B1_N(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__o31a_1 _4145_ (.A1(_1693_),
    .A2(_1744_),
    .A3(_1745_),
    .B1(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__nand2_1 _4146_ (.A(net188),
    .B(_1566_),
    .Y(_1751_));
 sky130_fd_sc_hd__a31o_1 _4147_ (.A1(_1493_),
    .A2(_1559_),
    .A3(_1565_),
    .B1(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__a211o_1 _4148_ (.A1(_1533_),
    .A2(_1534_),
    .B1(_1535_),
    .C1(_1542_),
    .X(_1753_));
 sky130_fd_sc_hd__nand2_1 _4149_ (.A(_1548_),
    .B(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__o211a_1 _4150_ (.A1(_1543_),
    .A2(_1754_),
    .B1(_1752_),
    .C1(_1750_),
    .X(_1755_));
 sky130_fd_sc_hd__o211a_1 _4151_ (.A1(_1583_),
    .A2(_1584_),
    .B1(_1586_),
    .C1(_1595_),
    .X(_1756_));
 sky130_fd_sc_hd__o21a_1 _4152_ (.A1(_1596_),
    .A2(_1756_),
    .B1(_1603_),
    .X(_1757_));
 sky130_fd_sc_hd__o211ai_4 _4153_ (.A1(net185),
    .A2(_0497_),
    .B1(_1743_),
    .C1(net171),
    .Y(_1758_));
 sky130_fd_sc_hd__o21ai_1 _4154_ (.A1(_1755_),
    .A2(_1757_),
    .B1(net175),
    .Y(_1759_));
 sky130_fd_sc_hd__a32o_1 _4155_ (.A1(_1670_),
    .A2(_1758_),
    .A3(_1759_),
    .B1(net194),
    .B2(net7),
    .X(_1760_));
 sky130_fd_sc_hd__mux2_1 _4156_ (.A0(net214),
    .A1(_1760_),
    .S(_1662_),
    .X(_0315_));
 sky130_fd_sc_hd__nor2_1 _4157_ (.A(net191),
    .B(_0997_),
    .Y(_1761_));
 sky130_fd_sc_hd__nand2_1 _4158_ (.A(net188),
    .B(_1617_),
    .Y(_1762_));
 sky130_fd_sc_hd__a31o_1 _4159_ (.A1(_1488_),
    .A2(_1557_),
    .A3(_1616_),
    .B1(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__a21oi_1 _4160_ (.A1(_1493_),
    .A2(_1737_),
    .B1(_1492_),
    .Y(_1764_));
 sky130_fd_sc_hd__nor2_1 _4161_ (.A(_1489_),
    .B(_1764_),
    .Y(_1765_));
 sky130_fd_sc_hd__a21o_1 _4162_ (.A1(_1489_),
    .A2(_1764_),
    .B1(_1980_),
    .X(_1766_));
 sky130_fd_sc_hd__a22o_1 _4163_ (.A1(net212),
    .A2(net157),
    .B1(net178),
    .B2(net214),
    .X(_1767_));
 sky130_fd_sc_hd__a2bb2o_1 _4164_ (.A1_N(_1257_),
    .A2_N(_1556_),
    .B1(_1489_),
    .B2(_1987_),
    .X(_1768_));
 sky130_fd_sc_hd__a2111o_1 _4165_ (.A1(_1507_),
    .A2(_1582_),
    .B1(_1508_),
    .C1(net202),
    .D1(_1976_),
    .X(_1769_));
 sky130_fd_sc_hd__o211ai_1 _4166_ (.A1(_1765_),
    .A2(_1766_),
    .B1(_1769_),
    .C1(_1763_),
    .Y(_1770_));
 sky130_fd_sc_hd__or4_1 _4167_ (.A(_1664_),
    .B(_1767_),
    .C(_1768_),
    .D(_1770_),
    .X(_1771_));
 sky130_fd_sc_hd__o311a_1 _4168_ (.A1(net213),
    .A2(net34),
    .A3(_1665_),
    .B1(_1771_),
    .C1(net191),
    .X(_1772_));
 sky130_fd_sc_hd__o21ai_2 _4169_ (.A1(_1761_),
    .A2(_1772_),
    .B1(net186),
    .Y(_1773_));
 sky130_fd_sc_hd__o211ai_4 _4170_ (.A1(net185),
    .A2(net79),
    .B1(_1773_),
    .C1(net171),
    .Y(_1774_));
 sky130_fd_sc_hd__a211o_1 _4171_ (.A1(_1491_),
    .A2(_1581_),
    .B1(_1583_),
    .C1(_1596_),
    .X(_1775_));
 sky130_fd_sc_hd__and3_1 _4172_ (.A(_1597_),
    .B(_1603_),
    .C(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__a211o_1 _4173_ (.A1(_1530_),
    .A2(_1531_),
    .B1(_1532_),
    .C1(_1543_),
    .X(_1777_));
 sky130_fd_sc_hd__a311o_1 _4174_ (.A1(_1544_),
    .A2(_1548_),
    .A3(_1777_),
    .B1(_1767_),
    .C1(net172),
    .X(_1778_));
 sky130_fd_sc_hd__o21ai_2 _4175_ (.A1(_1490_),
    .A2(_1744_),
    .B1(_1488_),
    .Y(_1779_));
 sky130_fd_sc_hd__o211a_1 _4176_ (.A1(_1581_),
    .A2(_1744_),
    .B1(_1779_),
    .C1(_1692_),
    .X(_1780_));
 sky130_fd_sc_hd__nand3_1 _4177_ (.A(_1488_),
    .B(_1557_),
    .C(_1566_),
    .Y(_1781_));
 sky130_fd_sc_hd__a31o_1 _4178_ (.A1(net188),
    .A2(_1567_),
    .A3(_1781_),
    .B1(_1780_),
    .X(_1782_));
 sky130_fd_sc_hd__o21ai_2 _4179_ (.A1(_1492_),
    .A2(_1746_),
    .B1(_1488_),
    .Y(_1783_));
 sky130_fd_sc_hd__o211a_1 _4180_ (.A1(_1531_),
    .A2(_1746_),
    .B1(_1783_),
    .C1(_1697_),
    .X(_1784_));
 sky130_fd_sc_hd__or4_2 _4181_ (.A(_1776_),
    .B(_1778_),
    .C(_1782_),
    .D(_1784_),
    .X(_1785_));
 sky130_fd_sc_hd__a32o_1 _4182_ (.A1(_1670_),
    .A2(_1774_),
    .A3(_1785_),
    .B1(net194),
    .B2(net8),
    .X(_1786_));
 sky130_fd_sc_hd__mux2_1 _4183_ (.A0(net213),
    .A1(_1786_),
    .S(_1662_),
    .X(_0316_));
 sky130_fd_sc_hd__nor2_1 _4184_ (.A(net191),
    .B(_1045_),
    .Y(_1787_));
 sky130_fd_sc_hd__nand3_1 _4185_ (.A(net182),
    .B(_1556_),
    .C(_1617_),
    .Y(_1788_));
 sky130_fd_sc_hd__o21a_1 _4186_ (.A1(_1487_),
    .A2(_1765_),
    .B1(net182),
    .X(_1789_));
 sky130_fd_sc_hd__o21ba_1 _4187_ (.A1(_1528_),
    .A2(_1765_),
    .B1_N(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__or3_1 _4188_ (.A(net182),
    .B(_1486_),
    .C(_1508_),
    .X(_1791_));
 sky130_fd_sc_hd__a22o_1 _4189_ (.A1(\as1802.D[6] ),
    .A2(net157),
    .B1(net178),
    .B2(\as1802.D[4] ),
    .X(_1792_));
 sky130_fd_sc_hd__o22a_1 _4190_ (.A1(_1986_),
    .A2(net182),
    .B1(_1555_),
    .B2(_1257_),
    .X(_1793_));
 sky130_fd_sc_hd__or3b_1 _4191_ (.A(_1664_),
    .B(_1792_),
    .C_N(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__a31o_1 _4192_ (.A1(_1981_),
    .A2(_1509_),
    .A3(_1791_),
    .B1(_1794_),
    .X(_1795_));
 sky130_fd_sc_hd__a21o_1 _4193_ (.A1(_1979_),
    .A2(_1790_),
    .B1(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__a31o_1 _4194_ (.A1(_1954_),
    .A2(_1618_),
    .A3(_1788_),
    .B1(_1796_),
    .X(_1797_));
 sky130_fd_sc_hd__o311a_1 _4195_ (.A1(net212),
    .A2(net35),
    .A3(_1665_),
    .B1(_1797_),
    .C1(net191),
    .X(_1798_));
 sky130_fd_sc_hd__o21ai_1 _4196_ (.A1(_1787_),
    .A2(_1798_),
    .B1(net185),
    .Y(_1799_));
 sky130_fd_sc_hd__o211ai_1 _4197_ (.A1(net185),
    .A2(_0610_),
    .B1(_1799_),
    .C1(net170),
    .Y(_1800_));
 sky130_fd_sc_hd__o211ai_1 _4198_ (.A1(_1579_),
    .A2(_1580_),
    .B1(_1597_),
    .C1(_1491_),
    .Y(_1801_));
 sky130_fd_sc_hd__o21a_1 _4199_ (.A1(_1485_),
    .A2(_1779_),
    .B1(_1578_),
    .X(_1802_));
 sky130_fd_sc_hd__nand2_1 _4200_ (.A(_1580_),
    .B(_1779_),
    .Y(_1803_));
 sky130_fd_sc_hd__o21a_1 _4201_ (.A1(_1485_),
    .A2(_1783_),
    .B1(_1527_),
    .X(_1804_));
 sky130_fd_sc_hd__nand2b_1 _4202_ (.A_N(_1528_),
    .B(_1783_),
    .Y(_1805_));
 sky130_fd_sc_hd__a311o_1 _4203_ (.A1(_1697_),
    .A2(_1804_),
    .A3(_1805_),
    .B1(_1792_),
    .C1(net172),
    .X(_1806_));
 sky130_fd_sc_hd__nand3_1 _4204_ (.A(_1529_),
    .B(_1530_),
    .C(_1544_),
    .Y(_1807_));
 sky130_fd_sc_hd__nand3_1 _4205_ (.A(net182),
    .B(_1556_),
    .C(_1567_),
    .Y(_1808_));
 sky130_fd_sc_hd__a31o_1 _4206_ (.A1(_1954_),
    .A2(_1568_),
    .A3(_1808_),
    .B1(_1806_),
    .X(_1809_));
 sky130_fd_sc_hd__a31o_1 _4207_ (.A1(_1545_),
    .A2(_1548_),
    .A3(_1807_),
    .B1(_1809_),
    .X(_1810_));
 sky130_fd_sc_hd__a31o_1 _4208_ (.A1(_1692_),
    .A2(_1802_),
    .A3(_1803_),
    .B1(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__a31o_1 _4209_ (.A1(_1598_),
    .A2(_1603_),
    .A3(_1801_),
    .B1(_1811_),
    .X(_1812_));
 sky130_fd_sc_hd__a32o_1 _4210_ (.A1(_1670_),
    .A2(_1800_),
    .A3(_1812_),
    .B1(net194),
    .B2(net9),
    .X(_1813_));
 sky130_fd_sc_hd__mux2_1 _4211_ (.A0(net212),
    .A1(_1813_),
    .S(_1662_),
    .X(_0317_));
 sky130_fd_sc_hd__nand3_1 _4212_ (.A(_1518_),
    .B(_1555_),
    .C(_1618_),
    .Y(_1814_));
 sky130_fd_sc_hd__or3b_1 _4213_ (.A(_1789_),
    .B(_1518_),
    .C_N(_1483_),
    .X(_1815_));
 sky130_fd_sc_hd__a21oi_1 _4214_ (.A1(_1518_),
    .A2(_1789_),
    .B1(_1525_),
    .Y(_1816_));
 sky130_fd_sc_hd__and3_1 _4215_ (.A(_1979_),
    .B(_1815_),
    .C(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__or2_1 _4216_ (.A(_1510_),
    .B(_1519_),
    .X(_1818_));
 sky130_fd_sc_hd__nand2_1 _4217_ (.A(_1509_),
    .B(_1577_),
    .Y(_1819_));
 sky130_fd_sc_hd__a22o_1 _4218_ (.A1(net210),
    .A2(net157),
    .B1(net178),
    .B2(net212),
    .X(_1820_));
 sky130_fd_sc_hd__o22a_1 _4219_ (.A1(_1986_),
    .A2(_1518_),
    .B1(_1554_),
    .B2(_1257_),
    .X(_1821_));
 sky130_fd_sc_hd__a31o_1 _4220_ (.A1(net188),
    .A2(_1619_),
    .A3(_1814_),
    .B1(_1820_),
    .X(_1822_));
 sky130_fd_sc_hd__or4b_1 _4221_ (.A(_1664_),
    .B(_1822_),
    .C(_1817_),
    .D_N(_1821_),
    .X(_1823_));
 sky130_fd_sc_hd__a31o_1 _4222_ (.A1(_1981_),
    .A2(_1818_),
    .A3(_1819_),
    .B1(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__o311a_1 _4223_ (.A1(\as1802.D[6] ),
    .A2(net205),
    .A3(_1665_),
    .B1(_1824_),
    .C1(net191),
    .X(_1825_));
 sky130_fd_sc_hd__nor2_1 _4224_ (.A(net191),
    .B(_1102_),
    .Y(_1826_));
 sky130_fd_sc_hd__o21ai_1 _4225_ (.A1(_1825_),
    .A2(_1826_),
    .B1(net186),
    .Y(_1827_));
 sky130_fd_sc_hd__o211a_1 _4226_ (.A1(net186),
    .A2(_0667_),
    .B1(_1827_),
    .C1(net170),
    .X(_1828_));
 sky130_fd_sc_hd__o211ai_1 _4227_ (.A1(_1575_),
    .A2(_1577_),
    .B1(_1578_),
    .C1(_1598_),
    .Y(_1829_));
 sky130_fd_sc_hd__and3_1 _4228_ (.A(_1599_),
    .B(_1603_),
    .C(_1829_),
    .X(_1830_));
 sky130_fd_sc_hd__nand2_1 _4229_ (.A(net188),
    .B(_1569_),
    .Y(_1831_));
 sky130_fd_sc_hd__a31o_1 _4230_ (.A1(_1518_),
    .A2(_1555_),
    .A3(_1568_),
    .B1(_1831_),
    .X(_1832_));
 sky130_fd_sc_hd__o211a_1 _4231_ (.A1(_1525_),
    .A2(_1526_),
    .B1(_1527_),
    .C1(_1545_),
    .X(_1833_));
 sky130_fd_sc_hd__o41a_1 _4232_ (.A1(net230),
    .A2(_1980_),
    .A3(_1546_),
    .A4(_1833_),
    .B1(_1832_),
    .X(_1834_));
 sky130_fd_sc_hd__nand2_1 _4233_ (.A(_1577_),
    .B(_1802_),
    .Y(_1835_));
 sky130_fd_sc_hd__a21o_1 _4234_ (.A1(_1482_),
    .A2(_1802_),
    .B1(_1519_),
    .X(_1836_));
 sky130_fd_sc_hd__and3_1 _4235_ (.A(_1692_),
    .B(_1835_),
    .C(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__a21oi_2 _4236_ (.A1(_1483_),
    .A2(_1804_),
    .B1(_1519_),
    .Y(_1838_));
 sky130_fd_sc_hd__a211o_1 _4237_ (.A1(_1526_),
    .A2(_1804_),
    .B1(_1838_),
    .C1(_1698_),
    .X(_1839_));
 sky130_fd_sc_hd__or4b_1 _4238_ (.A(net173),
    .B(_1820_),
    .C(_1837_),
    .D_N(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__or3b_1 _4239_ (.A(_1840_),
    .B(_1830_),
    .C_N(_1834_),
    .X(_1841_));
 sky130_fd_sc_hd__nand2_1 _4240_ (.A(_1670_),
    .B(_1841_),
    .Y(_1842_));
 sky130_fd_sc_hd__nand2_1 _4241_ (.A(net10),
    .B(net194),
    .Y(_1843_));
 sky130_fd_sc_hd__o21ai_1 _4242_ (.A1(_1828_),
    .A2(_1842_),
    .B1(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__mux2_1 _4243_ (.A0(\as1802.D[6] ),
    .A1(_1844_),
    .S(_1662_),
    .X(_0318_));
 sky130_fd_sc_hd__xnor2_1 _4244_ (.A(_1511_),
    .B(_1517_),
    .Y(_1845_));
 sky130_fd_sc_hd__and3_1 _4245_ (.A(_1516_),
    .B(_1554_),
    .C(_1619_),
    .X(_1846_));
 sky130_fd_sc_hd__nor2_1 _4246_ (.A(_1620_),
    .B(_1846_),
    .Y(_1847_));
 sky130_fd_sc_hd__mux2_1 _4247_ (.A0(_1517_),
    .A1(_1524_),
    .S(_1816_),
    .X(_1848_));
 sky130_fd_sc_hd__nor2_1 _4248_ (.A(_1986_),
    .B(_1516_),
    .Y(_1849_));
 sky130_fd_sc_hd__a31o_1 _4249_ (.A1(net210),
    .A2(net204),
    .A3(_1256_),
    .B1(_1849_),
    .X(_1850_));
 sky130_fd_sc_hd__a211o_1 _4250_ (.A1(\as1802.D[6] ),
    .A2(net178),
    .B1(_1664_),
    .C1(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__a31o_1 _4251_ (.A1(_1979_),
    .A2(_1523_),
    .A3(_1848_),
    .B1(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__a221o_1 _4252_ (.A1(_1981_),
    .A2(_1845_),
    .B1(_1847_),
    .B2(_1954_),
    .C1(_1852_),
    .X(_1853_));
 sky130_fd_sc_hd__o31a_1 _4253_ (.A1(net210),
    .A2(net204),
    .A3(_1665_),
    .B1(_2036_),
    .X(_1854_));
 sky130_fd_sc_hd__a22o_1 _4254_ (.A1(_2035_),
    .A2(_1150_),
    .B1(_1853_),
    .B2(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__o21ai_1 _4255_ (.A1(net186),
    .A2(_0716_),
    .B1(net170),
    .Y(_1856_));
 sky130_fd_sc_hd__a21o_1 _4256_ (.A1(net186),
    .A2(_1855_),
    .B1(_1856_),
    .X(_1857_));
 sky130_fd_sc_hd__a31o_1 _4257_ (.A1(_1574_),
    .A2(_1576_),
    .A3(_1599_),
    .B1(_1602_),
    .X(_1858_));
 sky130_fd_sc_hd__and2b_1 _4258_ (.A_N(_1858_),
    .B(_1600_),
    .X(_1859_));
 sky130_fd_sc_hd__a211o_1 _4259_ (.A1(_1523_),
    .A2(_1524_),
    .B1(_1525_),
    .C1(_1546_),
    .X(_1860_));
 sky130_fd_sc_hd__and3b_1 _4260_ (.A_N(_1547_),
    .B(_1548_),
    .C(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__and3_1 _4261_ (.A(_1516_),
    .B(_1554_),
    .C(_1569_),
    .X(_1862_));
 sky130_fd_sc_hd__or3_1 _4262_ (.A(_1955_),
    .B(_1570_),
    .C(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__mux2_1 _4263_ (.A0(_1524_),
    .A1(_1517_),
    .S(_1838_),
    .X(_1864_));
 sky130_fd_sc_hd__and3_1 _4264_ (.A(_1523_),
    .B(_1697_),
    .C(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(_1516_),
    .A1(_1573_),
    .S(_1836_),
    .X(_1866_));
 sky130_fd_sc_hd__or3_1 _4266_ (.A(_1572_),
    .B(_1693_),
    .C(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__a221o_1 _4267_ (.A1(\as1802.DF ),
    .A2(net157),
    .B1(net178),
    .B2(\as1802.D[6] ),
    .C1(net173),
    .X(_1868_));
 sky130_fd_sc_hd__or3b_1 _4268_ (.A(_1865_),
    .B(_1868_),
    .C_N(_1867_),
    .X(_1869_));
 sky130_fd_sc_hd__or4b_2 _4269_ (.A(_1859_),
    .B(_1861_),
    .C(_1869_),
    .D_N(_1863_),
    .X(_1870_));
 sky130_fd_sc_hd__and2_1 _4270_ (.A(net11),
    .B(net194),
    .X(_1871_));
 sky130_fd_sc_hd__a31o_1 _4271_ (.A1(_1670_),
    .A2(_1857_),
    .A3(_1870_),
    .B1(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__mux2_1 _4272_ (.A0(net210),
    .A1(_1872_),
    .S(_1662_),
    .X(_0319_));
 sky130_fd_sc_hd__o221a_1 _4273_ (.A1(_2023_),
    .A2(_2044_),
    .B1(_1650_),
    .B2(_1922_),
    .C1(_1448_),
    .X(_1873_));
 sky130_fd_sc_hd__o2111a_1 _4274_ (.A1(_1966_),
    .A2(_1210_),
    .B1(_1653_),
    .C1(_1655_),
    .D1(_1873_),
    .X(_1874_));
 sky130_fd_sc_hd__o41a_2 _4275_ (.A1(net272),
    .A2(_2017_),
    .A3(_2022_),
    .A4(_1255_),
    .B1(_1874_),
    .X(_1875_));
 sky130_fd_sc_hd__o31ai_4 _4276_ (.A1(net193),
    .A2(_1943_),
    .A3(_1460_),
    .B1(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__a22o_1 _4277_ (.A1(\as1802.P[0] ),
    .A2(_2092_),
    .B1(_1298_),
    .B2(\as1802.T[0] ),
    .X(_1877_));
 sky130_fd_sc_hd__nand2b_4 _4278_ (.A_N(_2091_),
    .B(_1207_),
    .Y(_1878_));
 sky130_fd_sc_hd__a22o_1 _4279_ (.A1(net158),
    .A2(_1877_),
    .B1(_1878_),
    .B2(net218),
    .X(_1879_));
 sky130_fd_sc_hd__mux2_1 _4280_ (.A0(net1),
    .A1(_1879_),
    .S(net196),
    .X(_1880_));
 sky130_fd_sc_hd__mux2_1 _4281_ (.A0(_1880_),
    .A1(net209),
    .S(_1876_),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _4282_ (.A1(\as1802.P[1] ),
    .A2(_2092_),
    .B1(_1298_),
    .B2(\as1802.T[1] ),
    .X(_1881_));
 sky130_fd_sc_hd__a22o_1 _4283_ (.A1(net217),
    .A2(_1878_),
    .B1(_1881_),
    .B2(net158),
    .X(_1882_));
 sky130_fd_sc_hd__mux2_1 _4284_ (.A0(net5),
    .A1(_1882_),
    .S(net196),
    .X(_1883_));
 sky130_fd_sc_hd__mux2_1 _4285_ (.A0(_1883_),
    .A1(net207),
    .S(_1876_),
    .X(_0325_));
 sky130_fd_sc_hd__a22o_1 _4286_ (.A1(\as1802.P[2] ),
    .A2(_2092_),
    .B1(_1298_),
    .B2(\as1802.T[2] ),
    .X(_1884_));
 sky130_fd_sc_hd__a22o_1 _4287_ (.A1(net215),
    .A2(_1878_),
    .B1(_1884_),
    .B2(net158),
    .X(_1885_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(net6),
    .A1(_1885_),
    .S(net196),
    .X(_1886_));
 sky130_fd_sc_hd__mux2_1 _4289_ (.A0(_1886_),
    .A1(net206),
    .S(_1876_),
    .X(_0326_));
 sky130_fd_sc_hd__a22o_1 _4290_ (.A1(\as1802.P[3] ),
    .A2(_2092_),
    .B1(_1298_),
    .B2(\as1802.T[3] ),
    .X(_1887_));
 sky130_fd_sc_hd__a22o_1 _4291_ (.A1(\as1802.D[3] ),
    .A2(_1878_),
    .B1(_1887_),
    .B2(net158),
    .X(_1888_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(net7),
    .A1(_1888_),
    .S(net196),
    .X(_1889_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(_1889_),
    .A1(net33),
    .S(_1876_),
    .X(_0327_));
 sky130_fd_sc_hd__a22o_1 _4294_ (.A1(\as1802.X[0] ),
    .A2(_2092_),
    .B1(_1298_),
    .B2(\as1802.T[4] ),
    .X(_1890_));
 sky130_fd_sc_hd__a22o_1 _4295_ (.A1(\as1802.D[4] ),
    .A2(_1878_),
    .B1(_1890_),
    .B2(net158),
    .X(_1891_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(net8),
    .A1(_1891_),
    .S(net196),
    .X(_1892_));
 sky130_fd_sc_hd__mux2_1 _4297_ (.A0(_1892_),
    .A1(net34),
    .S(_1876_),
    .X(_0328_));
 sky130_fd_sc_hd__a22o_1 _4298_ (.A1(\as1802.X[1] ),
    .A2(_2092_),
    .B1(_1298_),
    .B2(\as1802.T[5] ),
    .X(_1893_));
 sky130_fd_sc_hd__a22o_1 _4299_ (.A1(\as1802.D[5] ),
    .A2(_1878_),
    .B1(_1893_),
    .B2(net158),
    .X(_1894_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(net9),
    .A1(_1894_),
    .S(net196),
    .X(_1895_));
 sky130_fd_sc_hd__mux2_1 _4301_ (.A0(_1895_),
    .A1(net35),
    .S(_1876_),
    .X(_0329_));
 sky130_fd_sc_hd__a22o_1 _4302_ (.A1(\as1802.X[2] ),
    .A2(_2092_),
    .B1(_1298_),
    .B2(\as1802.T[6] ),
    .X(_1896_));
 sky130_fd_sc_hd__a22o_1 _4303_ (.A1(\as1802.D[6] ),
    .A2(_1878_),
    .B1(_1896_),
    .B2(net158),
    .X(_1897_));
 sky130_fd_sc_hd__a21bo_1 _4304_ (.A1(net195),
    .A2(_1897_),
    .B1_N(_1843_),
    .X(_1898_));
 sky130_fd_sc_hd__mux2_1 _4305_ (.A0(_1898_),
    .A1(net205),
    .S(_1876_),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _4306_ (.A1(\as1802.X[3] ),
    .A2(_2092_),
    .B1(_1298_),
    .B2(\as1802.T[7] ),
    .X(_1899_));
 sky130_fd_sc_hd__a22o_1 _4307_ (.A1(net210),
    .A2(_1878_),
    .B1(_1899_),
    .B2(_1207_),
    .X(_1900_));
 sky130_fd_sc_hd__a21o_1 _4308_ (.A1(net195),
    .A2(_1900_),
    .B1(_1871_),
    .X(_1901_));
 sky130_fd_sc_hd__mux2_2 _4309_ (.A0(_1901_),
    .A1(net37),
    .S(_1876_),
    .X(_0331_));
 sky130_fd_sc_hd__and3_4 _4310_ (.A(_0759_),
    .B(net70),
    .C(_1196_),
    .X(_1902_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(\as1802.regs[9][8] ),
    .A1(net52),
    .S(_1902_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _4312_ (.A0(\as1802.regs[9][9] ),
    .A1(net50),
    .S(_1902_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(\as1802.regs[9][10] ),
    .A1(net48),
    .S(_1902_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _4314_ (.A0(\as1802.regs[9][11] ),
    .A1(net46),
    .S(_1902_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _4315_ (.A0(\as1802.regs[9][12] ),
    .A1(net45),
    .S(_1902_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _4316_ (.A0(\as1802.regs[9][13] ),
    .A1(net42),
    .S(_1902_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _4317_ (.A0(\as1802.regs[9][14] ),
    .A1(net40),
    .S(_1902_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _4318_ (.A0(\as1802.regs[9][15] ),
    .A1(net38),
    .S(_1902_),
    .X(_0339_));
 sky130_fd_sc_hd__and3_4 _4319_ (.A(_0758_),
    .B(net71),
    .C(_1191_),
    .X(_1903_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(\as1802.regs[2][8] ),
    .A1(net52),
    .S(_1903_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(\as1802.regs[2][9] ),
    .A1(net51),
    .S(_1903_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _4322_ (.A0(\as1802.regs[2][10] ),
    .A1(net49),
    .S(_1903_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _4323_ (.A0(\as1802.regs[2][11] ),
    .A1(net47),
    .S(_1903_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _4324_ (.A0(\as1802.regs[2][12] ),
    .A1(net45),
    .S(_1903_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(\as1802.regs[2][13] ),
    .A1(net43),
    .S(_1903_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(\as1802.regs[2][14] ),
    .A1(net41),
    .S(_1903_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _4327_ (.A0(\as1802.regs[2][15] ),
    .A1(net38),
    .S(_1903_),
    .X(_0347_));
 sky130_fd_sc_hd__a2bb2o_1 _4328_ (.A1_N(net270),
    .A2_N(net158),
    .B1(_1255_),
    .B2(_2053_),
    .X(_1904_));
 sky130_fd_sc_hd__mux2_1 _4329_ (.A0(_1904_),
    .A1(\as1802.mem_write ),
    .S(net76),
    .X(_0348_));
 sky130_fd_sc_hd__and3_4 _4330_ (.A(net71),
    .B(_1191_),
    .C(_1196_),
    .X(_1905_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(\as1802.regs[1][8] ),
    .A1(net53),
    .S(_1905_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _4332_ (.A0(\as1802.regs[1][9] ),
    .A1(net51),
    .S(_1905_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _4333_ (.A0(\as1802.regs[1][10] ),
    .A1(net49),
    .S(_1905_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _4334_ (.A0(\as1802.regs[1][11] ),
    .A1(net47),
    .S(_1905_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _4335_ (.A0(\as1802.regs[1][12] ),
    .A1(net45),
    .S(_1905_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(\as1802.regs[1][13] ),
    .A1(net43),
    .S(_1905_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _4337_ (.A0(\as1802.regs[1][14] ),
    .A1(net41),
    .S(_1905_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(\as1802.regs[1][15] ),
    .A1(net38),
    .S(_1905_),
    .X(_0356_));
 sky130_fd_sc_hd__o211a_1 _4339_ (.A1(\as1802.IE ),
    .A2(_1203_),
    .B1(net196),
    .C1(net273),
    .X(_1906_));
 sky130_fd_sc_hd__o211a_1 _4340_ (.A1(_1652_),
    .A2(_1906_),
    .B1(_1650_),
    .C1(_1651_),
    .X(_1907_));
 sky130_fd_sc_hd__nand2_1 _4341_ (.A(_1273_),
    .B(_1907_),
    .Y(_1908_));
 sky130_fd_sc_hd__mux2_1 _4342_ (.A0(_2038_),
    .A1(net30),
    .S(_1908_),
    .X(_0357_));
 sky130_fd_sc_hd__a22o_1 _4343_ (.A1(_1274_),
    .A2(_1907_),
    .B1(_1908_),
    .B2(net31),
    .X(_0358_));
 sky130_fd_sc_hd__o211a_1 _4344_ (.A1(\as1802.P[0] ),
    .A2(_1223_),
    .B1(_1225_),
    .C1(net276),
    .X(_0320_));
 sky130_fd_sc_hd__o21a_1 _4345_ (.A1(\as1802.P[1] ),
    .A2(_1223_),
    .B1(_1228_),
    .X(_0321_));
 sky130_fd_sc_hd__and2_1 _4346_ (.A(net277),
    .B(_1231_),
    .X(_0322_));
 sky130_fd_sc_hd__and2_1 _4347_ (.A(net277),
    .B(_1234_),
    .X(_0323_));
 sky130_fd_sc_hd__dfxtp_1 _4348_ (.CLK(clknet_leaf_1_clk),
    .D(_0012_),
    .Q(\as1802.regs[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4349_ (.CLK(clknet_leaf_3_clk),
    .D(_0013_),
    .Q(\as1802.regs[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4350_ (.CLK(clknet_leaf_6_clk),
    .D(_0014_),
    .Q(\as1802.regs[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4351_ (.CLK(clknet_leaf_7_clk),
    .D(_0015_),
    .Q(\as1802.regs[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4352_ (.CLK(clknet_leaf_0_clk),
    .D(_0016_),
    .Q(\as1802.regs[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4353_ (.CLK(clknet_leaf_52_clk),
    .D(_0017_),
    .Q(\as1802.regs[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4354_ (.CLK(clknet_leaf_51_clk),
    .D(_0018_),
    .Q(\as1802.regs[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4355_ (.CLK(clknet_leaf_52_clk),
    .D(_0019_),
    .Q(\as1802.regs[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4356_ (.CLK(clknet_leaf_46_clk),
    .D(_0020_),
    .Q(\as1802.regs[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4357_ (.CLK(clknet_leaf_49_clk),
    .D(_0021_),
    .Q(\as1802.regs[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4358_ (.CLK(clknet_leaf_41_clk),
    .D(_0022_),
    .Q(\as1802.regs[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4359_ (.CLK(clknet_leaf_37_clk),
    .D(_0023_),
    .Q(\as1802.regs[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4360_ (.CLK(clknet_leaf_41_clk),
    .D(_0024_),
    .Q(\as1802.regs[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4361_ (.CLK(clknet_leaf_43_clk),
    .D(_0025_),
    .Q(\as1802.regs[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4362_ (.CLK(clknet_leaf_39_clk),
    .D(_0026_),
    .Q(\as1802.regs[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4363_ (.CLK(clknet_leaf_35_clk),
    .D(_0027_),
    .Q(\as1802.regs[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4364_ (.CLK(clknet_leaf_44_clk),
    .D(_0028_),
    .Q(\as1802.regs[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4365_ (.CLK(clknet_leaf_45_clk),
    .D(_0029_),
    .Q(\as1802.regs[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4366_ (.CLK(clknet_leaf_47_clk),
    .D(_0030_),
    .Q(\as1802.regs[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4367_ (.CLK(clknet_leaf_34_clk),
    .D(_0031_),
    .Q(\as1802.regs[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4368_ (.CLK(clknet_leaf_44_clk),
    .D(_0032_),
    .Q(\as1802.regs[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4369_ (.CLK(clknet_leaf_35_clk),
    .D(_0033_),
    .Q(\as1802.regs[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4370_ (.CLK(clknet_leaf_33_clk),
    .D(_0034_),
    .Q(\as1802.regs[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4371_ (.CLK(clknet_leaf_33_clk),
    .D(_0035_),
    .Q(\as1802.regs[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4372_ (.CLK(clknet_leaf_46_clk),
    .D(_0036_),
    .Q(\as1802.regs[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4373_ (.CLK(clknet_leaf_48_clk),
    .D(_0037_),
    .Q(\as1802.regs[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4374_ (.CLK(clknet_leaf_48_clk),
    .D(_0038_),
    .Q(\as1802.regs[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4375_ (.CLK(clknet_leaf_37_clk),
    .D(_0039_),
    .Q(\as1802.regs[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4376_ (.CLK(clknet_leaf_40_clk),
    .D(_0040_),
    .Q(\as1802.regs[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4377_ (.CLK(clknet_leaf_43_clk),
    .D(_0041_),
    .Q(\as1802.regs[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4378_ (.CLK(clknet_leaf_38_clk),
    .D(_0042_),
    .Q(\as1802.regs[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4379_ (.CLK(clknet_leaf_39_clk),
    .D(_0043_),
    .Q(\as1802.regs[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4380_ (.CLK(clknet_leaf_42_clk),
    .D(_0044_),
    .Q(\as1802.regs[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4381_ (.CLK(clknet_leaf_48_clk),
    .D(_0045_),
    .Q(\as1802.regs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4382_ (.CLK(clknet_leaf_41_clk),
    .D(_0046_),
    .Q(\as1802.regs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4383_ (.CLK(clknet_leaf_37_clk),
    .D(_0047_),
    .Q(\as1802.regs[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4384_ (.CLK(clknet_leaf_39_clk),
    .D(_0048_),
    .Q(\as1802.regs[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4385_ (.CLK(clknet_leaf_35_clk),
    .D(_0049_),
    .Q(\as1802.regs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4386_ (.CLK(clknet_leaf_36_clk),
    .D(_0050_),
    .Q(\as1802.regs[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4387_ (.CLK(clknet_leaf_36_clk),
    .D(_0051_),
    .Q(\as1802.regs[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4388_ (.CLK(clknet_leaf_42_clk),
    .D(_0052_),
    .Q(\as1802.regs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4389_ (.CLK(clknet_leaf_48_clk),
    .D(_0053_),
    .Q(\as1802.regs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4390_ (.CLK(clknet_leaf_41_clk),
    .D(_0054_),
    .Q(\as1802.regs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4391_ (.CLK(clknet_leaf_37_clk),
    .D(_0055_),
    .Q(\as1802.regs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4392_ (.CLK(clknet_leaf_39_clk),
    .D(_0056_),
    .Q(\as1802.regs[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4393_ (.CLK(clknet_leaf_35_clk),
    .D(_0057_),
    .Q(\as1802.regs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4394_ (.CLK(clknet_leaf_36_clk),
    .D(_0058_),
    .Q(\as1802.regs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4395_ (.CLK(clknet_leaf_36_clk),
    .D(_0059_),
    .Q(\as1802.regs[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4396_ (.CLK(clknet_leaf_42_clk),
    .D(_0060_),
    .Q(\as1802.regs[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4397_ (.CLK(clknet_leaf_47_clk),
    .D(_0061_),
    .Q(\as1802.regs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4398_ (.CLK(clknet_leaf_48_clk),
    .D(_0062_),
    .Q(\as1802.regs[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4399_ (.CLK(clknet_leaf_37_clk),
    .D(_0063_),
    .Q(\as1802.regs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4400_ (.CLK(clknet_leaf_41_clk),
    .D(_0064_),
    .Q(\as1802.regs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4401_ (.CLK(clknet_leaf_43_clk),
    .D(_0065_),
    .Q(\as1802.regs[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4402_ (.CLK(clknet_leaf_36_clk),
    .D(_0066_),
    .Q(\as1802.regs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4403_ (.CLK(clknet_leaf_36_clk),
    .D(_0067_),
    .Q(\as1802.regs[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4404_ (.CLK(clknet_leaf_44_clk),
    .D(_0068_),
    .Q(\as1802.regs[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4405_ (.CLK(clknet_leaf_48_clk),
    .D(_0069_),
    .Q(\as1802.regs[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4406_ (.CLK(clknet_leaf_47_clk),
    .D(_0070_),
    .Q(\as1802.regs[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4407_ (.CLK(clknet_leaf_37_clk),
    .D(_0071_),
    .Q(\as1802.regs[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4408_ (.CLK(clknet_leaf_42_clk),
    .D(_0072_),
    .Q(\as1802.regs[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4409_ (.CLK(clknet_leaf_43_clk),
    .D(_0073_),
    .Q(\as1802.regs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4410_ (.CLK(clknet_leaf_36_clk),
    .D(_0074_),
    .Q(\as1802.regs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4411_ (.CLK(clknet_leaf_35_clk),
    .D(_0075_),
    .Q(\as1802.regs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4412_ (.CLK(clknet_leaf_45_clk),
    .D(_0076_),
    .Q(\as1802.regs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4413_ (.CLK(clknet_leaf_45_clk),
    .D(_0077_),
    .Q(\as1802.regs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4414_ (.CLK(clknet_leaf_47_clk),
    .D(_0078_),
    .Q(\as1802.regs[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4415_ (.CLK(clknet_leaf_35_clk),
    .D(_0079_),
    .Q(\as1802.regs[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4416_ (.CLK(clknet_leaf_44_clk),
    .D(_0080_),
    .Q(\as1802.regs[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4417_ (.CLK(clknet_leaf_31_clk),
    .D(_0081_),
    .Q(\as1802.regs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4418_ (.CLK(clknet_leaf_34_clk),
    .D(_0082_),
    .Q(\as1802.regs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4419_ (.CLK(clknet_leaf_33_clk),
    .D(_0083_),
    .Q(\as1802.regs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4420_ (.CLK(clknet_leaf_2_clk),
    .D(_0084_),
    .Q(\as1802.regs[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4421_ (.CLK(clknet_leaf_3_clk),
    .D(_0085_),
    .Q(\as1802.regs[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4422_ (.CLK(clknet_leaf_6_clk),
    .D(_0086_),
    .Q(\as1802.regs[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4423_ (.CLK(clknet_leaf_7_clk),
    .D(_0087_),
    .Q(\as1802.regs[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4424_ (.CLK(clknet_leaf_3_clk),
    .D(_0088_),
    .Q(\as1802.regs[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4425_ (.CLK(clknet_leaf_0_clk),
    .D(_0089_),
    .Q(\as1802.regs[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4426_ (.CLK(clknet_leaf_50_clk),
    .D(_0090_),
    .Q(\as1802.regs[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4427_ (.CLK(clknet_leaf_2_clk),
    .D(_0091_),
    .Q(\as1802.regs[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4428_ (.CLK(clknet_leaf_1_clk),
    .D(_0092_),
    .Q(\as1802.regs[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4429_ (.CLK(clknet_leaf_3_clk),
    .D(_0093_),
    .Q(\as1802.regs[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4430_ (.CLK(clknet_leaf_6_clk),
    .D(_0094_),
    .Q(\as1802.regs[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4431_ (.CLK(clknet_leaf_7_clk),
    .D(_0095_),
    .Q(\as1802.regs[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4432_ (.CLK(clknet_leaf_3_clk),
    .D(_0096_),
    .Q(\as1802.regs[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4433_ (.CLK(clknet_leaf_0_clk),
    .D(_0097_),
    .Q(\as1802.regs[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4434_ (.CLK(clknet_leaf_46_clk),
    .D(_0098_),
    .Q(\as1802.regs[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4435_ (.CLK(clknet_leaf_2_clk),
    .D(_0099_),
    .Q(\as1802.regs[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4436_ (.CLK(clknet_leaf_25_clk),
    .D(_0004_),
    .Q(\as1802.instr_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_4 _4437_ (.CLK(clknet_leaf_27_clk),
    .D(_0005_),
    .Q(\as1802.instr_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4438_ (.CLK(clknet_leaf_28_clk),
    .D(_0006_),
    .Q(\as1802.instr_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4439_ (.CLK(clknet_leaf_26_clk),
    .D(_0007_),
    .Q(\as1802.instr_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_4 _4440_ (.CLK(clknet_leaf_11_clk),
    .D(_0100_),
    .Q(_0000_));
 sky130_fd_sc_hd__dfxtp_4 _4441_ (.CLK(clknet_leaf_10_clk),
    .D(_0101_),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_4 _4442_ (.CLK(clknet_leaf_11_clk),
    .D(_0102_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_1 _4443_ (.CLK(clknet_leaf_11_clk),
    .D(_0103_),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_1 _4444_ (.CLK(clknet_leaf_5_clk),
    .D(_0104_),
    .Q(\as1802.regs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4445_ (.CLK(clknet_leaf_14_clk),
    .D(_0105_),
    .Q(\as1802.regs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4446_ (.CLK(clknet_leaf_13_clk),
    .D(_0106_),
    .Q(\as1802.regs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4447_ (.CLK(clknet_leaf_16_clk),
    .D(_0107_),
    .Q(\as1802.regs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4448_ (.CLK(clknet_leaf_14_clk),
    .D(_0108_),
    .Q(\as1802.regs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4449_ (.CLK(clknet_leaf_4_clk),
    .D(_0109_),
    .Q(\as1802.regs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4450_ (.CLK(clknet_leaf_12_clk),
    .D(_0110_),
    .Q(\as1802.regs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4451_ (.CLK(clknet_leaf_4_clk),
    .D(_0111_),
    .Q(\as1802.regs[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4452_ (.CLK(clknet_leaf_4_clk),
    .D(_0112_),
    .Q(\as1802.regs[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4453_ (.CLK(clknet_leaf_15_clk),
    .D(_0113_),
    .Q(\as1802.regs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4454_ (.CLK(clknet_leaf_13_clk),
    .D(_0114_),
    .Q(\as1802.regs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4455_ (.CLK(clknet_leaf_16_clk),
    .D(_0115_),
    .Q(\as1802.regs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4456_ (.CLK(clknet_leaf_14_clk),
    .D(_0116_),
    .Q(\as1802.regs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4457_ (.CLK(clknet_leaf_4_clk),
    .D(_0117_),
    .Q(\as1802.regs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4458_ (.CLK(clknet_leaf_12_clk),
    .D(_0118_),
    .Q(\as1802.regs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4459_ (.CLK(clknet_leaf_4_clk),
    .D(_0119_),
    .Q(\as1802.regs[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4460_ (.CLK(clknet_leaf_5_clk),
    .D(_0120_),
    .Q(\as1802.regs[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4461_ (.CLK(clknet_leaf_15_clk),
    .D(_0121_),
    .Q(\as1802.regs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4462_ (.CLK(clknet_leaf_13_clk),
    .D(_0122_),
    .Q(\as1802.regs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4463_ (.CLK(clknet_leaf_16_clk),
    .D(_0123_),
    .Q(\as1802.regs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4464_ (.CLK(clknet_leaf_15_clk),
    .D(_0124_),
    .Q(\as1802.regs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4465_ (.CLK(clknet_leaf_13_clk),
    .D(_0125_),
    .Q(\as1802.regs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4466_ (.CLK(clknet_leaf_12_clk),
    .D(_0126_),
    .Q(\as1802.regs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4467_ (.CLK(clknet_leaf_4_clk),
    .D(_0127_),
    .Q(\as1802.regs[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4468_ (.CLK(clknet_leaf_12_clk),
    .D(_0128_),
    .Q(\as1802.regs[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4469_ (.CLK(clknet_leaf_16_clk),
    .D(_0129_),
    .Q(\as1802.regs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4470_ (.CLK(clknet_leaf_13_clk),
    .D(_0130_),
    .Q(\as1802.regs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4471_ (.CLK(clknet_leaf_16_clk),
    .D(_0131_),
    .Q(\as1802.regs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4472_ (.CLK(clknet_leaf_17_clk),
    .D(_0132_),
    .Q(\as1802.regs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4473_ (.CLK(clknet_leaf_13_clk),
    .D(_0133_),
    .Q(\as1802.regs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4474_ (.CLK(clknet_leaf_12_clk),
    .D(_0134_),
    .Q(\as1802.regs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4475_ (.CLK(clknet_leaf_4_clk),
    .D(_0135_),
    .Q(\as1802.regs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4476_ (.CLK(clknet_leaf_12_clk),
    .D(_0136_),
    .Q(\as1802.regs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4477_ (.CLK(clknet_leaf_11_clk),
    .D(_0137_),
    .Q(\as1802.regs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4478_ (.CLK(clknet_leaf_11_clk),
    .D(_0138_),
    .Q(\as1802.regs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4479_ (.CLK(clknet_leaf_11_clk),
    .D(_0139_),
    .Q(\as1802.regs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4480_ (.CLK(clknet_leaf_14_clk),
    .D(_0140_),
    .Q(\as1802.regs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4481_ (.CLK(clknet_leaf_13_clk),
    .D(_0141_),
    .Q(\as1802.regs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4482_ (.CLK(clknet_leaf_9_clk),
    .D(_0142_),
    .Q(\as1802.regs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4483_ (.CLK(clknet_leaf_4_clk),
    .D(_0143_),
    .Q(\as1802.regs[3][7] ));
 sky130_fd_sc_hd__dfxtp_4 _4484_ (.CLK(clknet_leaf_10_clk),
    .D(_0144_),
    .Q(\as1802.regs[2][0] ));
 sky130_fd_sc_hd__dfxtp_4 _4485_ (.CLK(clknet_leaf_9_clk),
    .D(_0145_),
    .Q(\as1802.regs[2][1] ));
 sky130_fd_sc_hd__dfxtp_4 _4486_ (.CLK(clknet_leaf_9_clk),
    .D(_0146_),
    .Q(\as1802.regs[2][2] ));
 sky130_fd_sc_hd__dfxtp_2 _4487_ (.CLK(clknet_leaf_10_clk),
    .D(_0147_),
    .Q(\as1802.regs[2][3] ));
 sky130_fd_sc_hd__dfxtp_4 _4488_ (.CLK(clknet_leaf_10_clk),
    .D(_0148_),
    .Q(\as1802.regs[2][4] ));
 sky130_fd_sc_hd__dfxtp_2 _4489_ (.CLK(clknet_leaf_9_clk),
    .D(_0149_),
    .Q(\as1802.regs[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4490_ (.CLK(clknet_leaf_9_clk),
    .D(_0150_),
    .Q(\as1802.regs[2][6] ));
 sky130_fd_sc_hd__dfxtp_2 _4491_ (.CLK(clknet_leaf_8_clk),
    .D(_0151_),
    .Q(\as1802.regs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4492_ (.CLK(clknet_leaf_12_clk),
    .D(_0152_),
    .Q(\as1802.regs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4493_ (.CLK(clknet_leaf_14_clk),
    .D(_0153_),
    .Q(\as1802.regs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4494_ (.CLK(clknet_leaf_11_clk),
    .D(_0154_),
    .Q(\as1802.regs[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4495_ (.CLK(clknet_leaf_11_clk),
    .D(_0155_),
    .Q(\as1802.regs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4496_ (.CLK(clknet_leaf_14_clk),
    .D(_0156_),
    .Q(\as1802.regs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4497_ (.CLK(clknet_leaf_12_clk),
    .D(_0157_),
    .Q(\as1802.regs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4498_ (.CLK(clknet_leaf_8_clk),
    .D(_0158_),
    .Q(\as1802.regs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4499_ (.CLK(clknet_leaf_4_clk),
    .D(_0159_),
    .Q(\as1802.regs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4500_ (.CLK(clknet_leaf_46_clk),
    .D(_0160_),
    .Q(\as1802.regs[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4501_ (.CLK(clknet_leaf_49_clk),
    .D(_0161_),
    .Q(\as1802.regs[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4502_ (.CLK(clknet_leaf_47_clk),
    .D(_0162_),
    .Q(\as1802.regs[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4503_ (.CLK(clknet_leaf_40_clk),
    .D(_0163_),
    .Q(\as1802.regs[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4504_ (.CLK(clknet_leaf_41_clk),
    .D(_0164_),
    .Q(\as1802.regs[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4505_ (.CLK(clknet_leaf_42_clk),
    .D(_0165_),
    .Q(\as1802.regs[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4506_ (.CLK(clknet_leaf_40_clk),
    .D(_0166_),
    .Q(\as1802.regs[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4507_ (.CLK(clknet_leaf_39_clk),
    .D(_0167_),
    .Q(\as1802.regs[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4508_ (.CLK(clknet_leaf_1_clk),
    .D(_0168_),
    .Q(\as1802.regs[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4509_ (.CLK(clknet_leaf_3_clk),
    .D(_0169_),
    .Q(\as1802.regs[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4510_ (.CLK(clknet_leaf_6_clk),
    .D(_0170_),
    .Q(\as1802.regs[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4511_ (.CLK(clknet_leaf_7_clk),
    .D(_0171_),
    .Q(\as1802.regs[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4512_ (.CLK(clknet_leaf_0_clk),
    .D(_0172_),
    .Q(\as1802.regs[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4513_ (.CLK(clknet_leaf_52_clk),
    .D(_0173_),
    .Q(\as1802.regs[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4514_ (.CLK(clknet_leaf_51_clk),
    .D(_0174_),
    .Q(\as1802.regs[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4515_ (.CLK(clknet_leaf_51_clk),
    .D(_0175_),
    .Q(\as1802.regs[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4516_ (.CLK(clknet_leaf_50_clk),
    .D(_0176_),
    .Q(\as1802.regs[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4517_ (.CLK(clknet_leaf_2_clk),
    .D(_0177_),
    .Q(\as1802.regs[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4518_ (.CLK(clknet_leaf_6_clk),
    .D(_0178_),
    .Q(\as1802.regs[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4519_ (.CLK(clknet_leaf_7_clk),
    .D(_0179_),
    .Q(\as1802.regs[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4520_ (.CLK(clknet_leaf_0_clk),
    .D(_0180_),
    .Q(\as1802.regs[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4521_ (.CLK(clknet_leaf_52_clk),
    .D(_0181_),
    .Q(\as1802.regs[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4522_ (.CLK(clknet_leaf_49_clk),
    .D(_0182_),
    .Q(\as1802.regs[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4523_ (.CLK(clknet_leaf_51_clk),
    .D(_0183_),
    .Q(\as1802.regs[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4524_ (.CLK(clknet_leaf_47_clk),
    .D(_0184_),
    .Q(\as1802.regs[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4525_ (.CLK(clknet_leaf_49_clk),
    .D(_0185_),
    .Q(\as1802.regs[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4526_ (.CLK(clknet_leaf_41_clk),
    .D(_0186_),
    .Q(\as1802.regs[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4527_ (.CLK(clknet_leaf_38_clk),
    .D(_0187_),
    .Q(\as1802.regs[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4528_ (.CLK(clknet_leaf_40_clk),
    .D(_0188_),
    .Q(\as1802.regs[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4529_ (.CLK(clknet_leaf_39_clk),
    .D(_0189_),
    .Q(\as1802.regs[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4530_ (.CLK(clknet_leaf_40_clk),
    .D(_0190_),
    .Q(\as1802.regs[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4531_ (.CLK(clknet_leaf_39_clk),
    .D(_0191_),
    .Q(\as1802.regs[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4532_ (.CLK(clknet_leaf_1_clk),
    .D(_0192_),
    .Q(\as1802.regs[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4533_ (.CLK(clknet_leaf_3_clk),
    .D(_0193_),
    .Q(\as1802.regs[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4534_ (.CLK(clknet_leaf_6_clk),
    .D(_0194_),
    .Q(\as1802.regs[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4535_ (.CLK(clknet_leaf_7_clk),
    .D(_0195_),
    .Q(\as1802.regs[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4536_ (.CLK(clknet_leaf_3_clk),
    .D(_0196_),
    .Q(\as1802.regs[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4537_ (.CLK(clknet_leaf_0_clk),
    .D(_0197_),
    .Q(\as1802.regs[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4538_ (.CLK(clknet_leaf_49_clk),
    .D(_0198_),
    .Q(\as1802.regs[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4539_ (.CLK(clknet_leaf_1_clk),
    .D(_0199_),
    .Q(\as1802.regs[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4540_ (.CLK(clknet_leaf_1_clk),
    .D(_0200_),
    .Q(\as1802.regs[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4541_ (.CLK(clknet_leaf_3_clk),
    .D(_0201_),
    .Q(\as1802.regs[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4542_ (.CLK(clknet_leaf_6_clk),
    .D(_0202_),
    .Q(\as1802.regs[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4543_ (.CLK(clknet_leaf_7_clk),
    .D(_0203_),
    .Q(\as1802.regs[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4544_ (.CLK(clknet_leaf_3_clk),
    .D(_0204_),
    .Q(\as1802.regs[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4545_ (.CLK(clknet_leaf_52_clk),
    .D(_0205_),
    .Q(\as1802.regs[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4546_ (.CLK(clknet_leaf_50_clk),
    .D(_0206_),
    .Q(\as1802.regs[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4547_ (.CLK(clknet_leaf_2_clk),
    .D(_0207_),
    .Q(\as1802.regs[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4548_ (.CLK(clknet_leaf_5_clk),
    .D(_0208_),
    .Q(\as1802.regs[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4549_ (.CLK(clknet_leaf_11_clk),
    .D(_0209_),
    .Q(\as1802.regs[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4550_ (.CLK(clknet_leaf_10_clk),
    .D(_0210_),
    .Q(\as1802.regs[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4551_ (.CLK(clknet_leaf_10_clk),
    .D(_0211_),
    .Q(\as1802.regs[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4552_ (.CLK(clknet_leaf_14_clk),
    .D(_0212_),
    .Q(\as1802.regs[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4553_ (.CLK(clknet_leaf_12_clk),
    .D(_0213_),
    .Q(\as1802.regs[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4554_ (.CLK(clknet_leaf_8_clk),
    .D(_0214_),
    .Q(\as1802.regs[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4555_ (.CLK(clknet_leaf_4_clk),
    .D(_0215_),
    .Q(\as1802.regs[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4556_ (.CLK(clknet_leaf_46_clk),
    .D(_0216_),
    .Q(\as1802.regs[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4557_ (.CLK(clknet_leaf_49_clk),
    .D(_0217_),
    .Q(\as1802.regs[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4558_ (.CLK(clknet_leaf_47_clk),
    .D(_0218_),
    .Q(\as1802.regs[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4559_ (.CLK(clknet_leaf_40_clk),
    .D(_0219_),
    .Q(\as1802.regs[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4560_ (.CLK(clknet_leaf_41_clk),
    .D(_0220_),
    .Q(\as1802.regs[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4561_ (.CLK(clknet_leaf_42_clk),
    .D(_0221_),
    .Q(\as1802.regs[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4562_ (.CLK(clknet_leaf_40_clk),
    .D(_0222_),
    .Q(\as1802.regs[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4563_ (.CLK(clknet_leaf_39_clk),
    .D(_0223_),
    .Q(\as1802.regs[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4564_ (.CLK(clknet_leaf_46_clk),
    .D(_0224_),
    .Q(\as1802.regs[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4565_ (.CLK(clknet_leaf_49_clk),
    .D(_0225_),
    .Q(\as1802.regs[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4566_ (.CLK(clknet_leaf_48_clk),
    .D(_0226_),
    .Q(\as1802.regs[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4567_ (.CLK(clknet_leaf_38_clk),
    .D(_0227_),
    .Q(\as1802.regs[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4568_ (.CLK(clknet_leaf_40_clk),
    .D(_0228_),
    .Q(\as1802.regs[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4569_ (.CLK(clknet_leaf_42_clk),
    .D(_0229_),
    .Q(\as1802.regs[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4570_ (.CLK(clknet_leaf_40_clk),
    .D(_0230_),
    .Q(\as1802.regs[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4571_ (.CLK(clknet_leaf_39_clk),
    .D(_0231_),
    .Q(\as1802.regs[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4572_ (.CLK(clknet_leaf_50_clk),
    .D(_0232_),
    .Q(\as1802.regs[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4573_ (.CLK(clknet_leaf_2_clk),
    .D(_0233_),
    .Q(\as1802.regs[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4574_ (.CLK(clknet_leaf_6_clk),
    .D(_0234_),
    .Q(\as1802.regs[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4575_ (.CLK(clknet_leaf_45_clk),
    .D(_0235_),
    .Q(\as1802.regs[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4576_ (.CLK(clknet_leaf_1_clk),
    .D(_0236_),
    .Q(\as1802.regs[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4577_ (.CLK(clknet_leaf_51_clk),
    .D(_0237_),
    .Q(\as1802.regs[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4578_ (.CLK(clknet_leaf_49_clk),
    .D(_0238_),
    .Q(\as1802.regs[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4579_ (.CLK(clknet_leaf_51_clk),
    .D(_0239_),
    .Q(\as1802.regs[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4580_ (.CLK(clknet_leaf_46_clk),
    .D(_0240_),
    .Q(\as1802.regs[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4581_ (.CLK(clknet_leaf_49_clk),
    .D(_0241_),
    .Q(\as1802.regs[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4582_ (.CLK(clknet_leaf_41_clk),
    .D(_0242_),
    .Q(\as1802.regs[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4583_ (.CLK(clknet_leaf_37_clk),
    .D(_0243_),
    .Q(\as1802.regs[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4584_ (.CLK(clknet_leaf_42_clk),
    .D(_0244_),
    .Q(\as1802.regs[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4585_ (.CLK(clknet_leaf_31_clk),
    .D(_0245_),
    .Q(\as1802.regs[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4586_ (.CLK(clknet_leaf_39_clk),
    .D(_0246_),
    .Q(\as1802.regs[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4587_ (.CLK(clknet_leaf_36_clk),
    .D(_0247_),
    .Q(\as1802.regs[11][15] ));
 sky130_fd_sc_hd__dfxtp_4 _4588_ (.CLK(clknet_leaf_26_clk),
    .D(_0248_),
    .Q(\as1802.mem_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4589_ (.CLK(clknet_leaf_26_clk),
    .D(_0249_),
    .Q(\as1802.mem_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_4 _4590_ (.CLK(clknet_leaf_26_clk),
    .D(_0250_),
    .Q(\as1802.mem_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4591_ (.CLK(clknet_leaf_30_clk),
    .D(_0251_),
    .Q(\as1802.addr_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4592_ (.CLK(clknet_leaf_30_clk),
    .D(_0252_),
    .Q(\as1802.addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4593_ (.CLK(clknet_leaf_30_clk),
    .D(_0253_),
    .Q(\as1802.addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4594_ (.CLK(clknet_leaf_27_clk),
    .D(_0254_),
    .Q(\as1802.addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4595_ (.CLK(clknet_leaf_28_clk),
    .D(_0255_),
    .Q(\as1802.addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4596_ (.CLK(clknet_leaf_30_clk),
    .D(_0256_),
    .Q(\as1802.addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4597_ (.CLK(clknet_leaf_28_clk),
    .D(_0257_),
    .Q(\as1802.addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4598_ (.CLK(clknet_leaf_33_clk),
    .D(_0258_),
    .Q(\as1802.addr_buff[7] ));
 sky130_fd_sc_hd__dfxtp_2 _4599_ (.CLK(clknet_leaf_32_clk),
    .D(_0259_),
    .Q(\as1802.addr_buff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4600_ (.CLK(clknet_leaf_30_clk),
    .D(_0260_),
    .Q(\as1802.addr_buff[9] ));
 sky130_fd_sc_hd__dfxtp_2 _4601_ (.CLK(clknet_leaf_32_clk),
    .D(_0261_),
    .Q(\as1802.addr_buff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4602_ (.CLK(clknet_leaf_32_clk),
    .D(_0262_),
    .Q(\as1802.addr_buff[11] ));
 sky130_fd_sc_hd__dfxtp_2 _4603_ (.CLK(clknet_leaf_33_clk),
    .D(_0263_),
    .Q(\as1802.addr_buff[12] ));
 sky130_fd_sc_hd__dfxtp_2 _4604_ (.CLK(clknet_leaf_32_clk),
    .D(_0264_),
    .Q(\as1802.addr_buff[13] ));
 sky130_fd_sc_hd__dfxtp_2 _4605_ (.CLK(clknet_leaf_32_clk),
    .D(_0265_),
    .Q(\as1802.addr_buff[14] ));
 sky130_fd_sc_hd__dfxtp_2 _4606_ (.CLK(clknet_leaf_30_clk),
    .D(_0266_),
    .Q(\as1802.addr_buff[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4607_ (.CLK(clknet_leaf_32_clk),
    .D(_0267_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _4608_ (.CLK(clknet_leaf_29_clk),
    .D(_0268_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _4609_ (.CLK(clknet_leaf_29_clk),
    .D(_0269_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _4610_ (.CLK(clknet_leaf_28_clk),
    .D(_0270_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _4611_ (.CLK(clknet_leaf_28_clk),
    .D(_0271_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _4612_ (.CLK(clknet_leaf_28_clk),
    .D(_0272_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _4613_ (.CLK(clknet_leaf_27_clk),
    .D(_0273_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _4614_ (.CLK(clknet_leaf_26_clk),
    .D(_0274_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_4 _4615_ (.CLK(clknet_leaf_18_clk),
    .D(_0275_),
    .Q(\as1802.instr_latch[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4616_ (.CLK(clknet_leaf_18_clk),
    .D(_0276_),
    .Q(\as1802.instr_latch[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4617_ (.CLK(clknet_leaf_18_clk),
    .D(_0277_),
    .Q(\as1802.instr_latch[2] ));
 sky130_fd_sc_hd__dfxtp_4 _4618_ (.CLK(clknet_leaf_18_clk),
    .D(_0278_),
    .Q(\as1802.cond_inv ));
 sky130_fd_sc_hd__dfxtp_4 _4619_ (.CLK(clknet_leaf_19_clk),
    .D(_0279_),
    .Q(\as1802.instr_latch[4] ));
 sky130_fd_sc_hd__dfxtp_2 _4620_ (.CLK(clknet_leaf_22_clk),
    .D(_0280_),
    .Q(\as1802.instr_latch[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4621_ (.CLK(clknet_leaf_22_clk),
    .D(_0281_),
    .Q(\as1802.instr_latch[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4622_ (.CLK(clknet_leaf_22_clk),
    .D(_0282_),
    .Q(\as1802.instr_latch[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4623_ (.CLK(clknet_leaf_30_clk),
    .D(_0283_),
    .Q(\as1802.last_hi_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4624_ (.CLK(clknet_leaf_32_clk),
    .D(_0284_),
    .Q(\as1802.last_hi_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4625_ (.CLK(clknet_leaf_28_clk),
    .D(_0285_),
    .Q(\as1802.last_hi_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4626_ (.CLK(clknet_leaf_30_clk),
    .D(_0286_),
    .Q(\as1802.last_hi_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4627_ (.CLK(clknet_leaf_33_clk),
    .D(_0287_),
    .Q(\as1802.last_hi_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4628_ (.CLK(clknet_leaf_29_clk),
    .D(_0288_),
    .Q(\as1802.last_hi_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4629_ (.CLK(clknet_leaf_28_clk),
    .D(_0289_),
    .Q(\as1802.last_hi_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4630_ (.CLK(clknet_leaf_29_clk),
    .D(_0290_),
    .Q(\as1802.last_hi_addr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _4631_ (.CLK(clknet_leaf_25_clk),
    .D(_0291_),
    .Q(\as1802.will_interrupt ));
 sky130_fd_sc_hd__dfxtp_4 _4632_ (.CLK(clknet_leaf_25_clk),
    .D(_0292_),
    .Q(\as1802.IE ));
 sky130_fd_sc_hd__dfxtp_1 _4633_ (.CLK(clknet_leaf_25_clk),
    .D(_0293_),
    .Q(\as1802.idle ));
 sky130_fd_sc_hd__dfxtp_1 _4634_ (.CLK(clknet_leaf_25_clk),
    .D(_0294_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _4635_ (.CLK(clknet_leaf_26_clk),
    .D(_0295_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _4636_ (.CLK(clknet_leaf_26_clk),
    .D(_0296_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_2 _4637_ (.CLK(clknet_leaf_24_clk),
    .D(_0297_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _4638_ (.CLK(clknet_leaf_24_clk),
    .D(_0008_),
    .Q(\as1802.EF_l[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4639_ (.CLK(clknet_leaf_24_clk),
    .D(_0009_),
    .Q(\as1802.EF_l[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4640_ (.CLK(clknet_leaf_24_clk),
    .D(_0010_),
    .Q(\as1802.EF_l[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4641_ (.CLK(clknet_leaf_25_clk),
    .D(_0011_),
    .Q(\as1802.EF_l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4642_ (.CLK(clknet_leaf_25_clk),
    .D(_0298_),
    .Q(\as1802.lda ));
 sky130_fd_sc_hd__dfxtp_4 _4643_ (.CLK(clknet_leaf_24_clk),
    .D(_0299_),
    .Q(\as1802.DF ));
 sky130_fd_sc_hd__dfxtp_4 _4644_ (.CLK(clknet_leaf_21_clk),
    .D(_0300_),
    .Q(\as1802.X[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4645_ (.CLK(clknet_leaf_20_clk),
    .D(_0301_),
    .Q(\as1802.X[1] ));
 sky130_fd_sc_hd__dfxtp_4 _4646_ (.CLK(clknet_leaf_21_clk),
    .D(_0302_),
    .Q(\as1802.X[2] ));
 sky130_fd_sc_hd__dfxtp_4 _4647_ (.CLK(clknet_leaf_21_clk),
    .D(_0303_),
    .Q(\as1802.X[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4648_ (.CLK(clknet_leaf_16_clk),
    .D(_0304_),
    .Q(\as1802.T[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4649_ (.CLK(clknet_leaf_16_clk),
    .D(_0305_),
    .Q(\as1802.T[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4650_ (.CLK(clknet_leaf_16_clk),
    .D(_0306_),
    .Q(\as1802.T[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4651_ (.CLK(clknet_leaf_17_clk),
    .D(_0307_),
    .Q(\as1802.T[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4652_ (.CLK(clknet_leaf_16_clk),
    .D(_0308_),
    .Q(\as1802.T[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4653_ (.CLK(clknet_leaf_19_clk),
    .D(_0309_),
    .Q(\as1802.T[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4654_ (.CLK(clknet_leaf_20_clk),
    .D(_0310_),
    .Q(\as1802.T[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4655_ (.CLK(clknet_leaf_20_clk),
    .D(_0311_),
    .Q(\as1802.T[7] ));
 sky130_fd_sc_hd__dfxtp_2 _4656_ (.CLK(clknet_leaf_16_clk),
    .D(_0312_),
    .Q(\as1802.D[0] ));
 sky130_fd_sc_hd__dfxtp_4 _4657_ (.CLK(clknet_leaf_18_clk),
    .D(_0313_),
    .Q(\as1802.D[1] ));
 sky130_fd_sc_hd__dfxtp_4 _4658_ (.CLK(clknet_leaf_18_clk),
    .D(_0314_),
    .Q(\as1802.D[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4659_ (.CLK(clknet_leaf_18_clk),
    .D(_0315_),
    .Q(\as1802.D[3] ));
 sky130_fd_sc_hd__dfxtp_2 _4660_ (.CLK(clknet_leaf_19_clk),
    .D(_0316_),
    .Q(\as1802.D[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4661_ (.CLK(clknet_leaf_20_clk),
    .D(_0317_),
    .Q(\as1802.D[5] ));
 sky130_fd_sc_hd__dfxtp_4 _4662_ (.CLK(clknet_2_3__leaf_clk),
    .D(_0318_),
    .Q(\as1802.D[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4663_ (.CLK(clknet_leaf_22_clk),
    .D(_0319_),
    .Q(\as1802.D[7] ));
 sky130_fd_sc_hd__dfxtp_2 _4664_ (.CLK(clknet_leaf_19_clk),
    .D(_0320_),
    .Q(\as1802.P[0] ));
 sky130_fd_sc_hd__dfxtp_4 _4665_ (.CLK(clknet_leaf_21_clk),
    .D(_0321_),
    .Q(\as1802.P[1] ));
 sky130_fd_sc_hd__dfxtp_2 _4666_ (.CLK(clknet_leaf_16_clk),
    .D(_0322_),
    .Q(\as1802.P[2] ));
 sky130_fd_sc_hd__dfxtp_4 _4667_ (.CLK(clknet_leaf_16_clk),
    .D(_0323_),
    .Q(\as1802.P[3] ));
 sky130_fd_sc_hd__dfxtp_4 _4668_ (.CLK(clknet_leaf_19_clk),
    .D(_0324_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_4 _4669_ (.CLK(clknet_leaf_18_clk),
    .D(_0325_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_4 _4670_ (.CLK(clknet_leaf_18_clk),
    .D(_0326_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_4 _4671_ (.CLK(clknet_leaf_18_clk),
    .D(_0327_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_4 _4672_ (.CLK(clknet_leaf_19_clk),
    .D(_0328_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_4 _4673_ (.CLK(clknet_leaf_20_clk),
    .D(_0329_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_4 _4674_ (.CLK(clknet_leaf_22_clk),
    .D(_0330_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_4 _4675_ (.CLK(clknet_leaf_32_clk),
    .D(_0331_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _4676_ (.CLK(clknet_leaf_45_clk),
    .D(_0332_),
    .Q(\as1802.regs[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4677_ (.CLK(clknet_leaf_48_clk),
    .D(_0333_),
    .Q(\as1802.regs[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4678_ (.CLK(clknet_leaf_48_clk),
    .D(_0334_),
    .Q(\as1802.regs[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4679_ (.CLK(clknet_leaf_37_clk),
    .D(_0335_),
    .Q(\as1802.regs[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4680_ (.CLK(clknet_leaf_39_clk),
    .D(_0336_),
    .Q(\as1802.regs[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4681_ (.CLK(clknet_leaf_43_clk),
    .D(_0337_),
    .Q(\as1802.regs[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4682_ (.CLK(clknet_leaf_38_clk),
    .D(_0338_),
    .Q(\as1802.regs[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4683_ (.CLK(clknet_leaf_39_clk),
    .D(_0339_),
    .Q(\as1802.regs[9][15] ));
 sky130_fd_sc_hd__dfxtp_4 _4684_ (.CLK(clknet_leaf_8_clk),
    .D(_0340_),
    .Q(\as1802.regs[2][8] ));
 sky130_fd_sc_hd__dfxtp_2 _4685_ (.CLK(clknet_leaf_45_clk),
    .D(_0341_),
    .Q(\as1802.regs[2][9] ));
 sky130_fd_sc_hd__dfxtp_2 _4686_ (.CLK(clknet_leaf_44_clk),
    .D(_0342_),
    .Q(\as1802.regs[2][10] ));
 sky130_fd_sc_hd__dfxtp_2 _4687_ (.CLK(clknet_leaf_35_clk),
    .D(_0343_),
    .Q(\as1802.regs[2][11] ));
 sky130_fd_sc_hd__dfxtp_2 _4688_ (.CLK(clknet_leaf_44_clk),
    .D(_0344_),
    .Q(\as1802.regs[2][12] ));
 sky130_fd_sc_hd__dfxtp_2 _4689_ (.CLK(clknet_leaf_31_clk),
    .D(_0345_),
    .Q(\as1802.regs[2][13] ));
 sky130_fd_sc_hd__dfxtp_2 _4690_ (.CLK(clknet_leaf_34_clk),
    .D(_0346_),
    .Q(\as1802.regs[2][14] ));
 sky130_fd_sc_hd__dfxtp_2 _4691_ (.CLK(clknet_leaf_32_clk),
    .D(_0347_),
    .Q(\as1802.regs[2][15] ));
 sky130_fd_sc_hd__dfxtp_2 _4692_ (.CLK(clknet_leaf_26_clk),
    .D(_0348_),
    .Q(\as1802.mem_write ));
 sky130_fd_sc_hd__dfxtp_1 _4693_ (.CLK(clknet_leaf_45_clk),
    .D(_0349_),
    .Q(\as1802.regs[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4694_ (.CLK(clknet_leaf_45_clk),
    .D(_0350_),
    .Q(\as1802.regs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4695_ (.CLK(clknet_leaf_47_clk),
    .D(_0351_),
    .Q(\as1802.regs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4696_ (.CLK(clknet_leaf_34_clk),
    .D(_0352_),
    .Q(\as1802.regs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4697_ (.CLK(clknet_leaf_44_clk),
    .D(_0353_),
    .Q(\as1802.regs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4698_ (.CLK(clknet_leaf_35_clk),
    .D(_0354_),
    .Q(\as1802.regs[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4699_ (.CLK(clknet_leaf_33_clk),
    .D(_0355_),
    .Q(\as1802.regs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4700_ (.CLK(clknet_leaf_33_clk),
    .D(_0356_),
    .Q(\as1802.regs[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4701_ (.CLK(clknet_leaf_25_clk),
    .D(_0357_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _4702_ (.CLK(clknet_leaf_25_clk),
    .D(_0358_),
    .Q(net31));
 sky130_fd_sc_hd__clkbuf_2 _4708_ (.A(net15),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_opt_1_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_opt_1_0_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_opt_1_0_clk));
 sky130_fd_sc_hd__buf_4 fanout100 (.A(net111),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_8 fanout101 (.A(net104),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_8 fanout102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_6 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__buf_6 fanout104 (.A(net111),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__buf_6 fanout106 (.A(net110),
    .X(net106));
 sky130_fd_sc_hd__buf_6 fanout107 (.A(net109),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_6 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_6 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__buf_6 fanout111 (.A(_2166_),
    .X(net111));
 sky130_fd_sc_hd__buf_6 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_6 fanout113 (.A(net118),
    .X(net113));
 sky130_fd_sc_hd__buf_6 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_8 fanout115 (.A(net118),
    .X(net115));
 sky130_fd_sc_hd__buf_6 fanout116 (.A(net118),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_6 fanout118 (.A(_2163_),
    .X(net118));
 sky130_fd_sc_hd__buf_6 fanout119 (.A(net125),
    .X(net119));
 sky130_fd_sc_hd__buf_6 fanout120 (.A(net125),
    .X(net120));
 sky130_fd_sc_hd__buf_6 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net125),
    .X(net122));
 sky130_fd_sc_hd__buf_6 fanout123 (.A(net125),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_8 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_8 fanout125 (.A(_2162_),
    .X(net125));
 sky130_fd_sc_hd__buf_6 fanout126 (.A(_2149_),
    .X(net126));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(_2149_),
    .X(net127));
 sky130_fd_sc_hd__buf_6 fanout128 (.A(_2095_),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(_2095_),
    .X(net129));
 sky130_fd_sc_hd__buf_6 fanout130 (.A(_2094_),
    .X(net130));
 sky130_fd_sc_hd__buf_4 fanout131 (.A(_2094_),
    .X(net131));
 sky130_fd_sc_hd__buf_4 fanout132 (.A(_2057_),
    .X(net132));
 sky130_fd_sc_hd__buf_6 fanout133 (.A(_2055_),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_8 fanout134 (.A(_2048_),
    .X(net134));
 sky130_fd_sc_hd__buf_6 fanout135 (.A(_1303_),
    .X(net135));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(_1302_),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(_1302_),
    .X(net137));
 sky130_fd_sc_hd__buf_4 fanout138 (.A(_1301_),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net141),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 fanout140 (.A(net141),
    .X(net140));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(net146),
    .X(net141));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_4 fanout143 (.A(net146),
    .X(net143));
 sky130_fd_sc_hd__buf_4 fanout144 (.A(net146),
    .X(net144));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_4 fanout146 (.A(_2165_),
    .X(net146));
 sky130_fd_sc_hd__buf_4 fanout147 (.A(net149),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_2 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__buf_4 fanout149 (.A(net154),
    .X(net149));
 sky130_fd_sc_hd__buf_4 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__buf_4 fanout151 (.A(net154),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net154),
    .X(net152));
 sky130_fd_sc_hd__buf_2 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__buf_4 fanout154 (.A(_2164_),
    .X(net154));
 sky130_fd_sc_hd__buf_6 fanout155 (.A(_2139_),
    .X(net155));
 sky130_fd_sc_hd__buf_6 fanout156 (.A(_2138_),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_8 fanout157 (.A(_1551_),
    .X(net157));
 sky130_fd_sc_hd__buf_6 fanout158 (.A(_1207_),
    .X(net158));
 sky130_fd_sc_hd__buf_6 fanout159 (.A(_1205_),
    .X(net159));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(_1205_),
    .X(net160));
 sky130_fd_sc_hd__buf_8 fanout161 (.A(_1204_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(_1204_),
    .X(net162));
 sky130_fd_sc_hd__buf_6 fanout163 (.A(_0628_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_8 fanout164 (.A(_0413_),
    .X(net164));
 sky130_fd_sc_hd__buf_6 fanout165 (.A(_0379_),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_8 fanout166 (.A(net168),
    .X(net166));
 sky130_fd_sc_hd__buf_6 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_8 fanout168 (.A(_2093_),
    .X(net168));
 sky130_fd_sc_hd__buf_6 fanout169 (.A(_1969_),
    .X(net169));
 sky130_fd_sc_hd__buf_4 fanout170 (.A(net172),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__buf_4 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_6 fanout173 (.A(_1969_),
    .X(net173));
 sky130_fd_sc_hd__buf_6 fanout174 (.A(net177),
    .X(net174));
 sky130_fd_sc_hd__buf_8 fanout175 (.A(net177),
    .X(net175));
 sky130_fd_sc_hd__buf_8 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__buf_6 fanout177 (.A(_1968_),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_8 fanout178 (.A(_1552_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 fanout179 (.A(_1498_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 fanout180 (.A(_1498_),
    .X(net180));
 sky130_fd_sc_hd__buf_6 fanout181 (.A(_1494_),
    .X(net181));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(_1484_),
    .X(net182));
 sky130_fd_sc_hd__buf_6 fanout183 (.A(_2156_),
    .X(net183));
 sky130_fd_sc_hd__buf_6 fanout184 (.A(_2046_),
    .X(net184));
 sky130_fd_sc_hd__buf_6 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(_2028_),
    .X(net187));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(_1954_),
    .X(net188));
 sky130_fd_sc_hd__buf_6 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_16 fanout190 (.A(_1951_),
    .X(net190));
 sky130_fd_sc_hd__buf_6 fanout191 (.A(_2036_),
    .X(net191));
 sky130_fd_sc_hd__buf_6 fanout192 (.A(net194),
    .X(net192));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__buf_6 fanout194 (.A(_1934_),
    .X(net194));
 sky130_fd_sc_hd__buf_6 fanout195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__buf_6 fanout196 (.A(_1933_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_16 fanout197 (.A(_1932_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_16 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__buf_12 fanout199 (.A(_1931_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_16 fanout200 (.A(_1927_),
    .X(net200));
 sky130_fd_sc_hd__buf_12 fanout201 (.A(_1927_),
    .X(net201));
 sky130_fd_sc_hd__buf_12 fanout202 (.A(_1926_),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_16 fanout203 (.A(_1912_),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(net37),
    .X(net204));
 sky130_fd_sc_hd__buf_6 fanout205 (.A(net36),
    .X(net205));
 sky130_fd_sc_hd__buf_8 fanout206 (.A(net32),
    .X(net206));
 sky130_fd_sc_hd__buf_6 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__buf_4 fanout208 (.A(net24),
    .X(net208));
 sky130_fd_sc_hd__buf_6 fanout209 (.A(net16),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_8 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 fanout211 (.A(\as1802.D[7] ),
    .X(net211));
 sky130_fd_sc_hd__buf_6 fanout212 (.A(\as1802.D[5] ),
    .X(net212));
 sky130_fd_sc_hd__buf_6 fanout213 (.A(\as1802.D[4] ),
    .X(net213));
 sky130_fd_sc_hd__buf_6 fanout214 (.A(\as1802.D[3] ),
    .X(net214));
 sky130_fd_sc_hd__buf_6 fanout215 (.A(\as1802.D[2] ),
    .X(net215));
 sky130_fd_sc_hd__buf_8 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(\as1802.D[1] ),
    .X(net217));
 sky130_fd_sc_hd__buf_6 fanout218 (.A(\as1802.D[0] ),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(\as1802.D[0] ),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_8 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__buf_6 fanout221 (.A(\as1802.instr_latch[7] ),
    .X(net221));
 sky130_fd_sc_hd__buf_6 fanout222 (.A(\as1802.instr_latch[6] ),
    .X(net222));
 sky130_fd_sc_hd__buf_2 fanout223 (.A(\as1802.instr_latch[6] ),
    .X(net223));
 sky130_fd_sc_hd__buf_8 fanout224 (.A(\as1802.instr_latch[5] ),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_6 fanout226 (.A(\as1802.cond_inv ),
    .X(net226));
 sky130_fd_sc_hd__buf_4 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__buf_6 fanout228 (.A(\as1802.cond_inv ),
    .X(net228));
 sky130_fd_sc_hd__buf_8 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__buf_8 fanout230 (.A(\as1802.cond_inv ),
    .X(net230));
 sky130_fd_sc_hd__buf_8 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__buf_8 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_6 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(\as1802.instr_latch[2] ),
    .X(net234));
 sky130_fd_sc_hd__buf_8 fanout235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__buf_12 fanout236 (.A(\as1802.instr_latch[1] ),
    .X(net236));
 sky130_fd_sc_hd__buf_12 fanout237 (.A(\as1802.instr_latch[0] ),
    .X(net237));
 sky130_fd_sc_hd__buf_6 fanout238 (.A(\as1802.mem_cycle[1] ),
    .X(net238));
 sky130_fd_sc_hd__buf_12 fanout239 (.A(net241),
    .X(net239));
 sky130_fd_sc_hd__buf_8 fanout240 (.A(net241),
    .X(net240));
 sky130_fd_sc_hd__buf_12 fanout241 (.A(_0003_),
    .X(net241));
 sky130_fd_sc_hd__buf_6 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__buf_12 fanout243 (.A(_0002_),
    .X(net243));
 sky130_fd_sc_hd__buf_6 fanout244 (.A(_0002_),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_8 fanout245 (.A(net248),
    .X(net245));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net248),
    .X(net246));
 sky130_fd_sc_hd__buf_6 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__buf_4 fanout248 (.A(_0001_),
    .X(net248));
 sky130_fd_sc_hd__buf_6 fanout249 (.A(net251),
    .X(net249));
 sky130_fd_sc_hd__buf_4 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(_0001_),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_8 fanout252 (.A(net255),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_8 fanout253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__buf_4 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(_0001_),
    .X(net255));
 sky130_fd_sc_hd__buf_6 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_6 fanout257 (.A(net263),
    .X(net257));
 sky130_fd_sc_hd__buf_6 fanout258 (.A(net263),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 fanout259 (.A(net263),
    .X(net259));
 sky130_fd_sc_hd__buf_8 fanout260 (.A(net262),
    .X(net260));
 sky130_fd_sc_hd__buf_6 fanout261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__buf_6 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__buf_4 fanout263 (.A(_0000_),
    .X(net263));
 sky130_fd_sc_hd__buf_6 fanout264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__buf_4 fanout265 (.A(_0000_),
    .X(net265));
 sky130_fd_sc_hd__buf_6 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__buf_8 fanout267 (.A(_0000_),
    .X(net267));
 sky130_fd_sc_hd__buf_6 fanout268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__buf_4 fanout269 (.A(\as1802.instr_cycle[2] ),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_8 fanout270 (.A(net274),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(net274),
    .X(net271));
 sky130_fd_sc_hd__buf_4 fanout272 (.A(net274),
    .X(net272));
 sky130_fd_sc_hd__buf_2 fanout273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__buf_8 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(\as1802.instr_cycle[0] ),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_4 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_4 fanout277 (.A(_1928_),
    .X(net277));
 sky130_fd_sc_hd__buf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 fanout279 (.A(_1928_),
    .X(net279));
 sky130_fd_sc_hd__buf_8 fanout280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__buf_6 fanout281 (.A(net14),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_16 fanout282 (.A(net14),
    .X(net282));
 sky130_fd_sc_hd__buf_4 fanout38 (.A(_1189_),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 fanout39 (.A(_1189_),
    .X(net39));
 sky130_fd_sc_hd__buf_4 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(_1134_),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(_1084_),
    .X(net42));
 sky130_fd_sc_hd__buf_2 fanout43 (.A(_1084_),
    .X(net43));
 sky130_fd_sc_hd__buf_4 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 fanout45 (.A(_1028_),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(_0980_),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(_0924_),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(_0872_),
    .X(net51));
 sky130_fd_sc_hd__buf_4 fanout52 (.A(_0819_),
    .X(net52));
 sky130_fd_sc_hd__buf_2 fanout53 (.A(_0819_),
    .X(net53));
 sky130_fd_sc_hd__buf_4 fanout54 (.A(_0757_),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(_0757_),
    .X(net55));
 sky130_fd_sc_hd__buf_4 fanout56 (.A(_0698_),
    .X(net56));
 sky130_fd_sc_hd__buf_2 fanout57 (.A(_0698_),
    .X(net57));
 sky130_fd_sc_hd__buf_4 fanout58 (.A(_0649_),
    .X(net58));
 sky130_fd_sc_hd__buf_2 fanout59 (.A(_0649_),
    .X(net59));
 sky130_fd_sc_hd__buf_6 fanout60 (.A(_0592_),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(_0592_),
    .X(net61));
 sky130_fd_sc_hd__buf_4 fanout62 (.A(_0534_),
    .X(net62));
 sky130_fd_sc_hd__buf_2 fanout63 (.A(_0534_),
    .X(net63));
 sky130_fd_sc_hd__buf_4 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 fanout65 (.A(_0478_),
    .X(net65));
 sky130_fd_sc_hd__buf_4 fanout66 (.A(_0427_),
    .X(net66));
 sky130_fd_sc_hd__buf_2 fanout67 (.A(_0427_),
    .X(net67));
 sky130_fd_sc_hd__buf_4 fanout68 (.A(_0377_),
    .X(net68));
 sky130_fd_sc_hd__buf_2 fanout69 (.A(_0377_),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(_0761_),
    .X(net71));
 sky130_fd_sc_hd__buf_4 fanout72 (.A(_2125_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 fanout73 (.A(_2125_),
    .X(net73));
 sky130_fd_sc_hd__buf_4 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__buf_2 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 fanout76 (.A(_1299_),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_8 fanout77 (.A(_1299_),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 fanout79 (.A(_0550_),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_8 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__buf_8 fanout81 (.A(_2078_),
    .X(net81));
 sky130_fd_sc_hd__buf_4 fanout82 (.A(_0374_),
    .X(net82));
 sky130_fd_sc_hd__buf_6 fanout83 (.A(_2090_),
    .X(net83));
 sky130_fd_sc_hd__buf_4 fanout84 (.A(_2090_),
    .X(net84));
 sky130_fd_sc_hd__buf_12 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_12 fanout86 (.A(_0362_),
    .X(net86));
 sky130_fd_sc_hd__buf_8 fanout87 (.A(_0361_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_8 fanout88 (.A(_0361_),
    .X(net88));
 sky130_fd_sc_hd__buf_8 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__buf_8 fanout90 (.A(net92),
    .X(net90));
 sky130_fd_sc_hd__buf_6 fanout91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__buf_8 fanout92 (.A(_2169_),
    .X(net92));
 sky130_fd_sc_hd__buf_8 fanout93 (.A(net95),
    .X(net93));
 sky130_fd_sc_hd__buf_6 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_16 fanout95 (.A(_2168_),
    .X(net95));
 sky130_fd_sc_hd__buf_6 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__buf_6 fanout97 (.A(net100),
    .X(net97));
 sky130_fd_sc_hd__buf_6 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__buf_6 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(io_in[6]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(io_in[7]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(io_in[8]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(io_in[9]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(rst),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(io_in[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(io_in[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(io_in[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(io_in[1]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[2]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(io_in[3]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(io_in[4]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(io_in[5]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 output15 (.A(net15),
    .X(io_oeb));
 sky130_fd_sc_hd__buf_4 output16 (.A(net16),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_4 output17 (.A(net17),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_4 output18 (.A(net18),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_4 output19 (.A(net19),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_4 output20 (.A(net20),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_4 output21 (.A(net21),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_4 output22 (.A(net22),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_4 output23 (.A(net23),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_4 output24 (.A(net24),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_4 output25 (.A(net25),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_4 output26 (.A(net26),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_4 output27 (.A(net27),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_4 output28 (.A(net28),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_4 output29 (.A(net29),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_4 output30 (.A(net30),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_4 output31 (.A(net31),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_4 output32 (.A(net32),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_4 output33 (.A(net33),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_4 output34 (.A(net34),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_4 output35 (.A(net35),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_4 output36 (.A(net36),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_4 output37 (.A(net37),
    .X(io_out[7]));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_283 (.LO(net283));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_284 (.LO(net284));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_285 (.LO(net285));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_286 (.LO(net286));
 sky130_fd_sc_hd__conb_1 wrapped_as1802_287 (.LO(net287));
 assign io_out[10] = net285;
 assign io_out[11] = net286;
 assign io_out[12] = net287;
 assign io_out[8] = net283;
 assign io_out[9] = net284;
endmodule

