VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tholin_avalonsemi_tbb1143
  CLASS BLOCK ;
  FOREIGN tholin_avalonsemi_tbb1143 ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 146.000 10.490 150.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 146.000 47.290 150.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 146.000 65.690 150.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 146.000 84.090 150.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 146.000 102.490 150.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 146.000 120.890 150.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 146.000 139.290 150.000 ;
    END
  END io_in[5]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 10.240 150.000 10.840 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 28.600 150.000 29.200 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 46.960 150.000 47.560 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 65.320 150.000 65.920 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 83.680 150.000 84.280 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 102.040 150.000 102.640 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 120.400 150.000 121.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 138.760 150.000 139.360 ;
    END
  END io_out[7]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 146.000 28.890 150.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.085 10.640 23.685 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.815 10.640 58.415 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.545 10.640 93.145 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.275 10.640 127.875 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.450 10.640 41.050 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.180 10.640 75.780 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.910 10.640 110.510 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.640 10.640 145.240 138.960 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 137.305 144.630 138.910 ;
        RECT 5.330 131.865 144.630 134.695 ;
        RECT 5.330 126.425 144.630 129.255 ;
        RECT 5.330 120.985 144.630 123.815 ;
        RECT 5.330 115.545 144.630 118.375 ;
        RECT 5.330 110.105 144.630 112.935 ;
        RECT 5.330 104.665 144.630 107.495 ;
        RECT 5.330 99.225 144.630 102.055 ;
        RECT 5.330 93.785 144.630 96.615 ;
        RECT 5.330 88.345 144.630 91.175 ;
        RECT 5.330 82.905 144.630 85.735 ;
        RECT 5.330 77.465 144.630 80.295 ;
        RECT 5.330 72.025 144.630 74.855 ;
        RECT 5.330 66.585 144.630 69.415 ;
        RECT 5.330 61.145 144.630 63.975 ;
        RECT 5.330 55.705 144.630 58.535 ;
        RECT 5.330 50.265 144.630 53.095 ;
        RECT 5.330 44.825 144.630 47.655 ;
        RECT 5.330 39.385 144.630 42.215 ;
        RECT 5.330 33.945 144.630 36.775 ;
        RECT 5.330 28.505 144.630 31.335 ;
        RECT 5.330 23.065 144.630 25.895 ;
        RECT 5.330 17.625 144.630 20.455 ;
        RECT 5.330 12.185 144.630 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 5.520 10.640 145.240 138.960 ;
      LAYER met2 ;
        RECT 7.920 145.720 9.930 146.610 ;
        RECT 10.770 145.720 28.330 146.610 ;
        RECT 29.170 145.720 46.730 146.610 ;
        RECT 47.570 145.720 65.130 146.610 ;
        RECT 65.970 145.720 83.530 146.610 ;
        RECT 84.370 145.720 101.930 146.610 ;
        RECT 102.770 145.720 120.330 146.610 ;
        RECT 121.170 145.720 138.730 146.610 ;
        RECT 139.570 145.720 145.210 146.610 ;
        RECT 7.920 10.695 145.210 145.720 ;
      LAYER met3 ;
        RECT 22.095 138.360 145.600 139.225 ;
        RECT 22.095 121.400 146.890 138.360 ;
        RECT 22.095 120.000 145.600 121.400 ;
        RECT 22.095 103.040 146.890 120.000 ;
        RECT 22.095 101.640 145.600 103.040 ;
        RECT 22.095 84.680 146.890 101.640 ;
        RECT 22.095 83.280 145.600 84.680 ;
        RECT 22.095 66.320 146.890 83.280 ;
        RECT 22.095 64.920 145.600 66.320 ;
        RECT 22.095 47.960 146.890 64.920 ;
        RECT 22.095 46.560 145.600 47.960 ;
        RECT 22.095 29.600 146.890 46.560 ;
        RECT 22.095 28.200 145.600 29.600 ;
        RECT 22.095 11.240 146.890 28.200 ;
        RECT 22.095 10.715 145.600 11.240 ;
  END
END tholin_avalonsemi_tbb1143
END LIBRARY

