VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO posit_unit
  CLASS BLOCK ;
  FOREIGN posit_unit ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END io_in[2]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 43.560 350.000 44.160 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 130.600 350.000 131.200 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 217.640 350.000 218.240 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 304.680 350.000 305.280 ;
    END
  END io_out[3]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 344.080 337.365 ;
      LAYER met1 ;
        RECT 4.670 10.640 345.390 337.520 ;
      LAYER met2 ;
        RECT 4.690 10.695 345.370 337.465 ;
      LAYER met3 ;
        RECT 4.000 313.840 346.000 337.445 ;
        RECT 4.400 312.440 346.000 313.840 ;
        RECT 4.000 305.680 346.000 312.440 ;
        RECT 4.000 304.280 345.600 305.680 ;
        RECT 4.000 244.480 346.000 304.280 ;
        RECT 4.400 243.080 346.000 244.480 ;
        RECT 4.000 218.640 346.000 243.080 ;
        RECT 4.000 217.240 345.600 218.640 ;
        RECT 4.000 175.120 346.000 217.240 ;
        RECT 4.400 173.720 346.000 175.120 ;
        RECT 4.000 131.600 346.000 173.720 ;
        RECT 4.000 130.200 345.600 131.600 ;
        RECT 4.000 105.760 346.000 130.200 ;
        RECT 4.400 104.360 346.000 105.760 ;
        RECT 4.000 44.560 346.000 104.360 ;
        RECT 4.000 43.160 345.600 44.560 ;
        RECT 4.000 36.400 346.000 43.160 ;
        RECT 4.400 35.000 346.000 36.400 ;
        RECT 4.000 10.715 346.000 35.000 ;
      LAYER met4 ;
        RECT 36.175 19.895 97.440 286.785 ;
        RECT 99.840 19.895 174.240 286.785 ;
        RECT 176.640 19.895 251.040 286.785 ;
        RECT 253.440 19.895 327.840 286.785 ;
        RECT 330.240 19.895 335.505 286.785 ;
  END
END posit_unit
END LIBRARY

