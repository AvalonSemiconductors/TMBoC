magic
tech sky130B
magscale 1 2
timestamp 1681463271
<< viali >>
rect 5181 61353 5215 61387
rect 44465 61353 44499 61387
rect 46857 61353 46891 61387
rect 49433 61353 49467 61387
rect 9689 61285 9723 61319
rect 11161 61285 11195 61319
rect 20729 61285 20763 61319
rect 22661 61285 22695 61319
rect 38485 61285 38519 61319
rect 43729 61285 43763 61319
rect 2237 61217 2271 61251
rect 10425 61217 10459 61251
rect 18153 61217 18187 61251
rect 35173 61217 35207 61251
rect 48053 61217 48087 61251
rect 1685 61149 1719 61183
rect 2789 61149 2823 61183
rect 4353 61149 4387 61183
rect 5089 61149 5123 61183
rect 5733 61149 5767 61183
rect 6653 61149 6687 61183
rect 7573 61149 7607 61183
rect 9505 61149 9539 61183
rect 10241 61149 10275 61183
rect 10977 61149 11011 61183
rect 11989 61149 12023 61183
rect 12725 61149 12759 61183
rect 14933 61149 14967 61183
rect 16129 61149 16163 61183
rect 17141 61149 17175 61183
rect 17969 61149 18003 61183
rect 18705 61149 18739 61183
rect 19809 61149 19843 61183
rect 20545 61149 20579 61183
rect 21281 61149 21315 61183
rect 22385 61149 22419 61183
rect 23857 61149 23891 61183
rect 25329 61149 25363 61183
rect 26249 61149 26283 61183
rect 27261 61149 27295 61183
rect 28273 61149 28307 61183
rect 29837 61149 29871 61183
rect 31217 61149 31251 61183
rect 32413 61149 32447 61183
rect 33333 61149 33367 61183
rect 33517 61149 33551 61183
rect 34989 61149 35023 61183
rect 36461 61149 36495 61183
rect 37565 61149 37599 61183
rect 38301 61149 38335 61183
rect 38945 61149 38979 61183
rect 40141 61149 40175 61183
rect 41613 61149 41647 61183
rect 42625 61149 42659 61183
rect 43545 61149 43579 61183
rect 44373 61149 44407 61183
rect 45293 61149 45327 61183
rect 46765 61149 46799 61183
rect 47869 61149 47903 61183
rect 48605 61149 48639 61183
rect 49341 61149 49375 61183
rect 50445 61149 50479 61183
rect 51365 61149 51399 61183
rect 52101 61149 52135 61183
rect 53205 61149 53239 61183
rect 54125 61149 54159 61183
rect 55505 61149 55539 61183
rect 56517 61149 56551 61183
rect 58173 61149 58207 61183
rect 3065 61081 3099 61115
rect 4537 61081 4571 61115
rect 6929 61081 6963 61115
rect 7849 61081 7883 61115
rect 13001 61081 13035 61115
rect 15209 61081 15243 61115
rect 16313 61081 16347 61115
rect 19993 61081 20027 61115
rect 24041 61081 24075 61115
rect 26433 61081 26467 61115
rect 34069 61081 34103 61115
rect 35725 61081 35759 61115
rect 35909 61081 35943 61115
rect 37749 61081 37783 61115
rect 40877 61081 40911 61115
rect 42901 61081 42935 61115
rect 46029 61081 46063 61115
rect 52285 61081 52319 61115
rect 53481 61081 53515 61115
rect 55781 61081 55815 61115
rect 58357 61081 58391 61115
rect 5917 61013 5951 61047
rect 12173 61013 12207 61047
rect 17325 61013 17359 61047
rect 18797 61013 18831 61047
rect 21373 61013 21407 61047
rect 25421 61013 25455 61047
rect 27353 61013 27387 61047
rect 28365 61013 28399 61047
rect 29929 61013 29963 61047
rect 31309 61013 31343 61047
rect 32505 61013 32539 61047
rect 34161 61013 34195 61047
rect 36553 61013 36587 61047
rect 39129 61013 39163 61047
rect 40233 61013 40267 61047
rect 40969 61013 41003 61047
rect 41705 61013 41739 61047
rect 45385 61013 45419 61047
rect 46121 61013 46155 61047
rect 48697 61013 48731 61047
rect 50537 61013 50571 61047
rect 51457 61013 51491 61047
rect 54309 61013 54343 61047
rect 56609 61013 56643 61047
rect 3249 60741 3283 60775
rect 3985 60741 4019 60775
rect 8401 60741 8435 60775
rect 13553 60741 13587 60775
rect 14289 60741 14323 60775
rect 15761 60741 15795 60775
rect 19441 60741 19475 60775
rect 22109 60741 22143 60775
rect 23489 60741 23523 60775
rect 24593 60741 24627 60775
rect 36369 60741 36403 60775
rect 41521 60741 41555 60775
rect 46673 60741 46707 60775
rect 50353 60741 50387 60775
rect 53021 60741 53055 60775
rect 1593 60673 1627 60707
rect 9045 60673 9079 60707
rect 23213 60673 23247 60707
rect 23397 60673 23431 60707
rect 23581 60673 23615 60707
rect 27537 60673 27571 60707
rect 29009 60673 29043 60707
rect 30481 60673 30515 60707
rect 54677 60673 54711 60707
rect 55413 60673 55447 60707
rect 56149 60673 56183 60707
rect 56885 60673 56919 60707
rect 58081 60673 58115 60707
rect 1869 60605 1903 60639
rect 8585 60605 8619 60639
rect 4169 60537 4203 60571
rect 14473 60537 14507 60571
rect 27721 60537 27755 60571
rect 30665 60537 30699 60571
rect 3341 60469 3375 60503
rect 9229 60469 9263 60503
rect 13645 60469 13679 60503
rect 15853 60469 15887 60503
rect 19533 60469 19567 60503
rect 22385 60469 22419 60503
rect 23765 60469 23799 60503
rect 24685 60469 24719 60503
rect 29101 60469 29135 60503
rect 30021 60469 30055 60503
rect 36461 60469 36495 60503
rect 41613 60469 41647 60503
rect 46765 60469 46799 60503
rect 50445 60469 50479 60503
rect 53113 60469 53147 60503
rect 54861 60469 54895 60503
rect 55597 60469 55631 60503
rect 56333 60469 56367 60503
rect 57069 60469 57103 60503
rect 58265 60469 58299 60503
rect 19993 60197 20027 60231
rect 21189 60197 21223 60231
rect 41245 60197 41279 60231
rect 17877 60129 17911 60163
rect 18337 60129 18371 60163
rect 42257 60129 42291 60163
rect 42717 60129 42751 60163
rect 2605 60061 2639 60095
rect 7389 60061 7423 60095
rect 7757 60061 7791 60095
rect 18061 60061 18095 60095
rect 18429 60061 18463 60095
rect 19441 60061 19475 60095
rect 19625 60061 19659 60095
rect 19717 60061 19751 60095
rect 19861 60061 19895 60095
rect 20637 60061 20671 60095
rect 21057 60061 21091 60095
rect 22201 60061 22235 60095
rect 22477 60061 22511 60095
rect 22569 60061 22603 60095
rect 22845 60061 22879 60095
rect 23029 60061 23063 60095
rect 23673 60061 23707 60095
rect 27813 60061 27847 60095
rect 28089 60061 28123 60095
rect 28182 60061 28216 60095
rect 28554 60061 28588 60095
rect 30640 60061 30674 60095
rect 30757 60061 30791 60095
rect 30977 60061 31011 60095
rect 31125 60061 31159 60095
rect 32413 60061 32447 60095
rect 32597 60061 32631 60095
rect 32965 60061 32999 60095
rect 33057 60061 33091 60095
rect 40693 60061 40727 60095
rect 40969 60061 41003 60095
rect 41113 60061 41147 60095
rect 42441 60061 42475 60095
rect 42809 60061 42843 60095
rect 56517 60061 56551 60095
rect 57253 60061 57287 60095
rect 57897 60061 57931 60095
rect 1685 59993 1719 60027
rect 2053 59993 2087 60027
rect 7573 59993 7607 60027
rect 7665 59993 7699 60027
rect 20821 59993 20855 60027
rect 20913 59993 20947 60027
rect 28365 59993 28399 60027
rect 28457 59993 28491 60027
rect 30113 59993 30147 60027
rect 30849 59993 30883 60027
rect 40877 59993 40911 60027
rect 41797 59993 41831 60027
rect 56701 59993 56735 60027
rect 58173 59993 58207 60027
rect 2697 59925 2731 59959
rect 7941 59925 7975 59959
rect 17693 59925 17727 59959
rect 21833 59925 21867 59959
rect 23857 59925 23891 59959
rect 28733 59925 28767 59959
rect 29101 59925 29135 59959
rect 30481 59925 30515 59959
rect 31677 59925 31711 59959
rect 32229 59925 32263 59959
rect 57345 59925 57379 59959
rect 57437 59721 57471 59755
rect 58265 59721 58299 59755
rect 2605 59653 2639 59687
rect 21097 59653 21131 59687
rect 22293 59653 22327 59687
rect 30113 59653 30147 59687
rect 57345 59653 57379 59687
rect 1685 59585 1719 59619
rect 20913 59585 20947 59619
rect 21189 59585 21223 59619
rect 21281 59585 21315 59619
rect 22109 59585 22143 59619
rect 22385 59585 22419 59619
rect 22529 59585 22563 59619
rect 23213 59585 23247 59619
rect 23397 59585 23431 59619
rect 23489 59585 23523 59619
rect 23586 59585 23620 59619
rect 28365 59585 28399 59619
rect 28641 59585 28675 59619
rect 29745 59585 29779 59619
rect 29838 59585 29872 59619
rect 30021 59585 30055 59619
rect 30210 59585 30244 59619
rect 43085 59585 43119 59619
rect 43269 59585 43303 59619
rect 43637 59585 43671 59619
rect 58081 59585 58115 59619
rect 42717 59517 42751 59551
rect 43545 59517 43579 59551
rect 21465 59449 21499 59483
rect 30389 59449 30423 59483
rect 1961 59381 1995 59415
rect 2697 59381 2731 59415
rect 22661 59381 22695 59415
rect 23765 59381 23799 59415
rect 29469 59381 29503 59415
rect 30665 59381 30699 59415
rect 57345 59177 57379 59211
rect 19993 59109 20027 59143
rect 41337 59041 41371 59075
rect 41797 59041 41831 59075
rect 1685 58973 1719 59007
rect 19441 58973 19475 59007
rect 19717 58973 19751 59007
rect 19861 58973 19895 59007
rect 41521 58973 41555 59007
rect 41889 58973 41923 59007
rect 57161 58973 57195 59007
rect 57897 58973 57931 59007
rect 19625 58905 19659 58939
rect 58173 58905 58207 58939
rect 1777 58837 1811 58871
rect 41153 58837 41187 58871
rect 58173 58565 58207 58599
rect 1593 58497 1627 58531
rect 35725 58497 35759 58531
rect 37933 58497 37967 58531
rect 38209 58497 38243 58531
rect 38301 58497 38335 58531
rect 38577 58497 38611 58531
rect 38853 58497 38887 58531
rect 41337 58497 41371 58531
rect 41521 58497 41555 58531
rect 41889 58497 41923 58531
rect 1869 58429 1903 58463
rect 36001 58429 36035 58463
rect 41797 58429 41831 58463
rect 37565 58293 37599 58327
rect 41153 58293 41187 58327
rect 58265 58293 58299 58327
rect 1593 57885 1627 57919
rect 35633 57885 35667 57919
rect 35725 57885 35759 57919
rect 36001 57885 36035 57919
rect 36277 57885 36311 57919
rect 36553 57885 36587 57919
rect 1869 57817 1903 57851
rect 35173 57817 35207 57851
rect 57989 57817 58023 57851
rect 58081 57749 58115 57783
rect 1593 57409 1627 57443
rect 1777 57205 1811 57239
rect 33333 56865 33367 56899
rect 32873 56797 32907 56831
rect 33057 56797 33091 56831
rect 33425 56797 33459 56831
rect 57897 56797 57931 56831
rect 1685 56729 1719 56763
rect 58173 56729 58207 56763
rect 1961 56661 1995 56695
rect 32689 56661 32723 56695
rect 58265 56457 58299 56491
rect 58173 56389 58207 56423
rect 41521 56321 41555 56355
rect 41889 56321 41923 56355
rect 41429 56253 41463 56287
rect 41797 56253 41831 56287
rect 41153 56117 41187 56151
rect 58357 55913 58391 55947
rect 25145 55777 25179 55811
rect 25237 55709 25271 55743
rect 25605 55709 25639 55743
rect 25697 55709 25731 55743
rect 30389 55709 30423 55743
rect 30481 55709 30515 55743
rect 30757 55709 30791 55743
rect 30849 55709 30883 55743
rect 1685 55641 1719 55675
rect 24593 55641 24627 55675
rect 29745 55641 29779 55675
rect 1777 55573 1811 55607
rect 1777 55369 1811 55403
rect 41153 55301 41187 55335
rect 1593 55233 1627 55267
rect 23765 55233 23799 55267
rect 24409 55233 24443 55267
rect 24777 55233 24811 55267
rect 24961 55233 24995 55267
rect 40877 55233 40911 55267
rect 41061 55233 41095 55267
rect 41250 55233 41284 55267
rect 41446 55233 41480 55267
rect 24317 55165 24351 55199
rect 23489 54621 23523 54655
rect 23581 54621 23615 54655
rect 23857 54621 23891 54655
rect 24041 54621 24075 54655
rect 58357 54621 58391 54655
rect 1685 54553 1719 54587
rect 22845 54553 22879 54587
rect 1777 54485 1811 54519
rect 1593 54145 1627 54179
rect 1777 53941 1811 53975
rect 40969 53669 41003 53703
rect 40417 53533 40451 53567
rect 40601 53533 40635 53567
rect 40837 53533 40871 53567
rect 40693 53465 40727 53499
rect 40049 53397 40083 53431
rect 23765 53125 23799 53159
rect 23857 53125 23891 53159
rect 1685 53057 1719 53091
rect 23581 53057 23615 53091
rect 23949 53057 23983 53091
rect 24593 53057 24627 53091
rect 24777 52989 24811 53023
rect 1777 52853 1811 52887
rect 24133 52853 24167 52887
rect 58357 52853 58391 52887
rect 24961 52649 24995 52683
rect 2053 52445 2087 52479
rect 1685 52377 1719 52411
rect 24685 52377 24719 52411
rect 21189 52105 21223 52139
rect 1869 52037 1903 52071
rect 8217 52037 8251 52071
rect 1685 51969 1719 52003
rect 8033 51969 8067 52003
rect 8309 51969 8343 52003
rect 21281 51969 21315 52003
rect 21005 51901 21039 51935
rect 20913 51833 20947 51867
rect 7849 51765 7883 51799
rect 20545 51765 20579 51799
rect 20821 51765 20855 51799
rect 58357 51357 58391 51391
rect 1685 51289 1719 51323
rect 1869 51289 1903 51323
rect 3893 50949 3927 50983
rect 3985 50949 4019 50983
rect 3709 50881 3743 50915
rect 4082 50881 4116 50915
rect 4261 50677 4295 50711
rect 57897 50269 57931 50303
rect 1685 50201 1719 50235
rect 1869 50201 1903 50235
rect 58173 50201 58207 50235
rect 1593 49793 1627 49827
rect 1777 49657 1811 49691
rect 1593 49181 1627 49215
rect 57989 49113 58023 49147
rect 58357 49113 58391 49147
rect 1777 49045 1811 49079
rect 1685 48705 1719 48739
rect 1869 48569 1903 48603
rect 2605 48229 2639 48263
rect 2053 48093 2087 48127
rect 2237 48093 2271 48127
rect 2426 48093 2460 48127
rect 57897 48093 57931 48127
rect 2329 48025 2363 48059
rect 58173 48025 58207 48059
rect 1685 47617 1719 47651
rect 58081 47617 58115 47651
rect 1777 47413 1811 47447
rect 58265 47413 58299 47447
rect 1777 47141 1811 47175
rect 1593 47005 1627 47039
rect 1593 46529 1627 46563
rect 1777 46325 1811 46359
rect 58173 45985 58207 46019
rect 57897 45917 57931 45951
rect 1685 45849 1719 45883
rect 1777 45781 1811 45815
rect 17509 45509 17543 45543
rect 36553 45509 36587 45543
rect 38209 45509 38243 45543
rect 38301 45509 38335 45543
rect 17141 45441 17175 45475
rect 17234 45441 17268 45475
rect 17417 45441 17451 45475
rect 17647 45441 17681 45475
rect 36369 45441 36403 45475
rect 36645 45441 36679 45475
rect 36737 45441 36771 45475
rect 38025 45441 38059 45475
rect 38445 45441 38479 45475
rect 58081 45441 58115 45475
rect 36921 45305 36955 45339
rect 38577 45305 38611 45339
rect 17785 45237 17819 45271
rect 58265 45237 58299 45271
rect 35449 45033 35483 45067
rect 1593 44829 1627 44863
rect 1869 44829 1903 44863
rect 34897 44829 34931 44863
rect 35081 44829 35115 44863
rect 35270 44829 35304 44863
rect 56977 44829 57011 44863
rect 57253 44829 57287 44863
rect 35173 44761 35207 44795
rect 57989 44761 58023 44795
rect 58265 44693 58299 44727
rect 1685 44353 1719 44387
rect 1869 44217 1903 44251
rect 34253 43877 34287 43911
rect 33701 43741 33735 43775
rect 34074 43741 34108 43775
rect 57897 43741 57931 43775
rect 1685 43673 1719 43707
rect 33885 43673 33919 43707
rect 33977 43673 34011 43707
rect 58173 43673 58207 43707
rect 1777 43605 1811 43639
rect 32597 43333 32631 43367
rect 1593 43265 1627 43299
rect 32321 43265 32355 43299
rect 32505 43265 32539 43299
rect 32694 43265 32728 43299
rect 1777 43061 1811 43095
rect 32873 43061 32907 43095
rect 33057 42653 33091 42687
rect 33149 42653 33183 42687
rect 33425 42653 33459 42687
rect 33701 42653 33735 42687
rect 33885 42653 33919 42687
rect 37289 42653 37323 42687
rect 37657 42653 37691 42687
rect 57069 42653 57103 42687
rect 32597 42585 32631 42619
rect 37473 42585 37507 42619
rect 37565 42585 37599 42619
rect 57989 42585 58023 42619
rect 58357 42585 58391 42619
rect 37841 42517 37875 42551
rect 57161 42517 57195 42551
rect 1593 42177 1627 42211
rect 1777 41973 1811 42007
rect 56977 41565 57011 41599
rect 57253 41565 57287 41599
rect 1685 41497 1719 41531
rect 2053 41497 2087 41531
rect 57989 41497 58023 41531
rect 58265 41429 58299 41463
rect 1685 41089 1719 41123
rect 1777 40885 1811 40919
rect 57897 40477 57931 40511
rect 1685 40409 1719 40443
rect 57069 40409 57103 40443
rect 58173 40409 58207 40443
rect 1777 40341 1811 40375
rect 57161 40341 57195 40375
rect 1685 40069 1719 40103
rect 21097 40069 21131 40103
rect 21189 40069 21223 40103
rect 20913 40001 20947 40035
rect 21281 40001 21315 40035
rect 1777 39797 1811 39831
rect 21465 39797 21499 39831
rect 2881 39525 2915 39559
rect 2329 39389 2363 39423
rect 2513 39389 2547 39423
rect 2605 39389 2639 39423
rect 2702 39389 2736 39423
rect 57069 39389 57103 39423
rect 1685 39321 1719 39355
rect 57989 39321 58023 39355
rect 58357 39321 58391 39355
rect 1777 39253 1811 39287
rect 57161 39253 57195 39287
rect 1685 38913 1719 38947
rect 22017 38913 22051 38947
rect 22293 38913 22327 38947
rect 22477 38845 22511 38879
rect 22109 38777 22143 38811
rect 23121 38777 23155 38811
rect 1777 38709 1811 38743
rect 20085 38505 20119 38539
rect 3065 38369 3099 38403
rect 2053 38301 2087 38335
rect 2421 38301 2455 38335
rect 3249 38301 3283 38335
rect 3433 38301 3467 38335
rect 20269 38301 20303 38335
rect 20361 38301 20395 38335
rect 22937 38301 22971 38335
rect 23085 38301 23119 38335
rect 23402 38301 23436 38335
rect 57897 38301 57931 38335
rect 2237 38233 2271 38267
rect 2329 38233 2363 38267
rect 20085 38233 20119 38267
rect 23213 38233 23247 38267
rect 23305 38233 23339 38267
rect 58173 38233 58207 38267
rect 2605 38165 2639 38199
rect 19809 38165 19843 38199
rect 20545 38165 20579 38199
rect 23581 38165 23615 38199
rect 20361 37961 20395 37995
rect 21005 37961 21039 37995
rect 23305 37961 23339 37995
rect 19714 37893 19748 37927
rect 22937 37893 22971 37927
rect 23765 37893 23799 37927
rect 25237 37893 25271 37927
rect 1685 37825 1719 37859
rect 16957 37825 16991 37859
rect 19349 37825 19383 37859
rect 19469 37825 19503 37859
rect 19625 37825 19659 37859
rect 19855 37825 19889 37859
rect 20821 37825 20855 37859
rect 21097 37825 21131 37859
rect 22753 37825 22787 37859
rect 23029 37825 23063 37859
rect 23121 37825 23155 37859
rect 23995 37825 24029 37859
rect 24961 37825 24995 37859
rect 25145 37825 25179 37859
rect 25329 37825 25363 37859
rect 58081 37825 58115 37859
rect 17509 37757 17543 37791
rect 22477 37757 22511 37791
rect 24133 37757 24167 37791
rect 1869 37689 1903 37723
rect 23930 37689 23964 37723
rect 25513 37689 25547 37723
rect 19993 37621 20027 37655
rect 20637 37621 20671 37655
rect 24225 37621 24259 37655
rect 58265 37621 58299 37655
rect 21097 37281 21131 37315
rect 5917 37213 5951 37247
rect 6009 37213 6043 37247
rect 6285 37213 6319 37247
rect 6561 37213 6595 37247
rect 6745 37213 6779 37247
rect 19625 37213 19659 37247
rect 20821 37213 20855 37247
rect 53757 37213 53791 37247
rect 54130 37213 54164 37247
rect 57897 37213 57931 37247
rect 20177 37145 20211 37179
rect 53941 37145 53975 37179
rect 54033 37145 54067 37179
rect 58173 37145 58207 37179
rect 5549 37077 5583 37111
rect 54317 37077 54351 37111
rect 18797 36805 18831 36839
rect 23489 36805 23523 36839
rect 23765 36805 23799 36839
rect 53941 36805 53975 36839
rect 1593 36737 1627 36771
rect 18521 36737 18555 36771
rect 18705 36737 18739 36771
rect 18889 36737 18923 36771
rect 19533 36737 19567 36771
rect 20361 36737 20395 36771
rect 21005 36737 21039 36771
rect 24041 36737 24075 36771
rect 53665 36737 53699 36771
rect 53849 36737 53883 36771
rect 54038 36737 54072 36771
rect 21097 36669 21131 36703
rect 23857 36669 23891 36703
rect 19073 36601 19107 36635
rect 1777 36533 1811 36567
rect 21005 36533 21039 36567
rect 21373 36533 21407 36567
rect 23765 36533 23799 36567
rect 24225 36533 24259 36567
rect 54217 36533 54251 36567
rect 1777 36329 1811 36363
rect 23857 36329 23891 36363
rect 3065 36261 3099 36295
rect 20269 36193 20303 36227
rect 20729 36193 20763 36227
rect 2513 36125 2547 36159
rect 2886 36125 2920 36159
rect 20177 36125 20211 36159
rect 20453 36125 20487 36159
rect 22293 36125 22327 36159
rect 22569 36125 22603 36159
rect 22661 36125 22695 36159
rect 23305 36125 23339 36159
rect 23673 36125 23707 36159
rect 24593 36125 24627 36159
rect 24777 36125 24811 36159
rect 1685 36057 1719 36091
rect 2697 36057 2731 36091
rect 2789 36057 2823 36091
rect 22477 36057 22511 36091
rect 23489 36057 23523 36091
rect 23581 36057 23615 36091
rect 25145 36057 25179 36091
rect 57989 36057 58023 36091
rect 58357 36057 58391 36091
rect 22845 35989 22879 36023
rect 1777 35785 1811 35819
rect 19809 35785 19843 35819
rect 19533 35717 19567 35751
rect 40417 35717 40451 35751
rect 1685 35649 1719 35683
rect 19257 35649 19291 35683
rect 19441 35649 19475 35683
rect 19625 35649 19659 35683
rect 22661 35649 22695 35683
rect 40233 35649 40267 35683
rect 40509 35649 40543 35683
rect 40601 35649 40635 35683
rect 23397 35581 23431 35615
rect 40785 35513 40819 35547
rect 18889 35445 18923 35479
rect 22753 35241 22787 35275
rect 1869 35173 1903 35207
rect 22661 35105 22695 35139
rect 22753 35037 22787 35071
rect 40049 35037 40083 35071
rect 40325 35037 40359 35071
rect 40417 35037 40451 35071
rect 57897 35037 57931 35071
rect 1685 34969 1719 35003
rect 22477 34969 22511 35003
rect 40233 34969 40267 35003
rect 58173 34969 58207 35003
rect 22937 34901 22971 34935
rect 40601 34901 40635 34935
rect 58265 34697 58299 34731
rect 58081 34561 58115 34595
rect 1685 33949 1719 33983
rect 21281 33949 21315 33983
rect 21429 33949 21463 33983
rect 21557 33949 21591 33983
rect 21787 33949 21821 33983
rect 22477 33949 22511 33983
rect 22937 33949 22971 33983
rect 24593 33949 24627 33983
rect 24741 33949 24775 33983
rect 24869 33949 24903 33983
rect 25058 33949 25092 33983
rect 1869 33881 1903 33915
rect 21649 33881 21683 33915
rect 23213 33881 23247 33915
rect 24961 33881 24995 33915
rect 21925 33813 21959 33847
rect 25237 33813 25271 33847
rect 1869 33541 1903 33575
rect 21189 33541 21223 33575
rect 22385 33541 22419 33575
rect 36001 33541 36035 33575
rect 36093 33541 36127 33575
rect 1685 33473 1719 33507
rect 20913 33473 20947 33507
rect 21097 33473 21131 33507
rect 21281 33473 21315 33507
rect 22017 33473 22051 33507
rect 22165 33473 22199 33507
rect 22293 33473 22327 33507
rect 22523 33473 22557 33507
rect 35725 33473 35759 33507
rect 35873 33473 35907 33507
rect 36231 33473 36265 33507
rect 21465 33337 21499 33371
rect 22661 33269 22695 33303
rect 36369 33269 36403 33303
rect 21833 32997 21867 33031
rect 58173 32929 58207 32963
rect 21741 32861 21775 32895
rect 22017 32861 22051 32895
rect 57897 32861 57931 32895
rect 1685 32793 1719 32827
rect 22477 32793 22511 32827
rect 57069 32793 57103 32827
rect 1777 32725 1811 32759
rect 57161 32725 57195 32759
rect 1685 32385 1719 32419
rect 24869 32385 24903 32419
rect 24961 32385 24995 32419
rect 25145 32385 25179 32419
rect 25329 32317 25363 32351
rect 1777 32181 1811 32215
rect 22753 31841 22787 31875
rect 23029 31773 23063 31807
rect 23213 31773 23247 31807
rect 23305 31773 23339 31807
rect 23397 31773 23431 31807
rect 57897 31773 57931 31807
rect 58173 31773 58207 31807
rect 23581 31637 23615 31671
rect 24869 31433 24903 31467
rect 1685 31297 1719 31331
rect 24225 31297 24259 31331
rect 24373 31297 24407 31331
rect 24501 31297 24535 31331
rect 24593 31297 24627 31331
rect 24690 31297 24724 31331
rect 58081 31297 58115 31331
rect 1777 31093 1811 31127
rect 58265 31093 58299 31127
rect 19533 30821 19567 30855
rect 19441 30685 19475 30719
rect 19717 30685 19751 30719
rect 22845 30685 22879 30719
rect 23121 30685 23155 30719
rect 23213 30685 23247 30719
rect 1685 30617 1719 30651
rect 23029 30617 23063 30651
rect 1777 30549 1811 30583
rect 19901 30549 19935 30583
rect 23397 30549 23431 30583
rect 19441 30345 19475 30379
rect 19165 30277 19199 30311
rect 22293 30277 22327 30311
rect 1593 30209 1627 30243
rect 18797 30209 18831 30243
rect 18945 30209 18979 30243
rect 19073 30209 19107 30243
rect 19262 30209 19296 30243
rect 22017 30209 22051 30243
rect 22201 30209 22235 30243
rect 22385 30209 22419 30243
rect 23397 30209 23431 30243
rect 23489 30209 23523 30243
rect 23673 30209 23707 30243
rect 23857 30209 23891 30243
rect 1777 30141 1811 30175
rect 22569 30005 22603 30039
rect 23121 30005 23155 30039
rect 23581 30005 23615 30039
rect 58173 29665 58207 29699
rect 1593 29597 1627 29631
rect 22569 29597 22603 29631
rect 22661 29597 22695 29631
rect 22845 29597 22879 29631
rect 57897 29597 57931 29631
rect 1869 29529 1903 29563
rect 57069 29529 57103 29563
rect 23029 29461 23063 29495
rect 57161 29461 57195 29495
rect 9781 29257 9815 29291
rect 9413 29121 9447 29155
rect 9567 29121 9601 29155
rect 1777 28577 1811 28611
rect 1593 28509 1627 28543
rect 2513 28509 2547 28543
rect 2606 28509 2640 28543
rect 57897 28509 57931 28543
rect 2881 28441 2915 28475
rect 58173 28441 58207 28475
rect 1593 28033 1627 28067
rect 1777 27965 1811 27999
rect 1593 27421 1627 27455
rect 57989 27421 58023 27455
rect 1869 27353 1903 27387
rect 58081 27285 58115 27319
rect 2881 27081 2915 27115
rect 24317 27013 24351 27047
rect 1593 26945 1627 26979
rect 2513 26945 2547 26979
rect 2606 26945 2640 26979
rect 22753 26945 22787 26979
rect 23029 26945 23063 26979
rect 23949 26945 23983 26979
rect 24097 26945 24131 26979
rect 24225 26945 24259 26979
rect 24414 26945 24448 26979
rect 1777 26877 1811 26911
rect 23213 26877 23247 26911
rect 22845 26809 22879 26843
rect 24593 26809 24627 26843
rect 23673 26537 23707 26571
rect 58173 26401 58207 26435
rect 23121 26333 23155 26367
rect 23397 26333 23431 26367
rect 23489 26333 23523 26367
rect 57897 26333 57931 26367
rect 23305 26265 23339 26299
rect 1593 25857 1627 25891
rect 10701 25857 10735 25891
rect 10855 25857 10889 25891
rect 58081 25857 58115 25891
rect 1777 25789 1811 25823
rect 10885 25653 10919 25687
rect 58265 25653 58299 25687
rect 2881 25313 2915 25347
rect 1593 25245 1627 25279
rect 2513 25245 2547 25279
rect 2667 25245 2701 25279
rect 57897 25245 57931 25279
rect 1869 25177 1903 25211
rect 58173 25177 58207 25211
rect 1593 24769 1627 24803
rect 58081 24769 58115 24803
rect 1777 24701 1811 24735
rect 58265 24565 58299 24599
rect 2881 24361 2915 24395
rect 1593 24157 1627 24191
rect 2697 24157 2731 24191
rect 2851 24157 2885 24191
rect 1869 24089 1903 24123
rect 12265 23681 12299 23715
rect 12817 23613 12851 23647
rect 12173 23273 12207 23307
rect 1777 23137 1811 23171
rect 11253 23137 11287 23171
rect 58173 23137 58207 23171
rect 1593 23069 1627 23103
rect 10885 23069 10919 23103
rect 11039 23069 11073 23103
rect 11989 23069 12023 23103
rect 12143 23069 12177 23103
rect 57897 23069 57931 23103
rect 58173 22661 58207 22695
rect 1593 22593 1627 22627
rect 17233 22593 17267 22627
rect 17417 22593 17451 22627
rect 1777 22525 1811 22559
rect 17233 22389 17267 22423
rect 58265 22389 58299 22423
rect 17233 22117 17267 22151
rect 17969 22117 18003 22151
rect 9781 22049 9815 22083
rect 1593 21981 1627 22015
rect 9413 21981 9447 22015
rect 9567 21981 9601 22015
rect 17049 21981 17083 22015
rect 17785 21981 17819 22015
rect 18521 21981 18555 22015
rect 57897 21981 57931 22015
rect 1869 21913 1903 21947
rect 58173 21913 58207 21947
rect 18705 21845 18739 21879
rect 11069 21641 11103 21675
rect 18521 21641 18555 21675
rect 19257 21641 19291 21675
rect 23765 21641 23799 21675
rect 28825 21641 28859 21675
rect 1685 21505 1719 21539
rect 10701 21505 10735 21539
rect 10855 21505 10889 21539
rect 16037 21505 16071 21539
rect 17049 21505 17083 21539
rect 18337 21505 18371 21539
rect 18613 21505 18647 21539
rect 19073 21505 19107 21539
rect 19809 21505 19843 21539
rect 19993 21505 20027 21539
rect 20729 21505 20763 21539
rect 22845 21505 22879 21539
rect 23581 21505 23615 21539
rect 24317 21505 24351 21539
rect 25973 21505 26007 21539
rect 28641 21505 28675 21539
rect 38761 21505 38795 21539
rect 38853 21505 38887 21539
rect 42809 21505 42843 21539
rect 58081 21505 58115 21539
rect 16957 21437 16991 21471
rect 17417 21437 17451 21471
rect 38945 21437 38979 21471
rect 42625 21437 42659 21471
rect 18337 21369 18371 21403
rect 23029 21369 23063 21403
rect 24501 21369 24535 21403
rect 1777 21301 1811 21335
rect 16221 21301 16255 21335
rect 19809 21301 19843 21335
rect 20913 21301 20947 21335
rect 26157 21301 26191 21335
rect 38393 21301 38427 21335
rect 42993 21301 43027 21335
rect 58265 21301 58299 21335
rect 18429 21097 18463 21131
rect 19625 21097 19659 21131
rect 21097 21097 21131 21131
rect 26065 21097 26099 21131
rect 34989 21097 35023 21131
rect 12265 21029 12299 21063
rect 16773 21029 16807 21063
rect 20361 21029 20395 21063
rect 23949 21029 23983 21063
rect 27445 21029 27479 21063
rect 31585 21029 31619 21063
rect 53389 21029 53423 21063
rect 26433 20961 26467 20995
rect 27997 20961 28031 20995
rect 36369 20961 36403 20995
rect 42257 20961 42291 20995
rect 12081 20893 12115 20927
rect 12817 20893 12851 20927
rect 14289 20893 14323 20927
rect 15209 20893 15243 20927
rect 15393 20893 15427 20927
rect 15853 20893 15887 20927
rect 16589 20893 16623 20927
rect 17325 20893 17359 20927
rect 18153 20893 18187 20927
rect 18245 20893 18279 20927
rect 19441 20893 19475 20927
rect 20177 20893 20211 20927
rect 20913 20893 20947 20927
rect 21649 20893 21683 20927
rect 23765 20893 23799 20927
rect 24593 20893 24627 20927
rect 24777 20893 24811 20927
rect 25881 20893 25915 20927
rect 26617 20893 26651 20927
rect 27813 20893 27847 20927
rect 30665 20893 30699 20927
rect 30757 20893 30791 20927
rect 30941 20893 30975 20927
rect 31401 20893 31435 20927
rect 34805 20893 34839 20927
rect 35449 20893 35483 20927
rect 36921 20893 36955 20927
rect 38485 20893 38519 20927
rect 38577 20893 38611 20927
rect 42165 20893 42199 20927
rect 47501 20893 47535 20927
rect 47869 20893 47903 20927
rect 52837 20893 52871 20927
rect 53205 20893 53239 20927
rect 53941 20893 53975 20927
rect 54033 20893 54067 20927
rect 55873 20893 55907 20927
rect 56057 20893 56091 20927
rect 57897 20893 57931 20927
rect 43361 20825 43395 20859
rect 47685 20825 47719 20859
rect 47777 20825 47811 20859
rect 53021 20825 53055 20859
rect 53113 20825 53147 20859
rect 58173 20825 58207 20859
rect 13001 20757 13035 20791
rect 14473 20757 14507 20791
rect 15301 20757 15335 20791
rect 16037 20757 16071 20791
rect 17509 20757 17543 20791
rect 21833 20757 21867 20791
rect 24961 20757 24995 20791
rect 26801 20757 26835 20791
rect 27169 20757 27203 20791
rect 27905 20757 27939 20791
rect 35725 20757 35759 20791
rect 36093 20757 36127 20791
rect 36185 20757 36219 20791
rect 37105 20757 37139 20791
rect 38761 20757 38795 20791
rect 41705 20757 41739 20791
rect 42073 20757 42107 20791
rect 43637 20757 43671 20791
rect 48053 20757 48087 20791
rect 52561 20757 52595 20791
rect 54217 20757 54251 20791
rect 56241 20757 56275 20791
rect 16221 20553 16255 20587
rect 19181 20553 19215 20587
rect 19349 20553 19383 20587
rect 22477 20553 22511 20587
rect 25605 20553 25639 20587
rect 28549 20553 28583 20587
rect 30113 20553 30147 20587
rect 30665 20553 30699 20587
rect 31033 20553 31067 20587
rect 40049 20553 40083 20587
rect 49617 20553 49651 20587
rect 56333 20553 56367 20587
rect 18521 20485 18555 20519
rect 18981 20485 19015 20519
rect 19809 20485 19843 20519
rect 20025 20485 20059 20519
rect 24032 20485 24066 20519
rect 25973 20485 26007 20519
rect 27414 20485 27448 20519
rect 34805 20485 34839 20519
rect 35510 20485 35544 20519
rect 37841 20485 37875 20519
rect 42901 20485 42935 20519
rect 43131 20485 43165 20519
rect 44215 20485 44249 20519
rect 1593 20417 1627 20451
rect 8033 20417 8067 20451
rect 10241 20417 10275 20451
rect 11989 20417 12023 20451
rect 13185 20417 13219 20451
rect 13277 20417 13311 20451
rect 14013 20417 14047 20451
rect 15301 20417 15335 20451
rect 16037 20417 16071 20451
rect 16865 20417 16899 20451
rect 17141 20417 17175 20451
rect 21189 20417 21223 20451
rect 22385 20417 22419 20451
rect 26065 20417 26099 20451
rect 29193 20417 29227 20451
rect 29929 20417 29963 20451
rect 33241 20417 33275 20451
rect 33425 20417 33459 20451
rect 33609 20417 33643 20451
rect 34621 20417 34655 20451
rect 37657 20417 37691 20451
rect 38761 20417 38795 20451
rect 41613 20417 41647 20451
rect 42809 20417 42843 20451
rect 42993 20417 43027 20451
rect 43729 20417 43763 20451
rect 43913 20417 43947 20451
rect 44005 20417 44039 20451
rect 44097 20417 44131 20451
rect 44373 20417 44407 20451
rect 46029 20417 46063 20451
rect 48504 20417 48538 20451
rect 50445 20417 50479 20451
rect 51641 20417 51675 20451
rect 53113 20417 53147 20451
rect 53380 20417 53414 20451
rect 55209 20417 55243 20451
rect 1777 20349 1811 20383
rect 12817 20349 12851 20383
rect 13001 20349 13035 20383
rect 13093 20349 13127 20383
rect 21005 20349 21039 20383
rect 22661 20349 22695 20383
rect 23765 20349 23799 20383
rect 26157 20349 26191 20383
rect 27169 20349 27203 20383
rect 31125 20349 31159 20383
rect 31217 20349 31251 20383
rect 34437 20349 34471 20383
rect 35265 20349 35299 20383
rect 37473 20349 37507 20383
rect 38485 20349 38519 20383
rect 41429 20349 41463 20383
rect 43269 20349 43303 20383
rect 48237 20349 48271 20383
rect 50261 20349 50295 20383
rect 51457 20349 51491 20383
rect 54953 20349 54987 20383
rect 22017 20281 22051 20315
rect 54493 20281 54527 20315
rect 8217 20213 8251 20247
rect 10425 20213 10459 20247
rect 12173 20213 12207 20247
rect 14197 20213 14231 20247
rect 15485 20213 15519 20247
rect 19165 20213 19199 20247
rect 19993 20213 20027 20247
rect 20177 20213 20211 20247
rect 21373 20213 21407 20247
rect 25145 20213 25179 20247
rect 29377 20213 29411 20247
rect 36645 20213 36679 20247
rect 41797 20213 41831 20247
rect 42625 20213 42659 20247
rect 46305 20213 46339 20247
rect 50629 20213 50663 20247
rect 51825 20213 51859 20247
rect 9321 20009 9355 20043
rect 18337 20009 18371 20043
rect 20177 20009 20211 20043
rect 32045 20009 32079 20043
rect 40877 20009 40911 20043
rect 44649 20009 44683 20043
rect 47593 20009 47627 20043
rect 48513 20009 48547 20043
rect 51825 20009 51859 20043
rect 53757 20009 53791 20043
rect 56057 20009 56091 20043
rect 8125 19941 8159 19975
rect 11897 19941 11931 19975
rect 13737 19941 13771 19975
rect 16405 19941 16439 19975
rect 19625 19941 19659 19975
rect 24593 19941 24627 19975
rect 42717 19941 42751 19975
rect 8217 19873 8251 19907
rect 11621 19873 11655 19907
rect 16957 19873 16991 19907
rect 20729 19873 20763 19907
rect 24041 19873 24075 19907
rect 25237 19873 25271 19907
rect 26801 19873 26835 19907
rect 28273 19873 28307 19907
rect 32873 19873 32907 19907
rect 38393 19873 38427 19907
rect 46213 19873 46247 19907
rect 48145 19873 48179 19907
rect 50445 19873 50479 19907
rect 52377 19873 52411 19907
rect 1593 19805 1627 19839
rect 7021 19805 7055 19839
rect 9137 19805 9171 19839
rect 9873 19805 9907 19839
rect 10609 19805 10643 19839
rect 11529 19805 11563 19839
rect 12357 19805 12391 19839
rect 14289 19805 14323 19839
rect 15025 19805 15059 19839
rect 17224 19805 17258 19839
rect 19993 19805 20027 19839
rect 20996 19805 21030 19839
rect 23305 19805 23339 19839
rect 23397 19805 23431 19839
rect 23581 19805 23615 19839
rect 25789 19805 25823 19839
rect 25973 19805 26007 19839
rect 26985 19805 27019 19839
rect 28089 19805 28123 19839
rect 30665 19805 30699 19839
rect 33140 19805 33174 19839
rect 35817 19805 35851 19839
rect 38117 19805 38151 19839
rect 41337 19805 41371 19839
rect 43269 19805 43303 19839
rect 45385 19805 45419 19839
rect 45569 19805 45603 19839
rect 48329 19805 48363 19839
rect 52633 19805 52667 19839
rect 54309 19805 54343 19839
rect 54585 19805 54619 19839
rect 54677 19805 54711 19839
rect 55505 19805 55539 19839
rect 55873 19805 55907 19839
rect 56885 19805 56919 19839
rect 57141 19805 57175 19839
rect 1869 19737 1903 19771
rect 7757 19737 7791 19771
rect 12602 19737 12636 19771
rect 15292 19737 15326 19771
rect 19809 19737 19843 19771
rect 24961 19737 24995 19771
rect 25053 19737 25087 19771
rect 30932 19737 30966 19771
rect 36084 19737 36118 19771
rect 40509 19737 40543 19771
rect 40693 19737 40727 19771
rect 41604 19737 41638 19771
rect 43514 19737 43548 19771
rect 45753 19737 45787 19771
rect 46458 19737 46492 19771
rect 50690 19737 50724 19771
rect 54493 19737 54527 19771
rect 55689 19737 55723 19771
rect 55781 19737 55815 19771
rect 7205 19669 7239 19703
rect 10057 19669 10091 19703
rect 10793 19669 10827 19703
rect 14473 19669 14507 19703
rect 19901 19669 19935 19703
rect 22109 19669 22143 19703
rect 26157 19669 26191 19703
rect 27169 19669 27203 19703
rect 27629 19669 27663 19703
rect 27997 19669 28031 19703
rect 34253 19669 34287 19703
rect 37197 19669 37231 19703
rect 37749 19669 37783 19703
rect 38209 19669 38243 19703
rect 54861 19669 54895 19703
rect 58265 19669 58299 19703
rect 8217 19465 8251 19499
rect 10149 19465 10183 19499
rect 11161 19465 11195 19499
rect 13829 19465 13863 19499
rect 15761 19465 15795 19499
rect 19073 19465 19107 19499
rect 24777 19465 24811 19499
rect 31677 19465 31711 19499
rect 33609 19465 33643 19499
rect 33977 19465 34011 19499
rect 34069 19465 34103 19499
rect 35909 19465 35943 19499
rect 44281 19465 44315 19499
rect 46857 19465 46891 19499
rect 51641 19465 51675 19499
rect 54953 19465 54987 19499
rect 1869 19397 1903 19431
rect 10701 19397 10735 19431
rect 27690 19397 27724 19431
rect 36277 19397 36311 19431
rect 42073 19397 42107 19431
rect 43146 19397 43180 19431
rect 48053 19397 48087 19431
rect 51273 19397 51307 19431
rect 51365 19397 51399 19431
rect 1593 19329 1627 19363
rect 7104 19329 7138 19363
rect 8769 19329 8803 19363
rect 9036 19329 9070 19363
rect 11713 19329 11747 19363
rect 12449 19329 12483 19363
rect 12716 19329 12750 19363
rect 14381 19329 14415 19363
rect 14648 19329 14682 19363
rect 17305 19329 17339 19363
rect 19165 19329 19199 19363
rect 19257 19329 19291 19363
rect 20085 19329 20119 19363
rect 20352 19329 20386 19363
rect 22017 19329 22051 19363
rect 23397 19329 23431 19363
rect 23664 19329 23698 19363
rect 25605 19329 25639 19363
rect 26341 19329 26375 19363
rect 27445 19329 27479 19363
rect 30297 19329 30331 19363
rect 30564 19329 30598 19363
rect 36369 19329 36403 19363
rect 41705 19329 41739 19363
rect 41889 19329 41923 19363
rect 42901 19329 42935 19363
rect 45477 19329 45511 19363
rect 45744 19329 45778 19363
rect 47777 19329 47811 19363
rect 49801 19329 49835 19363
rect 49985 19329 50019 19363
rect 50077 19329 50111 19363
rect 50193 19329 50227 19363
rect 51089 19329 51123 19363
rect 51457 19329 51491 19363
rect 54769 19329 54803 19363
rect 6837 19261 6871 19295
rect 17049 19261 17083 19295
rect 19441 19261 19475 19295
rect 34253 19261 34287 19295
rect 36553 19261 36587 19295
rect 54585 19261 54619 19295
rect 10977 19193 11011 19227
rect 18889 19193 18923 19227
rect 26525 19193 26559 19227
rect 11897 19125 11931 19159
rect 18429 19125 18463 19159
rect 21465 19125 21499 19159
rect 22201 19125 22235 19159
rect 25789 19125 25823 19159
rect 28825 19125 28859 19159
rect 50353 19125 50387 19159
rect 8033 18921 8067 18955
rect 10609 18921 10643 18955
rect 11529 18921 11563 18955
rect 13461 18921 13495 18955
rect 16589 18921 16623 18955
rect 18797 18921 18831 18955
rect 21005 18921 21039 18955
rect 22385 18921 22419 18955
rect 30481 18921 30515 18955
rect 36737 18921 36771 18955
rect 44005 18921 44039 18955
rect 45661 18921 45695 18955
rect 46673 18921 46707 18955
rect 7481 18853 7515 18887
rect 9137 18853 9171 18887
rect 15853 18853 15887 18887
rect 18061 18853 18095 18887
rect 24685 18853 24719 18887
rect 25973 18853 26007 18887
rect 28917 18853 28951 18887
rect 6101 18785 6135 18819
rect 9689 18785 9723 18819
rect 10241 18785 10275 18819
rect 12081 18785 12115 18819
rect 14565 18785 14599 18819
rect 14841 18785 14875 18819
rect 19441 18785 19475 18819
rect 21649 18785 21683 18819
rect 26525 18785 26559 18819
rect 31401 18785 31435 18819
rect 31493 18785 31527 18819
rect 37381 18785 37415 18819
rect 38761 18785 38795 18819
rect 41245 18785 41279 18819
rect 55505 18785 55539 18819
rect 1593 18717 1627 18751
rect 5365 18717 5399 18751
rect 8217 18717 8251 18751
rect 8309 18717 8343 18751
rect 8401 18717 8435 18751
rect 8493 18717 8527 18751
rect 10333 18717 10367 18751
rect 11437 18717 11471 18751
rect 11621 18717 11655 18751
rect 14473 18717 14507 18751
rect 15669 18717 15703 18751
rect 16405 18717 16439 18751
rect 17141 18717 17175 18751
rect 17877 18717 17911 18751
rect 18613 18717 18647 18751
rect 19625 18717 19659 18751
rect 19901 18717 19935 18751
rect 20085 18717 20119 18751
rect 21373 18717 21407 18751
rect 22201 18717 22235 18751
rect 22937 18717 22971 18751
rect 23765 18717 23799 18751
rect 25789 18717 25823 18751
rect 28365 18717 28399 18751
rect 28641 18717 28675 18751
rect 28785 18717 28819 18751
rect 30205 18717 30239 18751
rect 30297 18717 30331 18751
rect 31309 18717 31343 18751
rect 32413 18717 32447 18751
rect 37105 18717 37139 18751
rect 38945 18717 38979 18751
rect 40969 18717 41003 18751
rect 42533 18717 42567 18751
rect 42626 18717 42660 18751
rect 42998 18717 43032 18751
rect 45385 18717 45419 18751
rect 45477 18717 45511 18751
rect 46121 18717 46155 18751
rect 46489 18717 46523 18751
rect 47225 18717 47259 18751
rect 48513 18717 48547 18751
rect 48697 18717 48731 18751
rect 55689 18717 55723 18751
rect 56977 18717 57011 18751
rect 57989 18717 58023 18751
rect 1869 18649 1903 18683
rect 6368 18649 6402 18683
rect 9413 18649 9447 18683
rect 12326 18649 12360 18683
rect 24961 18649 24995 18683
rect 25237 18649 25271 18683
rect 26792 18649 26826 18683
rect 28549 18649 28583 18683
rect 42809 18649 42843 18683
rect 42901 18649 42935 18683
rect 43637 18649 43671 18683
rect 43821 18649 43855 18683
rect 46305 18649 46339 18683
rect 46397 18649 46431 18683
rect 57253 18649 57287 18683
rect 5549 18581 5583 18615
rect 9321 18581 9355 18615
rect 9505 18581 9539 18615
rect 17325 18581 17359 18615
rect 21465 18581 21499 18615
rect 23121 18581 23155 18615
rect 23949 18581 23983 18615
rect 25145 18581 25179 18615
rect 27905 18581 27939 18615
rect 30941 18581 30975 18615
rect 32597 18581 32631 18615
rect 37197 18581 37231 18615
rect 39129 18581 39163 18615
rect 40601 18581 40635 18615
rect 41061 18581 41095 18615
rect 43177 18581 43211 18615
rect 47501 18581 47535 18615
rect 48881 18581 48915 18615
rect 55873 18581 55907 18615
rect 58081 18581 58115 18615
rect 10517 18377 10551 18411
rect 12173 18377 12207 18411
rect 14657 18377 14691 18411
rect 16221 18377 16255 18411
rect 18521 18377 18555 18411
rect 26525 18377 26559 18411
rect 27261 18377 27295 18411
rect 27629 18377 27663 18411
rect 46489 18377 46523 18411
rect 50077 18377 50111 18411
rect 55137 18377 55171 18411
rect 57253 18377 57287 18411
rect 13093 18309 13127 18343
rect 30849 18309 30883 18343
rect 30941 18309 30975 18343
rect 34345 18309 34379 18343
rect 42809 18309 42843 18343
rect 42901 18309 42935 18343
rect 46121 18309 46155 18343
rect 46213 18309 46247 18343
rect 54861 18309 54895 18343
rect 56140 18309 56174 18343
rect 5733 18241 5767 18275
rect 6745 18241 6779 18275
rect 8217 18241 8251 18275
rect 10333 18241 10367 18275
rect 11989 18241 12023 18275
rect 12909 18241 12943 18275
rect 13001 18241 13035 18275
rect 13277 18241 13311 18275
rect 14473 18241 14507 18275
rect 15301 18241 15335 18275
rect 16037 18241 16071 18275
rect 17141 18241 17175 18275
rect 17408 18241 17442 18275
rect 19533 18241 19567 18275
rect 20453 18241 20487 18275
rect 21189 18241 21223 18275
rect 22017 18241 22051 18275
rect 23121 18241 23155 18275
rect 23305 18241 23339 18275
rect 24317 18241 24351 18275
rect 26341 18241 26375 18275
rect 29469 18241 29503 18275
rect 29561 18241 29595 18275
rect 29745 18241 29779 18275
rect 29837 18241 29871 18275
rect 39129 18241 39163 18275
rect 42625 18241 42659 18275
rect 42993 18241 43027 18275
rect 45937 18241 45971 18275
rect 46305 18241 46339 18275
rect 48964 18241 48998 18275
rect 54585 18241 54619 18275
rect 54769 18241 54803 18275
rect 54953 18241 54987 18275
rect 6837 18173 6871 18207
rect 7113 18173 7147 18207
rect 8493 18173 8527 18207
rect 19349 18173 19383 18207
rect 27721 18173 27755 18207
rect 27905 18173 27939 18207
rect 30757 18173 30791 18207
rect 32321 18173 32355 18207
rect 32505 18173 32539 18207
rect 32597 18173 32631 18207
rect 32689 18173 32723 18207
rect 32781 18173 32815 18207
rect 34437 18173 34471 18207
rect 34621 18173 34655 18207
rect 38853 18173 38887 18207
rect 40233 18173 40267 18207
rect 48697 18173 48731 18207
rect 55873 18173 55907 18207
rect 9781 18105 9815 18139
rect 12725 18105 12759 18139
rect 22201 18105 22235 18139
rect 23489 18105 23523 18139
rect 24501 18105 24535 18139
rect 30389 18105 30423 18139
rect 43177 18105 43211 18139
rect 5917 18037 5951 18071
rect 15485 18037 15519 18071
rect 19717 18037 19751 18071
rect 20637 18037 20671 18071
rect 21373 18037 21407 18071
rect 29285 18037 29319 18071
rect 33977 18037 34011 18071
rect 9965 17833 9999 17867
rect 14473 17833 14507 17867
rect 15301 17833 15335 17867
rect 16773 17833 16807 17867
rect 18613 17833 18647 17867
rect 32045 17833 32079 17867
rect 53021 17833 53055 17867
rect 58265 17833 58299 17867
rect 29837 17765 29871 17799
rect 38761 17765 38795 17799
rect 41613 17765 41647 17799
rect 48513 17765 48547 17799
rect 1777 17697 1811 17731
rect 8125 17697 8159 17731
rect 8585 17697 8619 17731
rect 19533 17697 19567 17731
rect 25605 17697 25639 17731
rect 31677 17697 31711 17731
rect 32505 17697 32539 17731
rect 34069 17697 34103 17731
rect 35081 17697 35115 17731
rect 39405 17697 39439 17731
rect 40233 17697 40267 17731
rect 55689 17697 55723 17731
rect 56885 17697 56919 17731
rect 1593 17629 1627 17663
rect 6561 17629 6595 17663
rect 8217 17629 8251 17663
rect 9137 17629 9171 17663
rect 9873 17629 9907 17663
rect 10057 17629 10091 17663
rect 14289 17629 14323 17663
rect 15117 17629 15151 17663
rect 15853 17629 15887 17663
rect 16589 17629 16623 17663
rect 17693 17629 17727 17663
rect 18429 17629 18463 17663
rect 19441 17629 19475 17663
rect 19625 17629 19659 17663
rect 20085 17629 20119 17663
rect 20913 17629 20947 17663
rect 21005 17629 21039 17663
rect 24777 17629 24811 17663
rect 25145 17629 25179 17663
rect 25789 17629 25823 17663
rect 27077 17629 27111 17663
rect 27353 17629 27387 17663
rect 27445 17629 27479 17663
rect 28181 17629 28215 17663
rect 28329 17629 28363 17663
rect 28549 17629 28583 17663
rect 28646 17629 28680 17663
rect 29745 17629 29779 17663
rect 30021 17629 30055 17663
rect 31861 17629 31895 17663
rect 32689 17629 32723 17663
rect 33793 17629 33827 17663
rect 34897 17629 34931 17663
rect 40500 17629 40534 17663
rect 47961 17629 47995 17663
rect 48329 17629 48363 17663
rect 50629 17629 50663 17663
rect 50997 17629 51031 17663
rect 51641 17629 51675 17663
rect 55505 17629 55539 17663
rect 27261 17561 27295 17595
rect 28457 17561 28491 17595
rect 39129 17561 39163 17595
rect 39221 17561 39255 17595
rect 48145 17561 48179 17595
rect 48237 17561 48271 17595
rect 50813 17561 50847 17595
rect 50905 17561 50939 17595
rect 51908 17561 51942 17595
rect 57130 17561 57164 17595
rect 6745 17493 6779 17527
rect 9321 17493 9355 17527
rect 16037 17493 16071 17527
rect 17877 17493 17911 17527
rect 20269 17493 20303 17527
rect 21189 17493 21223 17527
rect 24685 17493 24719 17527
rect 24869 17493 24903 17527
rect 24961 17493 24995 17527
rect 25973 17493 26007 17527
rect 27629 17493 27663 17527
rect 28825 17493 28859 17527
rect 30205 17493 30239 17527
rect 32873 17493 32907 17527
rect 33425 17493 33459 17527
rect 33885 17493 33919 17527
rect 51181 17493 51215 17527
rect 8769 17289 8803 17323
rect 15393 17289 15427 17323
rect 17233 17289 17267 17323
rect 17969 17289 18003 17323
rect 18797 17289 18831 17323
rect 20729 17289 20763 17323
rect 24961 17289 24995 17323
rect 25237 17289 25271 17323
rect 38301 17289 38335 17323
rect 51825 17289 51859 17323
rect 56333 17289 56367 17323
rect 25421 17221 25455 17255
rect 28089 17221 28123 17255
rect 28181 17221 28215 17255
rect 33876 17221 33910 17255
rect 38669 17221 38703 17255
rect 1593 17153 1627 17187
rect 8585 17153 8619 17187
rect 15301 17153 15335 17187
rect 15485 17153 15519 17187
rect 16037 17153 16071 17187
rect 17049 17153 17083 17187
rect 17785 17153 17819 17187
rect 18613 17153 18647 17187
rect 19349 17153 19383 17187
rect 19901 17153 19935 17187
rect 20085 17153 20119 17187
rect 21097 17153 21131 17187
rect 22017 17153 22051 17187
rect 25053 17153 25087 17187
rect 25165 17153 25199 17187
rect 27905 17153 27939 17187
rect 28325 17153 28359 17187
rect 32781 17153 32815 17187
rect 33609 17153 33643 17187
rect 40969 17153 41003 17187
rect 51457 17153 51491 17187
rect 51641 17153 51675 17187
rect 54125 17153 54159 17187
rect 54953 17153 54987 17187
rect 55137 17153 55171 17187
rect 55229 17153 55263 17187
rect 55321 17153 55355 17187
rect 56149 17153 56183 17187
rect 57069 17153 57103 17187
rect 1777 17085 1811 17119
rect 19993 17085 20027 17119
rect 20453 17085 20487 17119
rect 21189 17085 21223 17119
rect 21373 17085 21407 17119
rect 32505 17085 32539 17119
rect 32597 17085 32631 17119
rect 32689 17085 32723 17119
rect 38761 17085 38795 17119
rect 38945 17085 38979 17119
rect 41061 17085 41095 17119
rect 41245 17085 41279 17119
rect 53941 17085 53975 17119
rect 55965 17085 55999 17119
rect 57345 17085 57379 17119
rect 28457 17017 28491 17051
rect 55505 17017 55539 17051
rect 2421 16949 2455 16983
rect 16221 16949 16255 16983
rect 19533 16949 19567 16983
rect 22201 16949 22235 16983
rect 32321 16949 32355 16983
rect 34989 16949 35023 16983
rect 40601 16949 40635 16983
rect 54309 16949 54343 16983
rect 16221 16745 16255 16779
rect 22661 16745 22695 16779
rect 57161 16745 57195 16779
rect 18705 16677 18739 16711
rect 19625 16677 19659 16711
rect 13461 16609 13495 16643
rect 13645 16609 13679 16643
rect 20821 16609 20855 16643
rect 25973 16609 26007 16643
rect 27721 16609 27755 16643
rect 28457 16609 28491 16643
rect 28641 16609 28675 16643
rect 32505 16609 32539 16643
rect 32965 16609 32999 16643
rect 36737 16609 36771 16643
rect 36921 16609 36955 16643
rect 37473 16609 37507 16643
rect 41521 16609 41555 16643
rect 45201 16609 45235 16643
rect 51457 16609 51491 16643
rect 53573 16609 53607 16643
rect 1593 16541 1627 16575
rect 12265 16541 12299 16575
rect 13369 16541 13403 16575
rect 13553 16541 13587 16575
rect 16221 16541 16255 16575
rect 16405 16541 16439 16575
rect 16865 16541 16899 16575
rect 17132 16541 17166 16575
rect 18705 16541 18739 16575
rect 18889 16541 18923 16575
rect 19441 16541 19475 16575
rect 20177 16541 20211 16575
rect 20361 16541 20395 16575
rect 21088 16541 21122 16575
rect 22661 16541 22695 16575
rect 22845 16541 22879 16575
rect 33232 16541 33266 16575
rect 37740 16541 37774 16575
rect 40693 16541 40727 16575
rect 40858 16541 40892 16575
rect 40969 16541 41003 16575
rect 41061 16541 41095 16575
rect 41705 16541 41739 16575
rect 41797 16541 41831 16575
rect 41981 16541 42015 16575
rect 42073 16541 42107 16575
rect 51641 16541 51675 16575
rect 53840 16541 53874 16575
rect 57989 16541 58023 16575
rect 1869 16473 1903 16507
rect 20269 16473 20303 16507
rect 26240 16473 26274 16507
rect 32137 16473 32171 16507
rect 32321 16473 32355 16507
rect 36645 16473 36679 16507
rect 45468 16473 45502 16507
rect 52377 16473 52411 16507
rect 57069 16473 57103 16507
rect 12449 16405 12483 16439
rect 13185 16405 13219 16439
rect 18245 16405 18279 16439
rect 22201 16405 22235 16439
rect 27353 16405 27387 16439
rect 27997 16405 28031 16439
rect 28365 16405 28399 16439
rect 34345 16405 34379 16439
rect 36277 16405 36311 16439
rect 38853 16405 38887 16439
rect 40509 16405 40543 16439
rect 46581 16405 46615 16439
rect 51825 16405 51859 16439
rect 52469 16405 52503 16439
rect 54953 16405 54987 16439
rect 58081 16405 58115 16439
rect 13553 16201 13587 16235
rect 22201 16201 22235 16235
rect 24133 16201 24167 16235
rect 27169 16201 27203 16235
rect 27537 16201 27571 16235
rect 29469 16201 29503 16235
rect 43177 16201 43211 16235
rect 45477 16201 45511 16235
rect 46397 16201 46431 16235
rect 46857 16201 46891 16235
rect 51641 16201 51675 16235
rect 53021 16201 53055 16235
rect 54217 16201 54251 16235
rect 18889 16133 18923 16167
rect 19257 16133 19291 16167
rect 19441 16133 19475 16167
rect 29561 16133 29595 16167
rect 31217 16133 31251 16167
rect 37473 16133 37507 16167
rect 38485 16133 38519 16167
rect 42901 16133 42935 16167
rect 46765 16133 46799 16167
rect 51273 16133 51307 16167
rect 53941 16133 53975 16167
rect 1593 16065 1627 16099
rect 2329 16065 2363 16099
rect 9873 16065 9907 16099
rect 11713 16065 11747 16099
rect 12449 16065 12483 16099
rect 13737 16065 13771 16099
rect 13829 16065 13863 16099
rect 13921 16065 13955 16099
rect 15761 16065 15795 16099
rect 17049 16065 17083 16099
rect 17316 16065 17350 16099
rect 19073 16065 19107 16099
rect 19165 16065 19199 16099
rect 20361 16065 20395 16099
rect 21097 16065 21131 16099
rect 22017 16065 22051 16099
rect 23121 16065 23155 16099
rect 23305 16065 23339 16099
rect 23949 16065 23983 16099
rect 25053 16065 25087 16099
rect 26341 16065 26375 16099
rect 31677 16065 31711 16099
rect 32597 16065 32631 16099
rect 32689 16065 32723 16099
rect 32873 16065 32907 16099
rect 32965 16065 32999 16099
rect 37657 16065 37691 16099
rect 38669 16065 38703 16099
rect 41521 16065 41555 16099
rect 41889 16065 41923 16099
rect 42625 16065 42659 16099
rect 42809 16065 42843 16099
rect 42993 16065 43027 16099
rect 44189 16065 44223 16099
rect 48033 16065 48067 16099
rect 51089 16065 51123 16099
rect 51365 16065 51399 16099
rect 51457 16065 51491 16099
rect 52101 16065 52135 16099
rect 52929 16065 52963 16099
rect 53113 16065 53147 16099
rect 53665 16065 53699 16099
rect 53849 16065 53883 16099
rect 54033 16065 54067 16099
rect 1777 15997 1811 16031
rect 14013 15997 14047 16031
rect 25329 15997 25363 16031
rect 27629 15997 27663 16031
rect 27813 15997 27847 16031
rect 29745 15997 29779 16031
rect 41613 15997 41647 16031
rect 41981 15997 42015 16031
rect 46949 15997 46983 16031
rect 47777 15997 47811 16031
rect 11897 15929 11931 15963
rect 18429 15929 18463 15963
rect 21281 15929 21315 15963
rect 26525 15929 26559 15963
rect 40969 15929 41003 15963
rect 10057 15861 10091 15895
rect 12633 15861 12667 15895
rect 15945 15861 15979 15895
rect 20545 15861 20579 15895
rect 23489 15861 23523 15895
rect 29101 15861 29135 15895
rect 32413 15861 32447 15895
rect 37749 15861 37783 15895
rect 38761 15861 38795 15895
rect 49157 15861 49191 15895
rect 50721 15861 50755 15895
rect 52285 15861 52319 15895
rect 10333 15657 10367 15691
rect 13093 15657 13127 15691
rect 17785 15657 17819 15691
rect 21741 15657 21775 15691
rect 23305 15657 23339 15691
rect 41705 15657 41739 15691
rect 48145 15657 48179 15691
rect 12449 15589 12483 15623
rect 18705 15589 18739 15623
rect 20637 15589 20671 15623
rect 23949 15589 23983 15623
rect 52929 15589 52963 15623
rect 11069 15521 11103 15555
rect 13461 15521 13495 15555
rect 18797 15521 18831 15555
rect 19625 15521 19659 15555
rect 19901 15521 19935 15555
rect 35449 15521 35483 15555
rect 9965 15453 9999 15487
rect 10149 15453 10183 15487
rect 13277 15453 13311 15487
rect 13369 15453 13403 15487
rect 13553 15453 13587 15487
rect 14289 15453 14323 15487
rect 15301 15453 15335 15487
rect 16129 15453 16163 15487
rect 16865 15453 16899 15487
rect 17601 15453 17635 15487
rect 19717 15453 19751 15487
rect 19809 15453 19843 15487
rect 20453 15453 20487 15487
rect 21557 15453 21591 15487
rect 22753 15453 22787 15487
rect 23173 15453 23207 15487
rect 23857 15453 23891 15487
rect 24593 15453 24627 15487
rect 26525 15453 26559 15487
rect 26709 15453 26743 15487
rect 27537 15453 27571 15487
rect 35265 15453 35299 15487
rect 36553 15453 36587 15487
rect 36809 15453 36843 15487
rect 41061 15453 41095 15487
rect 41209 15453 41243 15487
rect 41337 15453 41371 15487
rect 41429 15453 41463 15487
rect 41567 15453 41601 15487
rect 51549 15453 51583 15487
rect 57897 15453 57931 15487
rect 11336 15385 11370 15419
rect 18337 15385 18371 15419
rect 22937 15385 22971 15419
rect 23029 15385 23063 15419
rect 24860 15385 24894 15419
rect 26893 15385 26927 15419
rect 27804 15385 27838 15419
rect 46857 15385 46891 15419
rect 51816 15385 51850 15419
rect 58173 15385 58207 15419
rect 14473 15317 14507 15351
rect 15485 15317 15519 15351
rect 16313 15317 16347 15351
rect 17049 15317 17083 15351
rect 19441 15317 19475 15351
rect 25973 15317 26007 15351
rect 28917 15317 28951 15351
rect 34897 15317 34931 15351
rect 35357 15317 35391 15351
rect 37933 15317 37967 15351
rect 19089 15113 19123 15147
rect 19257 15113 19291 15147
rect 19901 15113 19935 15147
rect 22845 15113 22879 15147
rect 25329 15113 25363 15147
rect 27905 15113 27939 15147
rect 29837 15113 29871 15147
rect 38669 15113 38703 15147
rect 41797 15113 41831 15147
rect 43085 15113 43119 15147
rect 47777 15113 47811 15147
rect 17969 15045 18003 15079
rect 18153 15045 18187 15079
rect 18889 15045 18923 15079
rect 24317 15045 24351 15079
rect 24409 15045 24443 15079
rect 25697 15045 25731 15079
rect 28724 15045 28758 15079
rect 30941 15045 30975 15079
rect 41429 15045 41463 15079
rect 1593 14977 1627 15011
rect 9413 14977 9447 15011
rect 11897 14977 11931 15011
rect 12725 14977 12759 15011
rect 13461 14977 13495 15011
rect 16037 14977 16071 15011
rect 16865 14977 16899 15011
rect 19717 14977 19751 15011
rect 22017 14977 22051 15011
rect 22109 14977 22143 15011
rect 22786 14977 22820 15011
rect 23213 14977 23247 15011
rect 24133 14977 24167 15011
rect 24506 14977 24540 15011
rect 25789 14977 25823 15011
rect 27721 14977 27755 15011
rect 30389 14977 30423 15011
rect 32321 14977 32355 15011
rect 34437 14977 34471 15011
rect 34704 14977 34738 15011
rect 38666 14977 38700 15011
rect 41245 14977 41279 15011
rect 41521 14977 41555 15011
rect 41613 14977 41647 15011
rect 42993 14977 43027 15011
rect 48145 14977 48179 15011
rect 1777 14909 1811 14943
rect 9689 14909 9723 14943
rect 11989 14909 12023 14943
rect 13737 14909 13771 14943
rect 18245 14909 18279 14943
rect 23305 14909 23339 14943
rect 25881 14909 25915 14943
rect 27537 14909 27571 14943
rect 28457 14909 28491 14943
rect 32597 14909 32631 14943
rect 39129 14909 39163 14943
rect 48237 14909 48271 14943
rect 48329 14909 48363 14943
rect 12265 14841 12299 14875
rect 17693 14841 17727 14875
rect 24685 14841 24719 14875
rect 10977 14773 11011 14807
rect 12909 14773 12943 14807
rect 15025 14773 15059 14807
rect 16221 14773 16255 14807
rect 17049 14773 17083 14807
rect 19073 14773 19107 14807
rect 22661 14773 22695 14807
rect 33885 14773 33919 14807
rect 35817 14773 35851 14807
rect 38485 14773 38519 14807
rect 39037 14773 39071 14807
rect 12817 14569 12851 14603
rect 19809 14569 19843 14603
rect 21833 14569 21867 14603
rect 26617 14569 26651 14603
rect 31769 14569 31803 14603
rect 39405 14569 39439 14603
rect 58081 14569 58115 14603
rect 22845 14501 22879 14535
rect 32505 14501 32539 14535
rect 9321 14433 9355 14467
rect 11437 14433 11471 14467
rect 14381 14433 14415 14467
rect 16773 14433 16807 14467
rect 18797 14433 18831 14467
rect 23305 14433 23339 14467
rect 23949 14433 23983 14467
rect 28825 14433 28859 14467
rect 29745 14433 29779 14467
rect 42993 14433 43027 14467
rect 43269 14433 43303 14467
rect 1593 14365 1627 14399
rect 8309 14365 8343 14399
rect 9597 14365 9631 14399
rect 13461 14365 13495 14399
rect 14657 14365 14691 14399
rect 17029 14365 17063 14399
rect 18705 14365 18739 14399
rect 18889 14365 18923 14399
rect 19441 14365 19475 14399
rect 19625 14365 19659 14399
rect 20269 14365 20303 14399
rect 21649 14365 21683 14399
rect 23029 14365 23063 14399
rect 23121 14365 23155 14399
rect 23397 14365 23431 14399
rect 23857 14365 23891 14399
rect 24041 14365 24075 14399
rect 24961 14365 24995 14399
rect 25329 14365 25363 14399
rect 26433 14365 26467 14399
rect 29009 14365 29043 14399
rect 31769 14365 31803 14399
rect 31953 14365 31987 14399
rect 32689 14365 32723 14399
rect 32965 14365 32999 14399
rect 33149 14365 33183 14399
rect 33609 14365 33643 14399
rect 37381 14365 37415 14399
rect 37565 14365 37599 14399
rect 38025 14365 38059 14399
rect 40049 14365 40083 14399
rect 42073 14365 42107 14399
rect 42349 14365 42383 14399
rect 57989 14365 58023 14399
rect 1869 14297 1903 14331
rect 11704 14297 11738 14331
rect 25145 14297 25179 14331
rect 25237 14297 25271 14331
rect 29193 14297 29227 14331
rect 29990 14297 30024 14331
rect 34345 14297 34379 14331
rect 37473 14297 37507 14331
rect 38270 14297 38304 14331
rect 40294 14297 40328 14331
rect 8493 14229 8527 14263
rect 10701 14229 10735 14263
rect 13645 14229 13679 14263
rect 15761 14229 15795 14263
rect 18153 14229 18187 14263
rect 20453 14229 20487 14263
rect 25513 14229 25547 14263
rect 31125 14229 31159 14263
rect 41429 14229 41463 14263
rect 44557 14229 44591 14263
rect 8861 14025 8895 14059
rect 9965 14025 9999 14059
rect 11713 14025 11747 14059
rect 13737 14025 13771 14059
rect 18779 14025 18813 14059
rect 22017 14025 22051 14059
rect 22385 14025 22419 14059
rect 22477 14025 22511 14059
rect 26157 14025 26191 14059
rect 28825 14025 28859 14059
rect 29377 14025 29411 14059
rect 32597 14025 32631 14059
rect 34897 14025 34931 14059
rect 37841 14025 37875 14059
rect 38025 14025 38059 14059
rect 39037 14025 39071 14059
rect 42073 14025 42107 14059
rect 19073 13957 19107 13991
rect 19257 13957 19291 13991
rect 1593 13889 1627 13923
rect 8677 13889 8711 13923
rect 9597 13889 9631 13923
rect 12081 13889 12115 13923
rect 12173 13889 12207 13923
rect 13369 13889 13403 13923
rect 14197 13889 14231 13923
rect 16865 13889 16899 13923
rect 17132 13889 17166 13923
rect 20269 13889 20303 13923
rect 21189 13889 21223 13923
rect 24777 13889 24811 13923
rect 24961 13889 24995 13923
rect 25053 13889 25087 13923
rect 25237 13889 25271 13923
rect 25329 13889 25363 13923
rect 28733 13889 28767 13923
rect 29745 13889 29779 13923
rect 31217 13889 31251 13923
rect 31585 13889 31619 13923
rect 31769 13889 31803 13923
rect 32321 13889 32355 13923
rect 32781 13889 32815 13923
rect 38022 13889 38056 13923
rect 38945 13889 38979 13923
rect 39129 13889 39163 13923
rect 41521 13889 41555 13923
rect 41705 13889 41739 13923
rect 41797 13889 41831 13923
rect 41889 13889 41923 13923
rect 43085 13889 43119 13923
rect 1777 13821 1811 13855
rect 2421 13821 2455 13855
rect 9505 13821 9539 13855
rect 10701 13821 10735 13855
rect 11897 13821 11931 13855
rect 11989 13821 12023 13855
rect 13461 13821 13495 13855
rect 14473 13821 14507 13855
rect 15853 13821 15887 13855
rect 19349 13821 19383 13855
rect 21005 13821 21039 13855
rect 22569 13821 22603 13855
rect 26249 13821 26283 13855
rect 26433 13821 26467 13855
rect 29837 13821 29871 13855
rect 30021 13821 30055 13855
rect 30573 13821 30607 13855
rect 31125 13821 31159 13855
rect 34989 13821 35023 13855
rect 35173 13821 35207 13855
rect 38485 13821 38519 13855
rect 43361 13821 43395 13855
rect 44741 13821 44775 13855
rect 10977 13753 11011 13787
rect 18245 13753 18279 13787
rect 38393 13753 38427 13787
rect 11161 13685 11195 13719
rect 20453 13685 20487 13719
rect 21373 13685 21407 13719
rect 25789 13685 25823 13719
rect 34529 13685 34563 13719
rect 9873 13481 9907 13515
rect 10885 13481 10919 13515
rect 13645 13481 13679 13515
rect 15025 13481 15059 13515
rect 22385 13481 22419 13515
rect 27353 13481 27387 13515
rect 32505 13481 32539 13515
rect 32781 13481 32815 13515
rect 43545 13481 43579 13515
rect 14473 13413 14507 13447
rect 16313 13413 16347 13447
rect 19625 13413 19659 13447
rect 32137 13413 32171 13447
rect 11897 13345 11931 13379
rect 15209 13345 15243 13379
rect 17325 13345 17359 13379
rect 20177 13345 20211 13379
rect 21005 13345 21039 13379
rect 32873 13345 32907 13379
rect 38669 13345 38703 13379
rect 58173 13345 58207 13379
rect 1593 13277 1627 13311
rect 9689 13277 9723 13311
rect 12633 13277 12667 13311
rect 13461 13277 13495 13311
rect 14289 13277 14323 13311
rect 15301 13277 15335 13311
rect 15393 13277 15427 13311
rect 15485 13277 15519 13311
rect 16037 13277 16071 13311
rect 17233 13277 17267 13311
rect 18245 13277 18279 13311
rect 18429 13277 18463 13311
rect 18521 13277 18555 13311
rect 19441 13277 19475 13311
rect 20361 13277 20395 13311
rect 21272 13277 21306 13311
rect 24777 13277 24811 13311
rect 30849 13277 30883 13311
rect 31585 13277 31619 13311
rect 31953 13277 31987 13311
rect 33057 13277 33091 13311
rect 36369 13277 36403 13311
rect 36461 13277 36495 13311
rect 38301 13277 38335 13311
rect 38761 13277 38795 13311
rect 42165 13277 42199 13311
rect 42349 13277 42383 13311
rect 42441 13277 42475 13311
rect 42533 13277 42567 13311
rect 43177 13277 43211 13311
rect 43361 13277 43395 13311
rect 57897 13277 57931 13311
rect 1869 13209 1903 13243
rect 10517 13209 10551 13243
rect 10701 13209 10735 13243
rect 12265 13209 12299 13243
rect 26065 13209 26099 13243
rect 31125 13209 31159 13243
rect 31769 13209 31803 13243
rect 31861 13209 31895 13243
rect 32781 13209 32815 13243
rect 57069 13209 57103 13243
rect 12081 13141 12115 13175
rect 12173 13141 12207 13175
rect 16497 13141 16531 13175
rect 17601 13141 17635 13175
rect 18061 13141 18095 13175
rect 20545 13141 20579 13175
rect 24869 13141 24903 13175
rect 33241 13141 33275 13175
rect 36645 13141 36679 13175
rect 42717 13141 42751 13175
rect 57161 13141 57195 13175
rect 10701 12937 10735 12971
rect 11897 12937 11931 12971
rect 14013 12937 14047 12971
rect 15209 12937 15243 12971
rect 19441 12937 19475 12971
rect 20177 12937 20211 12971
rect 20729 12937 20763 12971
rect 22937 12937 22971 12971
rect 27353 12937 27387 12971
rect 29929 12937 29963 12971
rect 31217 12937 31251 12971
rect 35173 12937 35207 12971
rect 41981 12937 42015 12971
rect 43177 12937 43211 12971
rect 14565 12869 14599 12903
rect 14933 12869 14967 12903
rect 17693 12869 17727 12903
rect 25136 12869 25170 12903
rect 28641 12869 28675 12903
rect 34060 12869 34094 12903
rect 36093 12869 36127 12903
rect 36185 12869 36219 12903
rect 10517 12801 10551 12835
rect 11713 12801 11747 12835
rect 12449 12801 12483 12835
rect 13829 12801 13863 12835
rect 14841 12801 14875 12835
rect 16037 12801 16071 12835
rect 17325 12801 17359 12835
rect 17509 12801 17543 12835
rect 18153 12801 18187 12835
rect 19282 12801 19316 12835
rect 19993 12801 20027 12835
rect 21097 12801 21131 12835
rect 22017 12801 22051 12835
rect 22753 12801 22787 12835
rect 24869 12801 24903 12835
rect 27261 12801 27295 12835
rect 27445 12801 27479 12835
rect 31033 12801 31067 12835
rect 31309 12801 31343 12835
rect 32597 12801 32631 12835
rect 32873 12801 32907 12835
rect 33793 12801 33827 12835
rect 35909 12801 35943 12835
rect 36277 12801 36311 12835
rect 41889 12801 41923 12835
rect 42809 12801 42843 12835
rect 42993 12801 43027 12835
rect 15025 12733 15059 12767
rect 21189 12733 21223 12767
rect 21373 12733 21407 12767
rect 33241 12733 33275 12767
rect 26249 12665 26283 12699
rect 32689 12665 32723 12699
rect 36461 12665 36495 12699
rect 12633 12597 12667 12631
rect 16221 12597 16255 12631
rect 18337 12597 18371 12631
rect 22201 12597 22235 12631
rect 30849 12597 30883 12631
rect 10609 12393 10643 12427
rect 11621 12393 11655 12427
rect 16037 12393 16071 12427
rect 17141 12393 17175 12427
rect 18613 12393 18647 12427
rect 22201 12393 22235 12427
rect 27629 12393 27663 12427
rect 30021 12393 30055 12427
rect 35817 12393 35851 12427
rect 37841 12393 37875 12427
rect 2329 12325 2363 12359
rect 25145 12325 25179 12359
rect 31033 12325 31067 12359
rect 13645 12257 13679 12291
rect 14381 12257 14415 12291
rect 25697 12257 25731 12291
rect 26617 12257 26651 12291
rect 36277 12257 36311 12291
rect 36553 12257 36587 12291
rect 2145 12189 2179 12223
rect 2605 12189 2639 12223
rect 10517 12189 10551 12223
rect 10701 12189 10735 12223
rect 11437 12189 11471 12223
rect 13553 12189 13587 12223
rect 13737 12189 13771 12223
rect 14473 12189 14507 12223
rect 15853 12189 15887 12223
rect 16957 12189 16991 12223
rect 17693 12189 17727 12223
rect 18429 12189 18463 12223
rect 20821 12189 20855 12223
rect 21088 12189 21122 12223
rect 24869 12189 24903 12223
rect 25145 12189 25179 12223
rect 25881 12189 25915 12223
rect 26525 12189 26559 12223
rect 27629 12189 27663 12223
rect 27813 12189 27847 12223
rect 30205 12189 30239 12223
rect 30481 12189 30515 12223
rect 31217 12189 31251 12223
rect 31309 12189 31343 12223
rect 31769 12189 31803 12223
rect 31953 12189 31987 12223
rect 35265 12189 35299 12223
rect 35541 12189 35575 12223
rect 35633 12189 35667 12223
rect 40049 12189 40083 12223
rect 40197 12189 40231 12223
rect 40417 12189 40451 12223
rect 40555 12189 40589 12223
rect 41153 12189 41187 12223
rect 41291 12189 41325 12223
rect 41429 12189 41463 12223
rect 41521 12189 41555 12223
rect 41637 12189 41671 12223
rect 57897 12189 57931 12223
rect 26801 12121 26835 12155
rect 31033 12121 31067 12155
rect 31861 12121 31895 12155
rect 35449 12121 35483 12155
rect 40325 12121 40359 12155
rect 58173 12121 58207 12155
rect 14841 12053 14875 12087
rect 17877 12053 17911 12087
rect 26065 12053 26099 12087
rect 26525 12053 26559 12087
rect 30389 12053 30423 12087
rect 40693 12053 40727 12087
rect 41797 12053 41831 12087
rect 14657 11849 14691 11883
rect 17417 11849 17451 11883
rect 18153 11849 18187 11883
rect 24593 11849 24627 11883
rect 24685 11849 24719 11883
rect 25329 11849 25363 11883
rect 25789 11849 25823 11883
rect 31401 11849 31435 11883
rect 33425 11849 33459 11883
rect 1869 11781 1903 11815
rect 15485 11781 15519 11815
rect 15685 11781 15719 11815
rect 24869 11781 24903 11815
rect 27414 11781 27448 11815
rect 46673 11781 46707 11815
rect 1593 11713 1627 11747
rect 11989 11713 12023 11747
rect 14473 11713 14507 11747
rect 17233 11713 17267 11747
rect 17969 11713 18003 11747
rect 20361 11713 20395 11747
rect 24501 11713 24535 11747
rect 25697 11713 25731 11747
rect 29561 11713 29595 11747
rect 29653 11713 29687 11747
rect 29837 11713 29871 11747
rect 29929 11713 29963 11747
rect 30665 11713 30699 11747
rect 31309 11713 31343 11747
rect 31493 11713 31527 11747
rect 32965 11713 32999 11747
rect 33241 11713 33275 11747
rect 34621 11713 34655 11747
rect 34888 11713 34922 11747
rect 38761 11713 38795 11747
rect 57161 11713 57195 11747
rect 11713 11645 11747 11679
rect 11897 11645 11931 11679
rect 12081 11645 12115 11679
rect 12173 11645 12207 11679
rect 20453 11645 20487 11679
rect 20637 11645 20671 11679
rect 25973 11645 26007 11679
rect 27169 11645 27203 11679
rect 33057 11645 33091 11679
rect 46765 11645 46799 11679
rect 46857 11645 46891 11679
rect 24317 11577 24351 11611
rect 40049 11577 40083 11611
rect 15669 11509 15703 11543
rect 15853 11509 15887 11543
rect 19993 11509 20027 11543
rect 28549 11509 28583 11543
rect 29377 11509 29411 11543
rect 30757 11509 30791 11543
rect 36001 11509 36035 11543
rect 46305 11509 46339 11543
rect 57253 11509 57287 11543
rect 18797 11305 18831 11339
rect 21005 11305 21039 11339
rect 26433 11305 26467 11339
rect 35265 11305 35299 11339
rect 15117 11237 15151 11271
rect 21649 11237 21683 11271
rect 31309 11237 31343 11271
rect 46949 11237 46983 11271
rect 53665 11237 53699 11271
rect 56149 11237 56183 11271
rect 58265 11237 58299 11271
rect 1777 11169 1811 11203
rect 10977 11169 11011 11203
rect 11161 11169 11195 11203
rect 11253 11169 11287 11203
rect 11345 11169 11379 11203
rect 13185 11169 13219 11203
rect 16405 11169 16439 11203
rect 27813 11169 27847 11203
rect 30113 11169 30147 11203
rect 33425 11169 33459 11203
rect 35817 11169 35851 11203
rect 41429 11169 41463 11203
rect 43269 11169 43303 11203
rect 1593 11101 1627 11135
rect 11437 11101 11471 11135
rect 13001 11101 13035 11135
rect 14933 11101 14967 11135
rect 16313 11101 16347 11135
rect 16681 11101 16715 11135
rect 16865 11101 16899 11135
rect 18613 11101 18647 11135
rect 19625 11101 19659 11135
rect 21465 11101 21499 11135
rect 24777 11101 24811 11135
rect 26249 11101 26283 11135
rect 27353 11101 27387 11135
rect 29745 11101 29779 11135
rect 31585 11101 31619 11135
rect 32045 11101 32079 11135
rect 32137 11101 32171 11135
rect 32965 11101 32999 11135
rect 35633 11101 35667 11135
rect 38485 11101 38519 11135
rect 41521 11101 41555 11135
rect 41889 11101 41923 11135
rect 42073 11101 42107 11135
rect 43177 11101 43211 11135
rect 43545 11101 43579 11135
rect 43637 11101 43671 11135
rect 44189 11101 44223 11135
rect 45569 11101 45603 11135
rect 53113 11101 53147 11135
rect 53297 11101 53331 11135
rect 53481 11101 53515 11135
rect 56149 11101 56183 11135
rect 56425 11101 56459 11135
rect 56885 11101 56919 11135
rect 57141 11101 57175 11135
rect 15669 11033 15703 11067
rect 17509 11033 17543 11067
rect 19881 11033 19915 11067
rect 25605 11033 25639 11067
rect 31309 11033 31343 11067
rect 35725 11033 35759 11067
rect 38301 11033 38335 11067
rect 38853 11033 38887 11067
rect 40877 11033 40911 11067
rect 42533 11033 42567 11067
rect 44465 11033 44499 11067
rect 45836 11033 45870 11067
rect 53389 11033 53423 11067
rect 56333 11033 56367 11067
rect 17601 10965 17635 10999
rect 31493 10965 31527 10999
rect 9321 10761 9355 10795
rect 12173 10761 12207 10795
rect 18521 10761 18555 10795
rect 18889 10761 18923 10795
rect 21097 10761 21131 10795
rect 22017 10761 22051 10795
rect 22385 10761 22419 10795
rect 23581 10761 23615 10795
rect 31217 10761 31251 10795
rect 33793 10761 33827 10795
rect 34805 10761 34839 10795
rect 45477 10761 45511 10795
rect 57253 10761 57287 10795
rect 1869 10693 1903 10727
rect 17049 10693 17083 10727
rect 19962 10693 19996 10727
rect 26341 10693 26375 10727
rect 34437 10693 34471 10727
rect 34529 10693 34563 10727
rect 35265 10693 35299 10727
rect 38209 10693 38243 10727
rect 38301 10693 38335 10727
rect 1593 10625 1627 10659
rect 9505 10625 9539 10659
rect 9598 10625 9632 10659
rect 9781 10625 9815 10659
rect 11713 10625 11747 10659
rect 12909 10625 12943 10659
rect 13185 10625 13219 10659
rect 14749 10625 14783 10659
rect 14933 10625 14967 10659
rect 15669 10625 15703 10659
rect 17417 10625 17451 10659
rect 17509 10625 17543 10659
rect 19717 10625 19751 10659
rect 23397 10625 23431 10659
rect 23581 10625 23615 10659
rect 24501 10625 24535 10659
rect 24869 10625 24903 10659
rect 25697 10625 25731 10659
rect 27721 10625 27755 10659
rect 27905 10625 27939 10659
rect 28089 10625 28123 10659
rect 28556 10625 28590 10659
rect 28825 10625 28859 10659
rect 31158 10625 31192 10659
rect 33149 10625 33183 10659
rect 33297 10625 33331 10659
rect 33425 10625 33459 10659
rect 33517 10625 33551 10659
rect 33655 10625 33689 10659
rect 34253 10625 34287 10659
rect 34621 10625 34655 10659
rect 35449 10625 35483 10659
rect 35541 10625 35575 10659
rect 38025 10625 38059 10659
rect 38393 10625 38427 10659
rect 40960 10625 40994 10659
rect 44189 10625 44223 10659
rect 57161 10625 57195 10659
rect 57345 10625 57379 10659
rect 9689 10557 9723 10591
rect 13369 10557 13403 10591
rect 15945 10557 15979 10591
rect 16957 10557 16991 10591
rect 17969 10557 18003 10591
rect 18981 10557 19015 10591
rect 19165 10557 19199 10591
rect 22477 10557 22511 10591
rect 22569 10557 22603 10591
rect 24961 10557 24995 10591
rect 31585 10557 31619 10591
rect 31677 10557 31711 10591
rect 40693 10557 40727 10591
rect 11989 10489 12023 10523
rect 13001 10489 13035 10523
rect 15117 10489 15151 10523
rect 24317 10489 24351 10523
rect 31033 10489 31067 10523
rect 14841 10421 14875 10455
rect 29929 10421 29963 10455
rect 35541 10421 35575 10455
rect 35725 10421 35759 10455
rect 38577 10421 38611 10455
rect 42073 10421 42107 10455
rect 11529 10217 11563 10251
rect 31953 10217 31987 10251
rect 41337 10217 41371 10251
rect 11345 10149 11379 10183
rect 12909 10149 12943 10183
rect 16957 10149 16991 10183
rect 21189 10149 21223 10183
rect 24758 10149 24792 10183
rect 24869 10149 24903 10183
rect 27721 10149 27755 10183
rect 1777 10081 1811 10115
rect 18337 10081 18371 10115
rect 19809 10081 19843 10115
rect 22201 10081 22235 10115
rect 23673 10081 23707 10115
rect 24961 10081 24995 10115
rect 25789 10081 25823 10115
rect 29745 10081 29779 10115
rect 37657 10081 37691 10115
rect 41797 10081 41831 10115
rect 41981 10081 42015 10115
rect 45661 10081 45695 10115
rect 58173 10081 58207 10115
rect 1593 10013 1627 10047
rect 11069 10013 11103 10047
rect 12817 10013 12851 10047
rect 13093 10013 13127 10047
rect 14381 10013 14415 10047
rect 15853 10013 15887 10047
rect 16313 10013 16347 10047
rect 16405 10013 16439 10047
rect 16773 10013 16807 10047
rect 17693 10013 17727 10047
rect 20076 10013 20110 10047
rect 22109 10013 22143 10047
rect 23857 10013 23891 10047
rect 25329 10013 25363 10047
rect 26065 10013 26099 10047
rect 26341 10013 26375 10047
rect 26525 10013 26559 10047
rect 26801 10013 26835 10047
rect 27905 10013 27939 10047
rect 28017 10013 28051 10047
rect 28129 10013 28163 10047
rect 28733 10013 28767 10047
rect 32137 10013 32171 10047
rect 32413 10013 32447 10047
rect 35081 10013 35115 10047
rect 37381 10013 37415 10047
rect 38301 10013 38335 10047
rect 38439 10013 38473 10047
rect 38577 10013 38611 10047
rect 38766 10013 38800 10047
rect 44189 10013 44223 10047
rect 44281 10013 44315 10047
rect 44373 10013 44407 10047
rect 44557 10013 44591 10047
rect 45845 10013 45879 10047
rect 46121 10013 46155 10047
rect 57897 10013 57931 10047
rect 14933 9945 14967 9979
rect 24041 9945 24075 9979
rect 24593 9945 24627 9979
rect 28273 9945 28307 9979
rect 29009 9945 29043 9979
rect 29929 9945 29963 9979
rect 30297 9945 30331 9979
rect 35265 9945 35299 9979
rect 35449 9945 35483 9979
rect 38669 9945 38703 9979
rect 41705 9945 41739 9979
rect 46857 9945 46891 9979
rect 57069 9945 57103 9979
rect 13277 9877 13311 9911
rect 21649 9877 21683 9911
rect 22017 9877 22051 9911
rect 27169 9877 27203 9911
rect 30021 9877 30055 9911
rect 30113 9877 30147 9911
rect 32321 9877 32355 9911
rect 38945 9877 38979 9911
rect 43913 9877 43947 9911
rect 46029 9877 46063 9911
rect 48145 9877 48179 9911
rect 57161 9877 57195 9911
rect 27537 9673 27571 9707
rect 28825 9673 28859 9707
rect 29837 9673 29871 9707
rect 32505 9673 32539 9707
rect 46581 9673 46615 9707
rect 20076 9605 20110 9639
rect 24685 9605 24719 9639
rect 28743 9605 28777 9639
rect 29469 9605 29503 9639
rect 43729 9605 43763 9639
rect 45468 9605 45502 9639
rect 1593 9537 1627 9571
rect 13369 9537 13403 9571
rect 13461 9537 13495 9571
rect 13645 9537 13679 9571
rect 13737 9537 13771 9571
rect 15209 9537 15243 9571
rect 15485 9537 15519 9571
rect 15577 9537 15611 9571
rect 15853 9537 15887 9571
rect 16129 9537 16163 9571
rect 17049 9537 17083 9571
rect 18705 9537 18739 9571
rect 23949 9537 23983 9571
rect 25237 9537 25271 9571
rect 25329 9537 25363 9571
rect 25605 9537 25639 9571
rect 27169 9537 27203 9571
rect 28641 9537 28675 9571
rect 29009 9537 29043 9571
rect 29653 9537 29687 9571
rect 29791 9537 29825 9571
rect 30021 9537 30055 9571
rect 30941 9537 30975 9571
rect 32597 9537 32631 9571
rect 32781 9537 32815 9571
rect 33333 9537 33367 9571
rect 36001 9537 36035 9571
rect 36185 9537 36219 9571
rect 37473 9537 37507 9571
rect 37621 9537 37655 9571
rect 37749 9537 37783 9571
rect 37841 9537 37875 9571
rect 37938 9537 37972 9571
rect 40509 9537 40543 9571
rect 43913 9537 43947 9571
rect 44005 9537 44039 9571
rect 44097 9537 44131 9571
rect 45201 9537 45235 9571
rect 57069 9537 57103 9571
rect 57253 9537 57287 9571
rect 1777 9469 1811 9503
rect 8769 9469 8803 9503
rect 9229 9469 9263 9503
rect 17785 9469 17819 9503
rect 19809 9469 19843 9503
rect 25789 9469 25823 9503
rect 26065 9469 26099 9503
rect 27261 9469 27295 9503
rect 33517 9469 33551 9503
rect 9045 9401 9079 9435
rect 18797 9401 18831 9435
rect 24133 9401 24167 9435
rect 28457 9401 28491 9435
rect 13185 9333 13219 9367
rect 14841 9333 14875 9367
rect 21189 9333 21223 9367
rect 27353 9333 27387 9367
rect 31217 9333 31251 9367
rect 32321 9333 32355 9367
rect 36001 9333 36035 9367
rect 38117 9333 38151 9367
rect 40601 9333 40635 9367
rect 44281 9333 44315 9367
rect 57161 9333 57195 9367
rect 28457 9129 28491 9163
rect 37749 9129 37783 9163
rect 41429 9129 41463 9163
rect 13093 9061 13127 9095
rect 13277 9061 13311 9095
rect 16957 9061 16991 9095
rect 21557 9061 21591 9095
rect 33057 9061 33091 9095
rect 33977 9061 34011 9095
rect 38669 9061 38703 9095
rect 56149 9061 56183 9095
rect 18061 8993 18095 9027
rect 19533 8993 19567 9027
rect 24777 8993 24811 9027
rect 26433 8993 26467 9027
rect 29009 8993 29043 9027
rect 36277 8993 36311 9027
rect 40049 8993 40083 9027
rect 56885 8993 56919 9027
rect 1593 8925 1627 8959
rect 16037 8925 16071 8959
rect 16405 8925 16439 8959
rect 16681 8925 16715 8959
rect 17417 8925 17451 8959
rect 18429 8925 18463 8959
rect 21373 8925 21407 8959
rect 24041 8925 24075 8959
rect 24593 8925 24627 8959
rect 25145 8925 25179 8959
rect 25881 8925 25915 8959
rect 25973 8925 26007 8959
rect 27813 8925 27847 8959
rect 27997 8925 28031 8959
rect 31125 8925 31159 8959
rect 31309 8925 31343 8959
rect 32137 8925 32171 8959
rect 33333 8925 33367 8959
rect 33517 8925 33551 8959
rect 34161 8925 34195 8959
rect 34253 8925 34287 8959
rect 35817 8925 35851 8959
rect 36369 8925 36403 8959
rect 37197 8925 37231 8959
rect 37473 8925 37507 8959
rect 37565 8925 37599 8959
rect 38853 8925 38887 8959
rect 44465 8925 44499 8959
rect 45201 8925 45235 8959
rect 46121 8925 46155 8959
rect 46305 8925 46339 8959
rect 56149 8925 56183 8959
rect 56333 8925 56367 8959
rect 56425 8925 56459 8959
rect 57141 8925 57175 8959
rect 1869 8857 1903 8891
rect 12817 8857 12851 8891
rect 14933 8857 14967 8891
rect 15301 8857 15335 8891
rect 17969 8857 18003 8891
rect 18521 8857 18555 8891
rect 18613 8857 18647 8891
rect 19800 8857 19834 8891
rect 23489 8857 23523 8891
rect 23673 8857 23707 8891
rect 25329 8857 25363 8891
rect 28917 8857 28951 8891
rect 29745 8857 29779 8891
rect 30481 8857 30515 8891
rect 31677 8857 31711 8891
rect 32413 8857 32447 8891
rect 33977 8857 34011 8891
rect 37381 8857 37415 8891
rect 40316 8857 40350 8891
rect 43729 8857 43763 8891
rect 45477 8857 45511 8891
rect 14841 8789 14875 8823
rect 15025 8789 15059 8823
rect 15117 8789 15151 8823
rect 20913 8789 20947 8823
rect 23765 8789 23799 8823
rect 23857 8789 23891 8823
rect 25237 8789 25271 8823
rect 28825 8789 28859 8823
rect 31401 8789 31435 8823
rect 31493 8789 31527 8823
rect 33241 8789 33275 8823
rect 36001 8789 36035 8823
rect 46305 8789 46339 8823
rect 58265 8789 58299 8823
rect 14105 8585 14139 8619
rect 15025 8585 15059 8619
rect 17417 8585 17451 8619
rect 17509 8585 17543 8619
rect 19349 8585 19383 8619
rect 20269 8585 20303 8619
rect 20637 8585 20671 8619
rect 23581 8585 23615 8619
rect 23673 8585 23707 8619
rect 25329 8585 25363 8619
rect 25973 8585 26007 8619
rect 26157 8585 26191 8619
rect 31309 8585 31343 8619
rect 31401 8585 31435 8619
rect 33425 8585 33459 8619
rect 38761 8585 38795 8619
rect 40049 8585 40083 8619
rect 44281 8585 44315 8619
rect 16957 8517 16991 8551
rect 20729 8517 20763 8551
rect 23305 8517 23339 8551
rect 26267 8517 26301 8551
rect 26433 8517 26467 8551
rect 27537 8517 27571 8551
rect 28917 8517 28951 8551
rect 31033 8517 31067 8551
rect 31217 8517 31251 8551
rect 33149 8517 33183 8551
rect 39865 8517 39899 8551
rect 43177 8517 43211 8551
rect 57345 8517 57379 8551
rect 1593 8449 1627 8483
rect 14013 8449 14047 8483
rect 14933 8449 14967 8483
rect 15669 8449 15703 8483
rect 17693 8449 17727 8483
rect 18245 8449 18279 8483
rect 18613 8449 18647 8483
rect 18981 8449 19015 8483
rect 19809 8449 19843 8483
rect 23489 8449 23523 8483
rect 23857 8449 23891 8483
rect 24317 8449 24351 8483
rect 24501 8449 24535 8483
rect 25145 8449 25179 8483
rect 26065 8449 26099 8483
rect 27353 8449 27387 8483
rect 27629 8449 27663 8483
rect 27721 8449 27755 8483
rect 28457 8449 28491 8483
rect 29561 8449 29595 8483
rect 31585 8449 31619 8483
rect 32781 8449 32815 8483
rect 32874 8449 32908 8483
rect 33057 8449 33091 8483
rect 33246 8449 33280 8483
rect 33885 8449 33919 8483
rect 33978 8449 34012 8483
rect 34161 8449 34195 8483
rect 34253 8449 34287 8483
rect 34350 8449 34384 8483
rect 35909 8449 35943 8483
rect 36737 8449 36771 8483
rect 37473 8449 37507 8483
rect 37565 8449 37599 8483
rect 37749 8449 37783 8483
rect 38209 8449 38243 8483
rect 38945 8449 38979 8483
rect 39221 8449 39255 8483
rect 39405 8449 39439 8483
rect 40141 8449 40175 8483
rect 42809 8449 42843 8483
rect 44465 8449 44499 8483
rect 44557 8449 44591 8483
rect 44741 8449 44775 8483
rect 44833 8449 44867 8483
rect 45293 8449 45327 8483
rect 46397 8449 46431 8483
rect 56241 8449 56275 8483
rect 57069 8449 57103 8483
rect 1777 8381 1811 8415
rect 16221 8381 16255 8415
rect 20913 8381 20947 8415
rect 29929 8381 29963 8415
rect 35357 8381 35391 8415
rect 35725 8381 35759 8415
rect 35817 8381 35851 8415
rect 36553 8381 36587 8415
rect 45477 8381 45511 8415
rect 46581 8381 46615 8415
rect 16957 8313 16991 8347
rect 24593 8313 24627 8347
rect 34529 8313 34563 8347
rect 39037 8313 39071 8347
rect 39129 8313 39163 8347
rect 39865 8313 39899 8347
rect 56425 8313 56459 8347
rect 27905 8245 27939 8279
rect 36921 8245 36955 8279
rect 15945 8041 15979 8075
rect 25053 8041 25087 8075
rect 25789 8041 25823 8075
rect 28733 8041 28767 8075
rect 34161 8041 34195 8075
rect 38669 8041 38703 8075
rect 42717 8041 42751 8075
rect 44281 8041 44315 8075
rect 45385 8041 45419 8075
rect 12909 7973 12943 8007
rect 13093 7973 13127 8007
rect 17693 7973 17727 8007
rect 28622 7973 28656 8007
rect 56149 7973 56183 8007
rect 8585 7905 8619 7939
rect 12633 7905 12667 7939
rect 15577 7905 15611 7939
rect 23305 7905 23339 7939
rect 24961 7905 24995 7939
rect 28825 7905 28859 7939
rect 30205 7905 30239 7939
rect 30941 7905 30975 7939
rect 31493 7905 31527 7939
rect 32689 7905 32723 7939
rect 46581 7905 46615 7939
rect 56885 7905 56919 7939
rect 1593 7837 1627 7871
rect 7849 7837 7883 7871
rect 7941 7837 7975 7871
rect 8125 7837 8159 7871
rect 10057 7837 10091 7871
rect 10977 7837 11011 7871
rect 15301 7837 15335 7871
rect 15669 7837 15703 7871
rect 16589 7837 16623 7871
rect 17141 7837 17175 7871
rect 17509 7837 17543 7871
rect 18061 7837 18095 7871
rect 19533 7837 19567 7871
rect 24593 7837 24627 7871
rect 25605 7837 25639 7871
rect 26709 7837 26743 7871
rect 30021 7837 30055 7871
rect 30113 7837 30147 7871
rect 31401 7837 31435 7871
rect 31677 7837 31711 7871
rect 32873 7837 32907 7871
rect 34161 7837 34195 7871
rect 34345 7837 34379 7871
rect 34989 7837 35023 7871
rect 36093 7837 36127 7871
rect 36360 7837 36394 7871
rect 38025 7837 38059 7871
rect 38118 7837 38152 7871
rect 38393 7837 38427 7871
rect 38490 7837 38524 7871
rect 42625 7837 42659 7871
rect 43821 7837 43855 7871
rect 44005 7837 44039 7871
rect 44097 7837 44131 7871
rect 45569 7837 45603 7871
rect 46305 7837 46339 7871
rect 55505 7837 55539 7871
rect 55689 7837 55723 7871
rect 56425 7837 56459 7871
rect 57141 7837 57175 7871
rect 1869 7769 1903 7803
rect 9873 7769 9907 7803
rect 10333 7769 10367 7803
rect 11989 7769 12023 7803
rect 15761 7769 15795 7803
rect 19901 7769 19935 7803
rect 27537 7769 27571 7803
rect 28457 7769 28491 7803
rect 30481 7769 30515 7803
rect 33149 7769 33183 7803
rect 38301 7769 38335 7803
rect 45293 7769 45327 7803
rect 45477 7769 45511 7803
rect 56149 7769 56183 7803
rect 10241 7701 10275 7735
rect 22661 7701 22695 7735
rect 23029 7701 23063 7735
rect 23121 7701 23155 7735
rect 24777 7701 24811 7735
rect 29101 7701 29135 7735
rect 31861 7701 31895 7735
rect 33057 7701 33091 7735
rect 35081 7701 35115 7735
rect 37473 7701 37507 7735
rect 55689 7701 55723 7735
rect 56333 7701 56367 7735
rect 58265 7701 58299 7735
rect 10609 7497 10643 7531
rect 18613 7497 18647 7531
rect 22201 7497 22235 7531
rect 24685 7497 24719 7531
rect 25973 7497 26007 7531
rect 29929 7497 29963 7531
rect 35541 7497 35575 7531
rect 36185 7497 36219 7531
rect 37565 7497 37599 7531
rect 11989 7429 12023 7463
rect 15117 7429 15151 7463
rect 15209 7429 15243 7463
rect 15669 7429 15703 7463
rect 16957 7429 16991 7463
rect 18521 7429 18555 7463
rect 28641 7429 28675 7463
rect 36553 7429 36587 7463
rect 44557 7429 44591 7463
rect 46213 7429 46247 7463
rect 55781 7429 55815 7463
rect 56977 7429 57011 7463
rect 10793 7361 10827 7395
rect 10977 7361 11011 7395
rect 11805 7361 11839 7395
rect 12449 7361 12483 7395
rect 15577 7361 15611 7395
rect 16129 7361 16163 7395
rect 17417 7361 17451 7395
rect 17509 7361 17543 7395
rect 20352 7361 20386 7395
rect 22023 7361 22057 7395
rect 23397 7361 23431 7395
rect 27629 7361 27663 7395
rect 31217 7361 31251 7395
rect 34428 7361 34462 7395
rect 36645 7361 36679 7395
rect 37473 7361 37507 7395
rect 37657 7361 37691 7395
rect 44465 7361 44499 7395
rect 45201 7361 45235 7395
rect 45385 7361 45419 7395
rect 46305 7361 46339 7395
rect 55965 7361 55999 7395
rect 56057 7361 56091 7395
rect 56609 7361 56643 7395
rect 58081 7361 58115 7395
rect 58265 7361 58299 7395
rect 10885 7293 10919 7327
rect 11069 7293 11103 7327
rect 12909 7293 12943 7327
rect 17049 7293 17083 7327
rect 17969 7293 18003 7327
rect 20085 7293 20119 7327
rect 27721 7293 27755 7327
rect 31309 7293 31343 7327
rect 31493 7293 31527 7327
rect 34161 7293 34195 7327
rect 36829 7293 36863 7327
rect 45293 7293 45327 7327
rect 46489 7293 46523 7327
rect 12725 7225 12759 7259
rect 25605 7225 25639 7259
rect 58173 7225 58207 7259
rect 21465 7157 21499 7191
rect 25973 7157 26007 7191
rect 26157 7157 26191 7191
rect 27813 7157 27847 7191
rect 27997 7157 28031 7191
rect 30849 7157 30883 7191
rect 45845 7157 45879 7191
rect 55781 7157 55815 7191
rect 13645 6953 13679 6987
rect 20729 6953 20763 6987
rect 28135 6953 28169 6987
rect 28273 6953 28307 6987
rect 34345 6953 34379 6987
rect 46581 6953 46615 6987
rect 1777 6817 1811 6851
rect 10793 6817 10827 6851
rect 11069 6817 11103 6851
rect 16037 6817 16071 6851
rect 16129 6817 16163 6851
rect 17693 6817 17727 6851
rect 21281 6817 21315 6851
rect 22477 6817 22511 6851
rect 25421 6817 25455 6851
rect 26525 6817 26559 6851
rect 28365 6817 28399 6851
rect 30113 6817 30147 6851
rect 33977 6817 34011 6851
rect 35541 6817 35575 6851
rect 47409 6817 47443 6851
rect 56885 6817 56919 6851
rect 1593 6749 1627 6783
rect 9505 6749 9539 6783
rect 10977 6749 11011 6783
rect 11161 6749 11195 6783
rect 11253 6749 11287 6783
rect 16497 6749 16531 6783
rect 16589 6749 16623 6783
rect 17417 6749 17451 6783
rect 19625 6749 19659 6783
rect 22744 6749 22778 6783
rect 25973 6749 26007 6783
rect 26617 6749 26651 6783
rect 26985 6749 27019 6783
rect 27077 6749 27111 6783
rect 29745 6749 29779 6783
rect 31401 6749 31435 6783
rect 34161 6749 34195 6783
rect 45201 6749 45235 6783
rect 57141 6749 57175 6783
rect 13553 6681 13587 6715
rect 14381 6681 14415 6715
rect 16681 6681 16715 6715
rect 19993 6681 20027 6715
rect 21097 6681 21131 6715
rect 27997 6681 28031 6715
rect 31217 6681 31251 6715
rect 31769 6681 31803 6715
rect 45468 6681 45502 6715
rect 47133 6681 47167 6715
rect 9689 6613 9723 6647
rect 14473 6613 14507 6647
rect 21189 6613 21223 6647
rect 23857 6613 23891 6647
rect 24777 6613 24811 6647
rect 25145 6613 25179 6647
rect 25237 6613 25271 6647
rect 28641 6613 28675 6647
rect 31493 6613 31527 6647
rect 31585 6613 31619 6647
rect 34897 6613 34931 6647
rect 35265 6613 35299 6647
rect 35357 6613 35391 6647
rect 58265 6613 58299 6647
rect 9137 6409 9171 6443
rect 13185 6409 13219 6443
rect 23029 6409 23063 6443
rect 28089 6409 28123 6443
rect 35633 6409 35667 6443
rect 36553 6409 36587 6443
rect 38761 6409 38795 6443
rect 13737 6341 13771 6375
rect 15301 6341 15335 6375
rect 16865 6341 16899 6375
rect 18521 6341 18555 6375
rect 23489 6341 23523 6375
rect 25044 6341 25078 6375
rect 29009 6341 29043 6375
rect 34805 6341 34839 6375
rect 35541 6341 35575 6375
rect 1593 6273 1627 6307
rect 9413 6273 9447 6307
rect 13001 6273 13035 6307
rect 15393 6273 15427 6307
rect 15761 6273 15795 6307
rect 15853 6273 15887 6307
rect 16313 6273 16347 6307
rect 17601 6273 17635 6307
rect 18245 6273 18279 6307
rect 19441 6273 19475 6307
rect 19708 6273 19742 6307
rect 22017 6273 22051 6307
rect 23397 6273 23431 6307
rect 24777 6273 24811 6307
rect 27537 6273 27571 6307
rect 28641 6273 28675 6307
rect 29745 6273 29779 6307
rect 30021 6273 30055 6307
rect 30941 6273 30975 6307
rect 31125 6273 31159 6307
rect 34529 6273 34563 6307
rect 36461 6273 36495 6307
rect 38577 6273 38611 6307
rect 46305 6273 46339 6307
rect 46397 6273 46431 6307
rect 58081 6273 58115 6307
rect 1777 6205 1811 6239
rect 9321 6205 9355 6239
rect 9505 6205 9539 6239
rect 9597 6205 9631 6239
rect 23673 6205 23707 6239
rect 27813 6205 27847 6239
rect 30205 6205 30239 6239
rect 46581 6205 46615 6239
rect 14013 6137 14047 6171
rect 14197 6137 14231 6171
rect 20821 6137 20855 6171
rect 29837 6137 29871 6171
rect 22201 6069 22235 6103
rect 26157 6069 26191 6103
rect 27905 6069 27939 6103
rect 31309 6069 31343 6103
rect 58265 6069 58299 6103
rect 9137 5865 9171 5899
rect 10885 5865 10919 5899
rect 23581 5865 23615 5899
rect 25145 5865 25179 5899
rect 25789 5865 25823 5899
rect 32689 5865 32723 5899
rect 37381 5865 37415 5899
rect 38025 5865 38059 5899
rect 10701 5797 10735 5831
rect 17969 5797 18003 5831
rect 22017 5797 22051 5831
rect 29101 5797 29135 5831
rect 29837 5797 29871 5831
rect 30757 5797 30791 5831
rect 41613 5797 41647 5831
rect 9413 5729 9447 5763
rect 19809 5729 19843 5763
rect 22477 5729 22511 5763
rect 22661 5729 22695 5763
rect 26341 5729 26375 5763
rect 31309 5729 31343 5763
rect 33609 5729 33643 5763
rect 36461 5729 36495 5763
rect 36645 5729 36679 5763
rect 38393 5729 38427 5763
rect 39221 5729 39255 5763
rect 39405 5729 39439 5763
rect 57253 5729 57287 5763
rect 1593 5661 1627 5695
rect 9321 5661 9355 5695
rect 9505 5661 9539 5695
rect 9597 5661 9631 5695
rect 17049 5661 17083 5695
rect 17417 5661 17451 5695
rect 17785 5661 17819 5695
rect 18429 5661 18463 5695
rect 20076 5661 20110 5695
rect 23305 5661 23339 5695
rect 24961 5661 24995 5695
rect 28549 5661 28583 5695
rect 28922 5661 28956 5695
rect 29653 5661 29687 5695
rect 30297 5661 30331 5695
rect 30573 5661 30607 5695
rect 31565 5661 31599 5695
rect 34161 5661 34195 5695
rect 34345 5661 34379 5695
rect 56977 5661 57011 5695
rect 57897 5661 57931 5695
rect 58173 5661 58207 5695
rect 1869 5593 1903 5627
rect 10425 5593 10459 5627
rect 26157 5593 26191 5627
rect 28733 5593 28767 5627
rect 28825 5593 28859 5627
rect 33425 5593 33459 5627
rect 34989 5593 35023 5627
rect 35173 5593 35207 5627
rect 37289 5593 37323 5627
rect 37933 5593 37967 5627
rect 39129 5593 39163 5627
rect 41429 5593 41463 5627
rect 21189 5525 21223 5559
rect 22385 5525 22419 5559
rect 26249 5525 26283 5559
rect 35725 5525 35759 5559
rect 36001 5525 36035 5559
rect 36369 5525 36403 5559
rect 38761 5525 38795 5559
rect 9413 5321 9447 5355
rect 10241 5321 10275 5355
rect 13829 5321 13863 5355
rect 19625 5321 19659 5355
rect 25789 5321 25823 5355
rect 29377 5321 29411 5355
rect 30757 5321 30791 5355
rect 40601 5321 40635 5355
rect 42809 5321 42843 5355
rect 58265 5321 58299 5355
rect 19993 5253 20027 5287
rect 20085 5253 20119 5287
rect 30021 5253 30055 5287
rect 1593 5185 1627 5219
rect 8217 5185 8251 5219
rect 10425 5185 10459 5219
rect 12449 5185 12483 5219
rect 13369 5185 13403 5219
rect 14381 5185 14415 5219
rect 18705 5185 18739 5219
rect 21005 5185 21039 5219
rect 22569 5185 22603 5219
rect 23673 5185 23707 5219
rect 25605 5185 25639 5219
rect 28365 5185 28399 5219
rect 28457 5185 28491 5219
rect 29193 5185 29227 5219
rect 30665 5185 30699 5219
rect 30849 5185 30883 5219
rect 32873 5185 32907 5219
rect 33609 5185 33643 5219
rect 34345 5185 34379 5219
rect 35173 5185 35207 5219
rect 35817 5185 35851 5219
rect 37565 5185 37599 5219
rect 38752 5185 38786 5219
rect 40417 5185 40451 5219
rect 41245 5185 41279 5219
rect 42717 5185 42751 5219
rect 43453 5185 43487 5219
rect 44189 5185 44223 5219
rect 44925 5185 44959 5219
rect 45845 5185 45879 5219
rect 48513 5185 48547 5219
rect 48769 5185 48803 5219
rect 58081 5185 58115 5219
rect 1777 5117 1811 5151
rect 8953 5117 8987 5151
rect 10517 5117 10551 5151
rect 10609 5117 10643 5151
rect 10701 5117 10735 5151
rect 18889 5117 18923 5151
rect 20269 5117 20303 5151
rect 21189 5117 21223 5151
rect 22753 5117 22787 5151
rect 23857 5117 23891 5151
rect 28641 5117 28675 5151
rect 33057 5117 33091 5151
rect 34989 5117 35023 5151
rect 36001 5117 36035 5151
rect 38485 5117 38519 5151
rect 46029 5117 46063 5151
rect 9229 5049 9263 5083
rect 13645 5049 13679 5083
rect 17877 5049 17911 5083
rect 34529 5049 34563 5083
rect 43637 5049 43671 5083
rect 8401 4981 8435 5015
rect 12541 4981 12575 5015
rect 14473 4981 14507 5015
rect 16313 4981 16347 5015
rect 17233 4981 17267 5015
rect 26525 4981 26559 5015
rect 27997 4981 28031 5015
rect 30113 4981 30147 5015
rect 33701 4981 33735 5015
rect 35357 4981 35391 5015
rect 37657 4981 37691 5015
rect 39865 4981 39899 5015
rect 41337 4981 41371 5015
rect 44281 4981 44315 5015
rect 45017 4981 45051 5015
rect 49893 4981 49927 5015
rect 9689 4777 9723 4811
rect 11161 4777 11195 4811
rect 19441 4777 19475 4811
rect 37105 4777 37139 4811
rect 39129 4777 39163 4811
rect 40233 4777 40267 4811
rect 41705 4777 41739 4811
rect 58265 4777 58299 4811
rect 7113 4709 7147 4743
rect 8585 4709 8619 4743
rect 10977 4709 11011 4743
rect 13461 4709 13495 4743
rect 13645 4709 13679 4743
rect 14565 4709 14599 4743
rect 32321 4709 32355 4743
rect 44465 4709 44499 4743
rect 45477 4709 45511 4743
rect 6285 4641 6319 4675
rect 9873 4641 9907 4675
rect 9965 4641 9999 4675
rect 13185 4641 13219 4675
rect 14289 4641 14323 4675
rect 19993 4641 20027 4675
rect 21281 4641 21315 4675
rect 23857 4641 23891 4675
rect 24961 4641 24995 4675
rect 27629 4641 27663 4675
rect 28825 4641 28859 4675
rect 32873 4641 32907 4675
rect 38761 4641 38795 4675
rect 46213 4641 46247 4675
rect 50905 4641 50939 4675
rect 6929 4573 6963 4607
rect 8401 4573 8435 4607
rect 10057 4573 10091 4607
rect 10149 4573 10183 4607
rect 10701 4573 10735 4607
rect 11989 4573 12023 4607
rect 15393 4573 15427 4607
rect 17049 4573 17083 4607
rect 17509 4573 17543 4607
rect 18429 4573 18463 4607
rect 22385 4573 22419 4607
rect 23673 4573 23707 4607
rect 24685 4573 24719 4607
rect 26525 4573 26559 4607
rect 27813 4573 27847 4607
rect 28549 4573 28583 4607
rect 32689 4573 32723 4607
rect 32781 4573 32815 4607
rect 33609 4573 33643 4607
rect 33701 4573 33735 4607
rect 35725 4573 35759 4607
rect 37749 4573 37783 4607
rect 37841 4573 37875 4607
rect 38945 4573 38979 4607
rect 40049 4573 40083 4607
rect 41521 4573 41555 4607
rect 42717 4573 42751 4607
rect 42865 4573 42899 4607
rect 43085 4573 43119 4607
rect 43223 4573 43257 4607
rect 43913 4573 43947 4607
rect 44286 4573 44320 4607
rect 51089 4573 51123 4607
rect 58081 4573 58115 4607
rect 6101 4505 6135 4539
rect 7665 4505 7699 4539
rect 11805 4505 11839 4539
rect 12541 4505 12575 4539
rect 15669 4505 15703 4539
rect 17785 4505 17819 4539
rect 18705 4505 18739 4539
rect 21005 4505 21039 4539
rect 22661 4505 22695 4539
rect 30021 4505 30055 4539
rect 30205 4505 30239 4539
rect 34989 4505 35023 4539
rect 35173 4505 35207 4539
rect 35992 4505 36026 4539
rect 40877 4505 40911 4539
rect 42993 4505 43027 4539
rect 44097 4505 44131 4539
rect 44189 4505 44223 4539
rect 45293 4505 45327 4539
rect 46029 4505 46063 4539
rect 7757 4437 7791 4471
rect 12633 4437 12667 4471
rect 14749 4437 14783 4471
rect 19809 4437 19843 4471
rect 19901 4437 19935 4471
rect 20637 4437 20671 4471
rect 21097 4437 21131 4471
rect 23305 4437 23339 4471
rect 23765 4437 23799 4471
rect 26985 4437 27019 4471
rect 27997 4437 28031 4471
rect 33885 4437 33919 4471
rect 38025 4437 38059 4471
rect 40969 4437 41003 4471
rect 43361 4437 43395 4471
rect 51273 4437 51307 4471
rect 11069 4233 11103 4267
rect 11897 4233 11931 4267
rect 21189 4233 21223 4267
rect 24777 4233 24811 4267
rect 32689 4233 32723 4267
rect 37473 4233 37507 4267
rect 37933 4233 37967 4267
rect 53113 4233 53147 4267
rect 5825 4165 5859 4199
rect 6653 4165 6687 4199
rect 9965 4165 9999 4199
rect 10977 4165 11011 4199
rect 11805 4165 11839 4199
rect 12449 4165 12483 4199
rect 13369 4165 13403 4199
rect 14289 4165 14323 4199
rect 20076 4165 20110 4199
rect 26433 4165 26467 4199
rect 30757 4165 30791 4199
rect 31585 4165 31619 4199
rect 39957 4165 39991 4199
rect 40693 4165 40727 4199
rect 41429 4165 41463 4199
rect 44373 4165 44407 4199
rect 46581 4165 46615 4199
rect 52193 4165 52227 4199
rect 53021 4165 53055 4199
rect 53757 4165 53791 4199
rect 58173 4165 58207 4199
rect 1593 4097 1627 4131
rect 7389 4097 7423 4131
rect 8033 4097 8067 4131
rect 9229 4097 9263 4131
rect 17049 4097 17083 4131
rect 17969 4097 18003 4131
rect 18889 4097 18923 4131
rect 19809 4097 19843 4131
rect 22477 4097 22511 4131
rect 23397 4097 23431 4131
rect 23653 4097 23687 4131
rect 25237 4097 25271 4131
rect 27528 4097 27562 4131
rect 29101 4097 29135 4131
rect 29745 4097 29779 4131
rect 33517 4097 33551 4131
rect 34437 4097 34471 4131
rect 35357 4097 35391 4131
rect 36277 4097 36311 4131
rect 37841 4097 37875 4131
rect 38761 4097 38795 4131
rect 40877 4097 40911 4131
rect 41613 4097 41647 4131
rect 43269 4097 43303 4131
rect 43637 4097 43671 4131
rect 45109 4097 45143 4131
rect 45845 4097 45879 4131
rect 46029 4097 46063 4131
rect 46765 4097 46799 4131
rect 48237 4097 48271 4131
rect 53941 4097 53975 4131
rect 54585 4097 54619 4131
rect 1777 4029 1811 4063
rect 8953 4029 8987 4063
rect 9137 4029 9171 4063
rect 9321 4029 9355 4063
rect 9413 4029 9447 4063
rect 10425 4029 10459 4063
rect 12909 4029 12943 4063
rect 13829 4029 13863 4063
rect 14749 4029 14783 4063
rect 15485 4029 15519 4063
rect 17325 4029 17359 4063
rect 18245 4029 18279 4063
rect 19165 4029 19199 4063
rect 22753 4029 22787 4063
rect 25421 4029 25455 4063
rect 27261 4029 27295 4063
rect 29929 4029 29963 4063
rect 32781 4029 32815 4063
rect 32873 4029 32907 4063
rect 33701 4029 33735 4063
rect 34621 4029 34655 4063
rect 35541 4029 35575 4063
rect 36461 4029 36495 4063
rect 38117 4029 38151 4063
rect 39313 4029 39347 4063
rect 42625 4029 42659 4063
rect 43085 4029 43119 4063
rect 43545 4029 43579 4063
rect 58357 4029 58391 4063
rect 6009 3961 6043 3995
rect 6837 3961 6871 3995
rect 8401 3961 8435 3995
rect 8493 3961 8527 3995
rect 10241 3961 10275 3995
rect 12725 3961 12759 3995
rect 13645 3961 13679 3995
rect 14565 3961 14599 3995
rect 15761 3961 15795 3995
rect 31769 3961 31803 3995
rect 40141 3961 40175 3995
rect 48421 3961 48455 3995
rect 54769 3961 54803 3995
rect 7481 3893 7515 3927
rect 15945 3893 15979 3927
rect 28641 3893 28675 3927
rect 30849 3893 30883 3927
rect 32321 3893 32355 3927
rect 44465 3893 44499 3927
rect 45201 3893 45235 3927
rect 52285 3893 52319 3927
rect 10885 3689 10919 3723
rect 16221 3689 16255 3723
rect 24593 3689 24627 3723
rect 27813 3689 27847 3723
rect 33609 3689 33643 3723
rect 36553 3689 36587 3723
rect 45385 3689 45419 3723
rect 46121 3689 46155 3723
rect 47041 3689 47075 3723
rect 47961 3689 47995 3723
rect 48697 3689 48731 3723
rect 49433 3689 49467 3723
rect 50537 3689 50571 3723
rect 52009 3689 52043 3723
rect 54217 3689 54251 3723
rect 5273 3621 5307 3655
rect 6009 3621 6043 3655
rect 7573 3621 7607 3655
rect 8493 3621 8527 3655
rect 8585 3621 8619 3655
rect 10701 3621 10735 3655
rect 12081 3621 12115 3655
rect 13553 3621 13587 3655
rect 14565 3621 14599 3655
rect 16037 3621 16071 3655
rect 21097 3621 21131 3655
rect 38393 3621 38427 3655
rect 40417 3621 40451 3655
rect 42073 3621 42107 3655
rect 52837 3621 52871 3655
rect 55689 3621 55723 3655
rect 6745 3553 6779 3587
rect 9413 3553 9447 3587
rect 9689 3553 9723 3587
rect 13737 3553 13771 3587
rect 14749 3553 14783 3587
rect 15761 3553 15795 3587
rect 18613 3553 18647 3587
rect 18797 3553 18831 3587
rect 19717 3553 19751 3587
rect 25145 3553 25179 3587
rect 25973 3553 26007 3587
rect 28273 3553 28307 3587
rect 28457 3553 28491 3587
rect 32229 3553 32263 3587
rect 37013 3553 37047 3587
rect 37289 3553 37323 3587
rect 40877 3553 40911 3587
rect 42901 3553 42935 3587
rect 56885 3553 56919 3587
rect 1593 3485 1627 3519
rect 9597 3485 9631 3519
rect 9781 3485 9815 3519
rect 9873 3485 9907 3519
rect 12817 3485 12851 3519
rect 17233 3485 17267 3519
rect 18521 3485 18555 3519
rect 21741 3485 21775 3519
rect 22661 3485 22695 3519
rect 25789 3485 25823 3519
rect 27123 3485 27157 3519
rect 27353 3485 27387 3519
rect 30297 3485 30331 3519
rect 31401 3485 31435 3519
rect 31585 3485 31619 3519
rect 31769 3485 31803 3519
rect 32505 3485 32539 3519
rect 34897 3485 34931 3519
rect 35909 3485 35943 3519
rect 36057 3485 36091 3519
rect 36415 3485 36449 3519
rect 40785 3485 40819 3519
rect 41153 3485 41187 3519
rect 41245 3485 41279 3519
rect 43361 3485 43395 3519
rect 43637 3485 43671 3519
rect 43729 3485 43763 3519
rect 44005 3485 44039 3519
rect 44281 3485 44315 3519
rect 46029 3485 46063 3519
rect 48513 3485 48547 3519
rect 49249 3485 49283 3519
rect 51917 3485 51951 3519
rect 54125 3485 54159 3519
rect 55505 3485 55539 3519
rect 1869 3417 1903 3451
rect 5089 3417 5123 3451
rect 5825 3417 5859 3451
rect 6561 3417 6595 3451
rect 7205 3417 7239 3451
rect 8125 3417 8159 3451
rect 10425 3417 10459 3451
rect 11897 3417 11931 3451
rect 12633 3417 12667 3451
rect 13277 3417 13311 3451
rect 14289 3417 14323 3451
rect 17509 3417 17543 3451
rect 19962 3417 19996 3451
rect 22017 3417 22051 3451
rect 22928 3417 22962 3451
rect 24961 3417 24995 3451
rect 26801 3417 26835 3451
rect 26985 3417 27019 3451
rect 29009 3417 29043 3451
rect 30573 3417 30607 3451
rect 35173 3417 35207 3451
rect 36185 3417 36219 3451
rect 36277 3417 36311 3451
rect 39221 3417 39255 3451
rect 41889 3417 41923 3451
rect 45293 3417 45327 3451
rect 46949 3417 46983 3451
rect 47869 3417 47903 3451
rect 50445 3417 50479 3451
rect 51181 3417 51215 3451
rect 52653 3417 52687 3451
rect 53389 3417 53423 3451
rect 57130 3417 57164 3451
rect 7665 3349 7699 3383
rect 18153 3349 18187 3383
rect 24041 3349 24075 3383
rect 25053 3349 25087 3383
rect 27169 3349 27203 3383
rect 28181 3349 28215 3383
rect 39313 3349 39347 3383
rect 51273 3349 51307 3383
rect 53481 3349 53515 3383
rect 58265 3349 58299 3383
rect 8861 3145 8895 3179
rect 12541 3145 12575 3179
rect 13553 3145 13587 3179
rect 21097 3145 21131 3179
rect 23305 3145 23339 3179
rect 23673 3145 23707 3179
rect 34713 3145 34747 3179
rect 39773 3145 39807 3179
rect 40693 3145 40727 3179
rect 41797 3145 41831 3179
rect 44465 3145 44499 3179
rect 45201 3145 45235 3179
rect 47961 3145 47995 3179
rect 48881 3145 48915 3179
rect 49801 3145 49835 3179
rect 52193 3145 52227 3179
rect 54217 3145 54251 3179
rect 55321 3145 55355 3179
rect 57437 3145 57471 3179
rect 4353 3077 4387 3111
rect 6009 3077 6043 3111
rect 8401 3077 8435 3111
rect 23765 3077 23799 3111
rect 37933 3077 37967 3111
rect 42625 3077 42659 3111
rect 46765 3077 46799 3111
rect 50629 3077 50663 3111
rect 52101 3077 52135 3111
rect 56149 3077 56183 3111
rect 58173 3077 58207 3111
rect 1593 3009 1627 3043
rect 5089 3009 5123 3043
rect 5825 3009 5859 3043
rect 7021 3009 7055 3043
rect 7757 3009 7791 3043
rect 9505 3009 9539 3043
rect 9597 3009 9631 3043
rect 9781 3009 9815 3043
rect 12449 3009 12483 3043
rect 14013 3009 14047 3043
rect 14933 3009 14967 3043
rect 15853 3009 15887 3043
rect 16957 3009 16991 3043
rect 17877 3009 17911 3043
rect 18797 3009 18831 3043
rect 19717 3009 19751 3043
rect 19984 3009 20018 3043
rect 22385 3009 22419 3043
rect 25237 3009 25271 3043
rect 26157 3009 26191 3043
rect 27537 3009 27571 3043
rect 28457 3009 28491 3043
rect 28733 3009 28767 3043
rect 30849 3009 30883 3043
rect 32321 3009 32355 3043
rect 33333 3009 33367 3043
rect 35449 3009 35483 3043
rect 36369 3009 36403 3043
rect 37565 3009 37599 3043
rect 38669 3009 38703 3043
rect 39681 3009 39715 3043
rect 40601 3009 40635 3043
rect 41705 3009 41739 3043
rect 43269 3009 43303 3043
rect 43637 3009 43671 3043
rect 44373 3009 44407 3043
rect 45017 3009 45051 3043
rect 46397 3009 46431 3043
rect 47869 3009 47903 3043
rect 48789 3009 48823 3043
rect 49709 3009 49743 3043
rect 51365 3009 51399 3043
rect 53021 3009 53055 3043
rect 54125 3009 54159 3043
rect 55045 3009 55079 3043
rect 55873 3009 55907 3043
rect 57253 3009 57287 3043
rect 1777 2941 1811 2975
rect 9321 2941 9355 2975
rect 9689 2941 9723 2975
rect 10333 2941 10367 2975
rect 13093 2941 13127 2975
rect 14289 2941 14323 2975
rect 15209 2941 15243 2975
rect 16129 2941 16163 2975
rect 17233 2941 17267 2975
rect 18153 2941 18187 2975
rect 18981 2941 19015 2975
rect 22661 2941 22695 2975
rect 23949 2941 23983 2975
rect 25421 2941 25455 2975
rect 26433 2941 26467 2975
rect 27813 2941 27847 2975
rect 31033 2941 31067 2975
rect 32505 2941 32539 2975
rect 33609 2941 33643 2975
rect 35633 2941 35667 2975
rect 36553 2941 36587 2975
rect 38945 2941 38979 2975
rect 43361 2941 43395 2975
rect 43545 2941 43579 2975
rect 53205 2941 53239 2975
rect 57069 2941 57103 2975
rect 58357 2941 58391 2975
rect 5273 2873 5307 2907
rect 8677 2873 8711 2907
rect 10609 2873 10643 2907
rect 10793 2873 10827 2907
rect 13369 2873 13403 2907
rect 29837 2873 29871 2907
rect 50813 2873 50847 2907
rect 51549 2873 51583 2907
rect 4445 2805 4479 2839
rect 7113 2805 7147 2839
rect 7849 2805 7883 2839
rect 24777 2805 24811 2839
rect 3341 2601 3375 2635
rect 8493 2601 8527 2635
rect 14473 2601 14507 2635
rect 19993 2601 20027 2635
rect 22201 2601 22235 2635
rect 43085 2601 43119 2635
rect 45385 2601 45419 2635
rect 46213 2601 46247 2635
rect 47961 2601 47995 2635
rect 48881 2601 48915 2635
rect 52009 2601 52043 2635
rect 58265 2601 58299 2635
rect 6009 2533 6043 2567
rect 10425 2533 10459 2567
rect 11161 2533 11195 2567
rect 41245 2533 41279 2567
rect 4537 2465 4571 2499
rect 12633 2465 12667 2499
rect 17049 2465 17083 2499
rect 20453 2465 20487 2499
rect 20637 2465 20671 2499
rect 24593 2465 24627 2499
rect 54033 2465 54067 2499
rect 55689 2465 55723 2499
rect 1593 2397 1627 2431
rect 4353 2397 4387 2431
rect 8401 2397 8435 2431
rect 10241 2397 10275 2431
rect 12357 2397 12391 2431
rect 13277 2397 13311 2431
rect 14933 2397 14967 2431
rect 15853 2397 15887 2431
rect 17509 2397 17543 2431
rect 18429 2397 18463 2431
rect 20361 2397 20395 2431
rect 21281 2397 21315 2431
rect 22661 2397 22695 2431
rect 23581 2397 23615 2431
rect 25237 2397 25271 2431
rect 26157 2397 26191 2431
rect 27813 2397 27847 2431
rect 28733 2397 28767 2431
rect 30205 2397 30239 2431
rect 31125 2397 31159 2431
rect 32321 2397 32355 2431
rect 33241 2397 33275 2431
rect 34897 2397 34931 2431
rect 35817 2397 35851 2431
rect 37473 2397 37507 2431
rect 38393 2397 38427 2431
rect 40049 2397 40083 2431
rect 43269 2397 43303 2431
rect 43453 2397 43487 2431
rect 43821 2397 43855 2431
rect 43913 2397 43947 2431
rect 51365 2397 51399 2431
rect 53849 2397 53883 2431
rect 55505 2397 55539 2431
rect 57069 2397 57103 2431
rect 58173 2397 58207 2431
rect 1869 2329 1903 2363
rect 3249 2329 3283 2363
rect 5089 2329 5123 2363
rect 5825 2329 5859 2363
rect 6929 2329 6963 2363
rect 7113 2329 7147 2363
rect 7665 2329 7699 2363
rect 9505 2329 9539 2363
rect 9689 2329 9723 2363
rect 10977 2329 11011 2363
rect 13553 2329 13587 2363
rect 15209 2329 15243 2363
rect 16129 2329 16163 2363
rect 17785 2329 17819 2363
rect 18705 2329 18739 2363
rect 22937 2329 22971 2363
rect 23857 2329 23891 2363
rect 25513 2329 25547 2363
rect 26433 2329 26467 2363
rect 28089 2329 28123 2363
rect 29009 2329 29043 2363
rect 30481 2329 30515 2363
rect 31401 2329 31435 2363
rect 32597 2329 32631 2363
rect 33517 2329 33551 2363
rect 35173 2329 35207 2363
rect 36093 2329 36127 2363
rect 37749 2329 37783 2363
rect 38669 2329 38703 2363
rect 40325 2329 40359 2363
rect 41061 2329 41095 2363
rect 45293 2329 45327 2363
rect 46121 2329 46155 2363
rect 47041 2329 47075 2363
rect 47869 2329 47903 2363
rect 48789 2329 48823 2363
rect 50445 2329 50479 2363
rect 51181 2329 51215 2363
rect 51917 2329 51951 2363
rect 53021 2329 53055 2363
rect 57345 2329 57379 2363
rect 5181 2261 5215 2295
rect 7757 2261 7791 2295
rect 21373 2261 21407 2295
rect 27169 2261 27203 2295
rect 47133 2261 47167 2295
rect 50537 2261 50571 2295
rect 53113 2261 53147 2295
<< metal1 >>
rect 30190 63248 30196 63300
rect 30248 63288 30254 63300
rect 30466 63288 30472 63300
rect 30248 63260 30472 63288
rect 30248 63248 30254 63260
rect 30466 63248 30472 63260
rect 30524 63248 30530 63300
rect 32582 63248 32588 63300
rect 32640 63288 32646 63300
rect 33318 63288 33324 63300
rect 32640 63260 33324 63288
rect 32640 63248 32646 63260
rect 33318 63248 33324 63260
rect 33376 63248 33382 63300
rect 34054 63248 34060 63300
rect 34112 63288 34118 63300
rect 34790 63288 34796 63300
rect 34112 63260 34796 63288
rect 34112 63248 34118 63260
rect 34790 63248 34796 63260
rect 34848 63248 34854 63300
rect 39206 63248 39212 63300
rect 39264 63288 39270 63300
rect 40126 63288 40132 63300
rect 39264 63260 40132 63288
rect 39264 63248 39270 63260
rect 40126 63248 40132 63260
rect 40184 63248 40190 63300
rect 40678 63248 40684 63300
rect 40736 63288 40742 63300
rect 41598 63288 41604 63300
rect 40736 63260 41604 63288
rect 40736 63248 40742 63260
rect 41598 63248 41604 63260
rect 41656 63248 41662 63300
rect 43530 63112 43536 63164
rect 43588 63152 43594 63164
rect 44358 63152 44364 63164
rect 43588 63124 44364 63152
rect 43588 63112 43594 63124
rect 44358 63112 44364 63124
rect 44416 63112 44422 63164
rect 30282 61684 30288 61736
rect 30340 61724 30346 61736
rect 49418 61724 49424 61736
rect 30340 61696 49424 61724
rect 30340 61684 30346 61696
rect 49418 61684 49424 61696
rect 49476 61684 49482 61736
rect 9766 61616 9772 61668
rect 9824 61656 9830 61668
rect 23474 61656 23480 61668
rect 9824 61628 23480 61656
rect 9824 61616 9830 61628
rect 23474 61616 23480 61628
rect 23532 61616 23538 61668
rect 33502 61616 33508 61668
rect 33560 61656 33566 61668
rect 41782 61656 41788 61668
rect 33560 61628 41788 61656
rect 33560 61616 33566 61628
rect 41782 61616 41788 61628
rect 41840 61616 41846 61668
rect 5166 61548 5172 61600
rect 5224 61588 5230 61600
rect 17862 61588 17868 61600
rect 5224 61560 17868 61588
rect 5224 61548 5230 61560
rect 17862 61548 17868 61560
rect 17920 61548 17926 61600
rect 28902 61548 28908 61600
rect 28960 61588 28966 61600
rect 46842 61588 46848 61600
rect 28960 61560 46848 61588
rect 28960 61548 28966 61560
rect 46842 61548 46848 61560
rect 46900 61548 46906 61600
rect 1104 61498 58880 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 58880 61498
rect 1104 61424 58880 61446
rect 5166 61344 5172 61396
rect 5224 61344 5230 61396
rect 8202 61344 8208 61396
rect 8260 61384 8266 61396
rect 35986 61384 35992 61396
rect 8260 61356 35992 61384
rect 8260 61344 8266 61356
rect 35986 61344 35992 61356
rect 36044 61344 36050 61396
rect 36170 61344 36176 61396
rect 36228 61384 36234 61396
rect 44453 61387 44511 61393
rect 44453 61384 44465 61387
rect 36228 61356 44465 61384
rect 36228 61344 36234 61356
rect 44453 61353 44465 61356
rect 44499 61353 44511 61387
rect 44453 61347 44511 61353
rect 46842 61344 46848 61396
rect 46900 61344 46906 61396
rect 49418 61344 49424 61396
rect 49476 61344 49482 61396
rect 9677 61319 9735 61325
rect 9677 61285 9689 61319
rect 9723 61316 9735 61319
rect 9766 61316 9772 61328
rect 9723 61288 9772 61316
rect 9723 61285 9735 61288
rect 9677 61279 9735 61285
rect 9766 61276 9772 61288
rect 9824 61276 9830 61328
rect 11149 61319 11207 61325
rect 11149 61285 11161 61319
rect 11195 61316 11207 61319
rect 19334 61316 19340 61328
rect 11195 61288 19340 61316
rect 11195 61285 11207 61288
rect 11149 61279 11207 61285
rect 19334 61276 19340 61288
rect 19392 61276 19398 61328
rect 20717 61319 20775 61325
rect 20717 61285 20729 61319
rect 20763 61316 20775 61319
rect 22094 61316 22100 61328
rect 20763 61288 22100 61316
rect 20763 61285 20775 61288
rect 20717 61279 20775 61285
rect 22094 61276 22100 61288
rect 22152 61276 22158 61328
rect 22649 61319 22707 61325
rect 22649 61285 22661 61319
rect 22695 61316 22707 61319
rect 26878 61316 26884 61328
rect 22695 61288 26884 61316
rect 22695 61285 22707 61288
rect 22649 61279 22707 61285
rect 26878 61276 26884 61288
rect 26936 61276 26942 61328
rect 38473 61319 38531 61325
rect 38473 61316 38485 61319
rect 31036 61288 38485 61316
rect 2225 61251 2283 61257
rect 2225 61217 2237 61251
rect 2271 61248 2283 61251
rect 7650 61248 7656 61260
rect 2271 61220 7656 61248
rect 2271 61217 2283 61220
rect 2225 61211 2283 61217
rect 7650 61208 7656 61220
rect 7708 61208 7714 61260
rect 10413 61251 10471 61257
rect 10413 61217 10425 61251
rect 10459 61248 10471 61251
rect 18046 61248 18052 61260
rect 10459 61220 18052 61248
rect 10459 61217 10471 61220
rect 10413 61211 10471 61217
rect 18046 61208 18052 61220
rect 18104 61208 18110 61260
rect 18141 61251 18199 61257
rect 18141 61217 18153 61251
rect 18187 61248 18199 61251
rect 23014 61248 23020 61260
rect 18187 61220 23020 61248
rect 18187 61217 18199 61220
rect 18141 61211 18199 61217
rect 23014 61208 23020 61220
rect 23072 61208 23078 61260
rect 31036 61248 31064 61288
rect 38473 61285 38485 61288
rect 38519 61285 38531 61319
rect 38473 61279 38531 61285
rect 43717 61319 43775 61325
rect 43717 61285 43729 61319
rect 43763 61285 43775 61319
rect 43717 61279 43775 61285
rect 23584 61220 31064 61248
rect 934 61140 940 61192
rect 992 61180 998 61192
rect 1673 61183 1731 61189
rect 1673 61180 1685 61183
rect 992 61152 1685 61180
rect 992 61140 998 61152
rect 1673 61149 1685 61152
rect 1719 61149 1731 61183
rect 2777 61183 2835 61189
rect 2777 61180 2789 61183
rect 1673 61143 1731 61149
rect 1780 61152 2789 61180
rect 1026 61072 1032 61124
rect 1084 61112 1090 61124
rect 1780 61112 1808 61152
rect 2777 61149 2789 61152
rect 2823 61149 2835 61183
rect 2777 61143 2835 61149
rect 4341 61183 4399 61189
rect 4341 61149 4353 61183
rect 4387 61180 4399 61183
rect 4614 61180 4620 61192
rect 4387 61152 4620 61180
rect 4387 61149 4399 61152
rect 4341 61143 4399 61149
rect 4614 61140 4620 61152
rect 4672 61140 4678 61192
rect 5074 61140 5080 61192
rect 5132 61140 5138 61192
rect 5718 61140 5724 61192
rect 5776 61140 5782 61192
rect 6638 61140 6644 61192
rect 6696 61140 6702 61192
rect 7558 61140 7564 61192
rect 7616 61140 7622 61192
rect 9493 61183 9551 61189
rect 9493 61149 9505 61183
rect 9539 61180 9551 61183
rect 9674 61180 9680 61192
rect 9539 61152 9680 61180
rect 9539 61149 9551 61152
rect 9493 61143 9551 61149
rect 9674 61140 9680 61152
rect 9732 61140 9738 61192
rect 10226 61140 10232 61192
rect 10284 61140 10290 61192
rect 10965 61183 11023 61189
rect 10965 61149 10977 61183
rect 11011 61180 11023 61183
rect 11146 61180 11152 61192
rect 11011 61152 11152 61180
rect 11011 61149 11023 61152
rect 10965 61143 11023 61149
rect 11146 61140 11152 61152
rect 11204 61140 11210 61192
rect 11974 61140 11980 61192
rect 12032 61140 12038 61192
rect 12710 61140 12716 61192
rect 12768 61140 12774 61192
rect 14918 61140 14924 61192
rect 14976 61140 14982 61192
rect 16114 61140 16120 61192
rect 16172 61140 16178 61192
rect 17126 61140 17132 61192
rect 17184 61140 17190 61192
rect 17954 61140 17960 61192
rect 18012 61140 18018 61192
rect 18690 61140 18696 61192
rect 18748 61140 18754 61192
rect 19794 61140 19800 61192
rect 19852 61140 19858 61192
rect 20533 61183 20591 61189
rect 20533 61149 20545 61183
rect 20579 61180 20591 61183
rect 20714 61180 20720 61192
rect 20579 61152 20720 61180
rect 20579 61149 20591 61152
rect 20533 61143 20591 61149
rect 20714 61140 20720 61152
rect 20772 61140 20778 61192
rect 21266 61140 21272 61192
rect 21324 61140 21330 61192
rect 22186 61140 22192 61192
rect 22244 61180 22250 61192
rect 22373 61183 22431 61189
rect 22373 61180 22385 61183
rect 22244 61152 22385 61180
rect 22244 61140 22250 61152
rect 22373 61149 22385 61152
rect 22419 61149 22431 61183
rect 22373 61143 22431 61149
rect 1084 61084 1808 61112
rect 3053 61115 3111 61121
rect 1084 61072 1090 61084
rect 3053 61081 3065 61115
rect 3099 61081 3111 61115
rect 3053 61075 3111 61081
rect 4525 61115 4583 61121
rect 4525 61081 4537 61115
rect 4571 61112 4583 61115
rect 5626 61112 5632 61124
rect 4571 61084 5632 61112
rect 4571 61081 4583 61084
rect 4525 61075 4583 61081
rect 3068 61044 3096 61075
rect 5626 61072 5632 61084
rect 5684 61072 5690 61124
rect 6178 61112 6184 61124
rect 5828 61084 6184 61112
rect 5828 61044 5856 61084
rect 6178 61072 6184 61084
rect 6236 61072 6242 61124
rect 6914 61072 6920 61124
rect 6972 61072 6978 61124
rect 7837 61115 7895 61121
rect 7837 61081 7849 61115
rect 7883 61112 7895 61115
rect 9122 61112 9128 61124
rect 7883 61084 9128 61112
rect 7883 61081 7895 61084
rect 7837 61075 7895 61081
rect 9122 61072 9128 61084
rect 9180 61072 9186 61124
rect 12989 61115 13047 61121
rect 12989 61081 13001 61115
rect 13035 61112 13047 61115
rect 13630 61112 13636 61124
rect 13035 61084 13636 61112
rect 13035 61081 13047 61084
rect 12989 61075 13047 61081
rect 13630 61072 13636 61084
rect 13688 61072 13694 61124
rect 15194 61072 15200 61124
rect 15252 61072 15258 61124
rect 16301 61115 16359 61121
rect 16301 61081 16313 61115
rect 16347 61112 16359 61115
rect 17494 61112 17500 61124
rect 16347 61084 17500 61112
rect 16347 61081 16359 61084
rect 16301 61075 16359 61081
rect 17494 61072 17500 61084
rect 17552 61072 17558 61124
rect 19978 61072 19984 61124
rect 20036 61072 20042 61124
rect 21174 61072 21180 61124
rect 21232 61112 21238 61124
rect 23584 61112 23612 61220
rect 32950 61208 32956 61260
rect 33008 61248 33014 61260
rect 35161 61251 35219 61257
rect 35161 61248 35173 61251
rect 33008 61220 35173 61248
rect 33008 61208 33014 61220
rect 35161 61217 35173 61220
rect 35207 61217 35219 61251
rect 35161 61211 35219 61217
rect 35894 61208 35900 61260
rect 35952 61248 35958 61260
rect 43732 61248 43760 61279
rect 48041 61251 48099 61257
rect 48041 61248 48053 61251
rect 35952 61220 36492 61248
rect 35952 61208 35958 61220
rect 23658 61140 23664 61192
rect 23716 61180 23722 61192
rect 23845 61183 23903 61189
rect 23845 61180 23857 61183
rect 23716 61152 23857 61180
rect 23716 61140 23722 61152
rect 23845 61149 23857 61152
rect 23891 61149 23903 61183
rect 23845 61143 23903 61149
rect 25130 61140 25136 61192
rect 25188 61180 25194 61192
rect 25317 61183 25375 61189
rect 25317 61180 25329 61183
rect 25188 61152 25329 61180
rect 25188 61140 25194 61152
rect 25317 61149 25329 61152
rect 25363 61149 25375 61183
rect 25317 61143 25375 61149
rect 26234 61140 26240 61192
rect 26292 61140 26298 61192
rect 26602 61140 26608 61192
rect 26660 61180 26666 61192
rect 27249 61183 27307 61189
rect 27249 61180 27261 61183
rect 26660 61152 27261 61180
rect 26660 61140 26666 61152
rect 27249 61149 27261 61152
rect 27295 61149 27307 61183
rect 27249 61143 27307 61149
rect 28074 61140 28080 61192
rect 28132 61180 28138 61192
rect 28261 61183 28319 61189
rect 28261 61180 28273 61183
rect 28132 61152 28273 61180
rect 28132 61140 28138 61152
rect 28261 61149 28273 61152
rect 28307 61149 28319 61183
rect 28261 61143 28319 61149
rect 29822 61140 29828 61192
rect 29880 61140 29886 61192
rect 31202 61140 31208 61192
rect 31260 61140 31266 61192
rect 31754 61140 31760 61192
rect 31812 61180 31818 61192
rect 32401 61183 32459 61189
rect 32401 61180 32413 61183
rect 31812 61152 32413 61180
rect 31812 61140 31818 61152
rect 32401 61149 32413 61152
rect 32447 61149 32459 61183
rect 32401 61143 32459 61149
rect 33318 61140 33324 61192
rect 33376 61140 33382 61192
rect 33502 61140 33508 61192
rect 33560 61140 33566 61192
rect 34790 61140 34796 61192
rect 34848 61180 34854 61192
rect 36464 61189 36492 61220
rect 37200 61220 43760 61248
rect 43824 61220 48053 61248
rect 34977 61183 35035 61189
rect 34977 61180 34989 61183
rect 34848 61152 34989 61180
rect 34848 61140 34854 61152
rect 34977 61149 34989 61152
rect 35023 61149 35035 61183
rect 34977 61143 35035 61149
rect 36449 61183 36507 61189
rect 36449 61149 36461 61183
rect 36495 61149 36507 61183
rect 36449 61143 36507 61149
rect 21232 61084 23612 61112
rect 24029 61115 24087 61121
rect 21232 61072 21238 61084
rect 24029 61081 24041 61115
rect 24075 61112 24087 61115
rect 24762 61112 24768 61124
rect 24075 61084 24768 61112
rect 24075 61081 24087 61084
rect 24029 61075 24087 61081
rect 24762 61072 24768 61084
rect 24820 61072 24826 61124
rect 26421 61115 26479 61121
rect 26421 61081 26433 61115
rect 26467 61112 26479 61115
rect 28166 61112 28172 61124
rect 26467 61084 28172 61112
rect 26467 61081 26479 61084
rect 26421 61075 26479 61081
rect 28166 61072 28172 61084
rect 28224 61072 28230 61124
rect 33226 61072 33232 61124
rect 33284 61112 33290 61124
rect 34057 61115 34115 61121
rect 34057 61112 34069 61115
rect 33284 61084 34069 61112
rect 33284 61072 33290 61084
rect 34057 61081 34069 61084
rect 34103 61081 34115 61115
rect 34057 61075 34115 61081
rect 34698 61072 34704 61124
rect 34756 61112 34762 61124
rect 35713 61115 35771 61121
rect 35713 61112 35725 61115
rect 34756 61084 35725 61112
rect 34756 61072 34762 61084
rect 35713 61081 35725 61084
rect 35759 61081 35771 61115
rect 35713 61075 35771 61081
rect 35894 61072 35900 61124
rect 35952 61072 35958 61124
rect 35986 61072 35992 61124
rect 36044 61112 36050 61124
rect 37200 61112 37228 61220
rect 37274 61140 37280 61192
rect 37332 61180 37338 61192
rect 37553 61183 37611 61189
rect 37553 61180 37565 61183
rect 37332 61152 37565 61180
rect 37332 61140 37338 61152
rect 37553 61149 37565 61152
rect 37599 61149 37611 61183
rect 37553 61143 37611 61149
rect 37642 61140 37648 61192
rect 37700 61180 37706 61192
rect 38289 61183 38347 61189
rect 38289 61180 38301 61183
rect 37700 61152 38301 61180
rect 37700 61140 37706 61152
rect 38289 61149 38301 61152
rect 38335 61149 38347 61183
rect 38289 61143 38347 61149
rect 38746 61140 38752 61192
rect 38804 61180 38810 61192
rect 38933 61183 38991 61189
rect 38933 61180 38945 61183
rect 38804 61152 38945 61180
rect 38804 61140 38810 61152
rect 38933 61149 38945 61152
rect 38979 61149 38991 61183
rect 38933 61143 38991 61149
rect 40126 61140 40132 61192
rect 40184 61140 40190 61192
rect 41598 61140 41604 61192
rect 41656 61140 41662 61192
rect 42058 61140 42064 61192
rect 42116 61180 42122 61192
rect 42613 61183 42671 61189
rect 42613 61180 42625 61183
rect 42116 61152 42625 61180
rect 42116 61140 42122 61152
rect 42613 61149 42625 61152
rect 42659 61149 42671 61183
rect 42613 61143 42671 61149
rect 42794 61140 42800 61192
rect 42852 61180 42858 61192
rect 43533 61183 43591 61189
rect 43533 61180 43545 61183
rect 42852 61152 43545 61180
rect 42852 61140 42858 61152
rect 43533 61149 43545 61152
rect 43579 61149 43591 61183
rect 43533 61143 43591 61149
rect 36044 61084 37228 61112
rect 37737 61115 37795 61121
rect 36044 61072 36050 61084
rect 37737 61081 37749 61115
rect 37783 61112 37795 61115
rect 38194 61112 38200 61124
rect 37783 61084 38200 61112
rect 37783 61081 37795 61084
rect 37737 61075 37795 61081
rect 38194 61072 38200 61084
rect 38252 61072 38258 61124
rect 40034 61072 40040 61124
rect 40092 61112 40098 61124
rect 40865 61115 40923 61121
rect 40865 61112 40877 61115
rect 40092 61084 40877 61112
rect 40092 61072 40098 61084
rect 40865 61081 40877 61084
rect 40911 61081 40923 61115
rect 40865 61075 40923 61081
rect 41414 61072 41420 61124
rect 41472 61112 41478 61124
rect 42889 61115 42947 61121
rect 41472 61084 41828 61112
rect 41472 61072 41478 61084
rect 3068 61016 5856 61044
rect 5902 61004 5908 61056
rect 5960 61004 5966 61056
rect 12158 61004 12164 61056
rect 12216 61004 12222 61056
rect 17310 61004 17316 61056
rect 17368 61004 17374 61056
rect 18782 61004 18788 61056
rect 18840 61004 18846 61056
rect 20990 61004 20996 61056
rect 21048 61044 21054 61056
rect 21361 61047 21419 61053
rect 21361 61044 21373 61047
rect 21048 61016 21373 61044
rect 21048 61004 21054 61016
rect 21361 61013 21373 61016
rect 21407 61013 21419 61047
rect 21361 61007 21419 61013
rect 22002 61004 22008 61056
rect 22060 61044 22066 61056
rect 24670 61044 24676 61056
rect 22060 61016 24676 61044
rect 22060 61004 22066 61016
rect 24670 61004 24676 61016
rect 24728 61004 24734 61056
rect 25406 61004 25412 61056
rect 25464 61004 25470 61056
rect 27338 61004 27344 61056
rect 27396 61004 27402 61056
rect 28353 61047 28411 61053
rect 28353 61013 28365 61047
rect 28399 61044 28411 61047
rect 28442 61044 28448 61056
rect 28399 61016 28448 61044
rect 28399 61013 28411 61016
rect 28353 61007 28411 61013
rect 28442 61004 28448 61016
rect 28500 61004 28506 61056
rect 29914 61004 29920 61056
rect 29972 61004 29978 61056
rect 31294 61004 31300 61056
rect 31352 61004 31358 61056
rect 32493 61047 32551 61053
rect 32493 61013 32505 61047
rect 32539 61044 32551 61047
rect 32582 61044 32588 61056
rect 32539 61016 32588 61044
rect 32539 61013 32551 61016
rect 32493 61007 32551 61013
rect 32582 61004 32588 61016
rect 32640 61004 32646 61056
rect 33502 61004 33508 61056
rect 33560 61044 33566 61056
rect 34149 61047 34207 61053
rect 34149 61044 34161 61047
rect 33560 61016 34161 61044
rect 33560 61004 33566 61016
rect 34149 61013 34161 61016
rect 34195 61013 34207 61047
rect 34149 61007 34207 61013
rect 36078 61004 36084 61056
rect 36136 61044 36142 61056
rect 36541 61047 36599 61053
rect 36541 61044 36553 61047
rect 36136 61016 36553 61044
rect 36136 61004 36142 61016
rect 36541 61013 36553 61016
rect 36587 61013 36599 61047
rect 36541 61007 36599 61013
rect 39114 61004 39120 61056
rect 39172 61004 39178 61056
rect 40218 61004 40224 61056
rect 40276 61004 40282 61056
rect 40310 61004 40316 61056
rect 40368 61044 40374 61056
rect 40957 61047 41015 61053
rect 40957 61044 40969 61047
rect 40368 61016 40969 61044
rect 40368 61004 40374 61016
rect 40957 61013 40969 61016
rect 41003 61013 41015 61047
rect 40957 61007 41015 61013
rect 41690 61004 41696 61056
rect 41748 61004 41754 61056
rect 41800 61044 41828 61084
rect 42889 61081 42901 61115
rect 42935 61112 42947 61115
rect 42978 61112 42984 61124
rect 42935 61084 42984 61112
rect 42935 61081 42947 61084
rect 42889 61075 42947 61081
rect 42978 61072 42984 61084
rect 43036 61072 43042 61124
rect 43824 61044 43852 61220
rect 48041 61217 48053 61220
rect 48087 61217 48099 61251
rect 48041 61211 48099 61217
rect 56686 61208 56692 61260
rect 56744 61248 56750 61260
rect 58986 61248 58992 61260
rect 56744 61220 58992 61248
rect 56744 61208 56750 61220
rect 58986 61208 58992 61220
rect 59044 61208 59050 61260
rect 44358 61140 44364 61192
rect 44416 61140 44422 61192
rect 44542 61140 44548 61192
rect 44600 61180 44606 61192
rect 45281 61183 45339 61189
rect 45281 61180 45293 61183
rect 44600 61152 45293 61180
rect 44600 61140 44606 61152
rect 45281 61149 45293 61152
rect 45327 61149 45339 61183
rect 45281 61143 45339 61149
rect 45554 61140 45560 61192
rect 45612 61180 45618 61192
rect 45612 61152 45692 61180
rect 45612 61140 45618 61152
rect 44818 61072 44824 61124
rect 44876 61112 44882 61124
rect 45664 61112 45692 61152
rect 45738 61140 45744 61192
rect 45796 61180 45802 61192
rect 46753 61183 46811 61189
rect 46753 61180 46765 61183
rect 45796 61152 46765 61180
rect 45796 61140 45802 61152
rect 46753 61149 46765 61152
rect 46799 61149 46811 61183
rect 46753 61143 46811 61149
rect 47210 61140 47216 61192
rect 47268 61180 47274 61192
rect 47857 61183 47915 61189
rect 47857 61180 47869 61183
rect 47268 61152 47869 61180
rect 47268 61140 47274 61152
rect 47857 61149 47869 61152
rect 47903 61149 47915 61183
rect 47857 61143 47915 61149
rect 48314 61140 48320 61192
rect 48372 61180 48378 61192
rect 48593 61183 48651 61189
rect 48593 61180 48605 61183
rect 48372 61152 48605 61180
rect 48372 61140 48378 61152
rect 48593 61149 48605 61152
rect 48639 61149 48651 61183
rect 48593 61143 48651 61149
rect 48682 61140 48688 61192
rect 48740 61180 48746 61192
rect 49329 61183 49387 61189
rect 49329 61180 49341 61183
rect 48740 61152 49341 61180
rect 48740 61140 48746 61152
rect 49329 61149 49341 61152
rect 49375 61149 49387 61183
rect 49329 61143 49387 61149
rect 49786 61140 49792 61192
rect 49844 61180 49850 61192
rect 50433 61183 50491 61189
rect 50433 61180 50445 61183
rect 49844 61152 50445 61180
rect 49844 61140 49850 61152
rect 50433 61149 50445 61152
rect 50479 61149 50491 61183
rect 50433 61143 50491 61149
rect 51258 61140 51264 61192
rect 51316 61180 51322 61192
rect 51353 61183 51411 61189
rect 51353 61180 51365 61183
rect 51316 61152 51365 61180
rect 51316 61140 51322 61152
rect 51353 61149 51365 61152
rect 51399 61149 51411 61183
rect 51353 61143 51411 61149
rect 51626 61140 51632 61192
rect 51684 61180 51690 61192
rect 52089 61183 52147 61189
rect 52089 61180 52101 61183
rect 51684 61152 52101 61180
rect 51684 61140 51690 61152
rect 52089 61149 52101 61152
rect 52135 61149 52147 61183
rect 52089 61143 52147 61149
rect 53190 61140 53196 61192
rect 53248 61140 53254 61192
rect 54110 61140 54116 61192
rect 54168 61140 54174 61192
rect 55490 61140 55496 61192
rect 55548 61140 55554 61192
rect 56042 61140 56048 61192
rect 56100 61180 56106 61192
rect 56505 61183 56563 61189
rect 56505 61180 56517 61183
rect 56100 61152 56517 61180
rect 56100 61140 56106 61152
rect 56505 61149 56517 61152
rect 56551 61149 56563 61183
rect 56505 61143 56563 61149
rect 57514 61140 57520 61192
rect 57572 61180 57578 61192
rect 58161 61183 58219 61189
rect 58161 61180 58173 61183
rect 57572 61152 58173 61180
rect 57572 61140 57578 61152
rect 58161 61149 58173 61152
rect 58207 61149 58219 61183
rect 58161 61143 58219 61149
rect 46017 61115 46075 61121
rect 46017 61112 46029 61115
rect 44876 61084 45554 61112
rect 45664 61084 46029 61112
rect 44876 61072 44882 61084
rect 41800 61016 43852 61044
rect 45370 61004 45376 61056
rect 45428 61004 45434 61056
rect 45526 61044 45554 61084
rect 46017 61081 46029 61084
rect 46063 61081 46075 61115
rect 46017 61075 46075 61081
rect 49694 61072 49700 61124
rect 49752 61112 49758 61124
rect 52273 61115 52331 61121
rect 52273 61112 52285 61115
rect 49752 61084 52285 61112
rect 49752 61072 49758 61084
rect 52273 61081 52285 61084
rect 52319 61081 52331 61115
rect 52273 61075 52331 61081
rect 53466 61072 53472 61124
rect 53524 61072 53530 61124
rect 55766 61072 55772 61124
rect 55824 61072 55830 61124
rect 58342 61072 58348 61124
rect 58400 61072 58406 61124
rect 46109 61047 46167 61053
rect 46109 61044 46121 61047
rect 45526 61016 46121 61044
rect 46109 61013 46121 61016
rect 46155 61013 46167 61047
rect 46109 61007 46167 61013
rect 46842 61004 46848 61056
rect 46900 61044 46906 61056
rect 48685 61047 48743 61053
rect 48685 61044 48697 61047
rect 46900 61016 48697 61044
rect 46900 61004 46906 61016
rect 48685 61013 48697 61016
rect 48731 61013 48743 61047
rect 48685 61007 48743 61013
rect 50062 61004 50068 61056
rect 50120 61044 50126 61056
rect 50525 61047 50583 61053
rect 50525 61044 50537 61047
rect 50120 61016 50537 61044
rect 50120 61004 50126 61016
rect 50525 61013 50537 61016
rect 50571 61013 50583 61047
rect 50525 61007 50583 61013
rect 50614 61004 50620 61056
rect 50672 61044 50678 61056
rect 51445 61047 51503 61053
rect 51445 61044 51457 61047
rect 50672 61016 51457 61044
rect 50672 61004 50678 61016
rect 51445 61013 51457 61016
rect 51491 61013 51503 61047
rect 51445 61007 51503 61013
rect 54294 61004 54300 61056
rect 54352 61004 54358 61056
rect 56594 61004 56600 61056
rect 56652 61004 56658 61056
rect 1104 60954 58880 60976
rect 1104 60902 19574 60954
rect 19626 60902 19638 60954
rect 19690 60902 19702 60954
rect 19754 60902 19766 60954
rect 19818 60902 19830 60954
rect 19882 60902 50294 60954
rect 50346 60902 50358 60954
rect 50410 60902 50422 60954
rect 50474 60902 50486 60954
rect 50538 60902 50550 60954
rect 50602 60902 58880 60954
rect 1104 60880 58880 60902
rect 36170 60840 36176 60852
rect 23492 60812 36176 60840
rect 3234 60732 3240 60784
rect 3292 60732 3298 60784
rect 3970 60732 3976 60784
rect 4028 60732 4034 60784
rect 8386 60732 8392 60784
rect 8444 60732 8450 60784
rect 13538 60732 13544 60784
rect 13596 60732 13602 60784
rect 14274 60732 14280 60784
rect 14332 60732 14338 60784
rect 15746 60732 15752 60784
rect 15804 60732 15810 60784
rect 19426 60732 19432 60784
rect 19484 60732 19490 60784
rect 22097 60775 22155 60781
rect 22097 60741 22109 60775
rect 22143 60772 22155 60775
rect 22186 60772 22192 60784
rect 22143 60744 22192 60772
rect 22143 60741 22155 60744
rect 22097 60735 22155 60741
rect 22186 60732 22192 60744
rect 22244 60732 22250 60784
rect 23492 60781 23520 60812
rect 36170 60800 36176 60812
rect 36228 60800 36234 60852
rect 40218 60840 40224 60852
rect 36280 60812 40224 60840
rect 23477 60775 23535 60781
rect 23477 60741 23489 60775
rect 23523 60741 23535 60775
rect 23477 60735 23535 60741
rect 24394 60732 24400 60784
rect 24452 60772 24458 60784
rect 24581 60775 24639 60781
rect 24581 60772 24593 60775
rect 24452 60744 24593 60772
rect 24452 60732 24458 60744
rect 24581 60741 24593 60744
rect 24627 60741 24639 60775
rect 24581 60735 24639 60741
rect 24670 60732 24676 60784
rect 24728 60772 24734 60784
rect 36280 60772 36308 60812
rect 40218 60800 40224 60812
rect 40276 60800 40282 60852
rect 58894 60840 58900 60852
rect 56704 60812 58900 60840
rect 24728 60744 36308 60772
rect 24728 60732 24734 60744
rect 36354 60732 36360 60784
rect 36412 60732 36418 60784
rect 41506 60732 41512 60784
rect 41564 60732 41570 60784
rect 46658 60732 46664 60784
rect 46716 60732 46722 60784
rect 50154 60732 50160 60784
rect 50212 60772 50218 60784
rect 50341 60775 50399 60781
rect 50341 60772 50353 60775
rect 50212 60744 50353 60772
rect 50212 60732 50218 60744
rect 50341 60741 50353 60744
rect 50387 60741 50399 60775
rect 50341 60735 50399 60741
rect 52638 60732 52644 60784
rect 52696 60772 52702 60784
rect 53009 60775 53067 60781
rect 53009 60772 53021 60775
rect 52696 60744 53021 60772
rect 52696 60732 52702 60744
rect 53009 60741 53021 60744
rect 53055 60741 53067 60775
rect 53009 60735 53067 60741
rect 934 60664 940 60716
rect 992 60704 998 60716
rect 1581 60707 1639 60713
rect 1581 60704 1593 60707
rect 992 60676 1593 60704
rect 992 60664 998 60676
rect 1581 60673 1593 60676
rect 1627 60673 1639 60707
rect 1581 60667 1639 60673
rect 9030 60664 9036 60716
rect 9088 60664 9094 60716
rect 17862 60664 17868 60716
rect 17920 60704 17926 60716
rect 23201 60707 23259 60713
rect 23201 60704 23213 60707
rect 17920 60676 23213 60704
rect 17920 60664 17926 60676
rect 23201 60673 23213 60676
rect 23247 60673 23259 60707
rect 23201 60667 23259 60673
rect 23385 60707 23443 60713
rect 23385 60673 23397 60707
rect 23431 60673 23443 60707
rect 23385 60667 23443 60673
rect 23569 60707 23627 60713
rect 23569 60673 23581 60707
rect 23615 60704 23627 60707
rect 23658 60704 23664 60716
rect 23615 60676 23664 60704
rect 23615 60673 23627 60676
rect 23569 60667 23627 60673
rect 1857 60639 1915 60645
rect 1857 60605 1869 60639
rect 1903 60636 1915 60639
rect 7926 60636 7932 60648
rect 1903 60608 7932 60636
rect 1903 60605 1915 60608
rect 1857 60599 1915 60605
rect 7926 60596 7932 60608
rect 7984 60596 7990 60648
rect 8573 60639 8631 60645
rect 8573 60605 8585 60639
rect 8619 60636 8631 60639
rect 18414 60636 18420 60648
rect 8619 60608 18420 60636
rect 8619 60605 8631 60608
rect 8573 60599 8631 60605
rect 18414 60596 18420 60608
rect 18472 60596 18478 60648
rect 19610 60596 19616 60648
rect 19668 60636 19674 60648
rect 22186 60636 22192 60648
rect 19668 60608 22192 60636
rect 19668 60596 19674 60608
rect 22186 60596 22192 60608
rect 22244 60636 22250 60648
rect 23400 60636 23428 60667
rect 23658 60664 23664 60676
rect 23716 60664 23722 60716
rect 27522 60664 27528 60716
rect 27580 60664 27586 60716
rect 28994 60664 29000 60716
rect 29052 60664 29058 60716
rect 30466 60664 30472 60716
rect 30524 60664 30530 60716
rect 30558 60664 30564 60716
rect 30616 60704 30622 60716
rect 30616 60676 31754 60704
rect 30616 60664 30622 60676
rect 31202 60636 31208 60648
rect 22244 60608 23428 60636
rect 26896 60608 31208 60636
rect 22244 60596 22250 60608
rect 4157 60571 4215 60577
rect 4157 60537 4169 60571
rect 4203 60568 4215 60571
rect 4614 60568 4620 60580
rect 4203 60540 4620 60568
rect 4203 60537 4215 60540
rect 4157 60531 4215 60537
rect 4614 60528 4620 60540
rect 4672 60528 4678 60580
rect 14461 60571 14519 60577
rect 14461 60537 14473 60571
rect 14507 60568 14519 60571
rect 26896 60568 26924 60608
rect 31202 60596 31208 60608
rect 31260 60596 31266 60648
rect 31726 60636 31754 60676
rect 54662 60664 54668 60716
rect 54720 60664 54726 60716
rect 55401 60707 55459 60713
rect 55401 60673 55413 60707
rect 55447 60673 55459 60707
rect 55401 60667 55459 60673
rect 56137 60707 56195 60713
rect 56137 60673 56149 60707
rect 56183 60704 56195 60707
rect 56704 60704 56732 60812
rect 58894 60800 58900 60812
rect 58952 60800 58958 60852
rect 56778 60732 56784 60784
rect 56836 60772 56842 60784
rect 58986 60772 58992 60784
rect 56836 60744 58992 60772
rect 56836 60732 56842 60744
rect 58986 60732 58992 60744
rect 59044 60732 59050 60784
rect 56183 60676 56732 60704
rect 56183 60673 56195 60676
rect 56137 60667 56195 60673
rect 55416 60636 55444 60667
rect 56870 60664 56876 60716
rect 56928 60664 56934 60716
rect 58066 60664 58072 60716
rect 58124 60664 58130 60716
rect 56686 60636 56692 60648
rect 31726 60608 51074 60636
rect 55416 60608 56692 60636
rect 14507 60540 26924 60568
rect 27709 60571 27767 60577
rect 14507 60537 14519 60540
rect 14461 60531 14519 60537
rect 27709 60537 27721 60571
rect 27755 60568 27767 60571
rect 30653 60571 30711 60577
rect 27755 60540 30604 60568
rect 27755 60537 27767 60540
rect 27709 60531 27767 60537
rect 3326 60460 3332 60512
rect 3384 60460 3390 60512
rect 9214 60460 9220 60512
rect 9272 60460 9278 60512
rect 13633 60503 13691 60509
rect 13633 60469 13645 60503
rect 13679 60500 13691 60503
rect 15102 60500 15108 60512
rect 13679 60472 15108 60500
rect 13679 60469 13691 60472
rect 13633 60463 13691 60469
rect 15102 60460 15108 60472
rect 15160 60460 15166 60512
rect 15841 60503 15899 60509
rect 15841 60469 15853 60503
rect 15887 60500 15899 60503
rect 17862 60500 17868 60512
rect 15887 60472 17868 60500
rect 15887 60469 15899 60472
rect 15841 60463 15899 60469
rect 17862 60460 17868 60472
rect 17920 60460 17926 60512
rect 19521 60503 19579 60509
rect 19521 60469 19533 60503
rect 19567 60500 19579 60503
rect 20070 60500 20076 60512
rect 19567 60472 20076 60500
rect 19567 60469 19579 60472
rect 19521 60463 19579 60469
rect 20070 60460 20076 60472
rect 20128 60460 20134 60512
rect 22278 60460 22284 60512
rect 22336 60500 22342 60512
rect 22373 60503 22431 60509
rect 22373 60500 22385 60503
rect 22336 60472 22385 60500
rect 22336 60460 22342 60472
rect 22373 60469 22385 60472
rect 22419 60469 22431 60503
rect 22373 60463 22431 60469
rect 23753 60503 23811 60509
rect 23753 60469 23765 60503
rect 23799 60500 23811 60503
rect 24394 60500 24400 60512
rect 23799 60472 24400 60500
rect 23799 60469 23811 60472
rect 23753 60463 23811 60469
rect 24394 60460 24400 60472
rect 24452 60460 24458 60512
rect 24670 60460 24676 60512
rect 24728 60460 24734 60512
rect 24854 60460 24860 60512
rect 24912 60500 24918 60512
rect 28994 60500 29000 60512
rect 24912 60472 29000 60500
rect 24912 60460 24918 60472
rect 28994 60460 29000 60472
rect 29052 60460 29058 60512
rect 29089 60503 29147 60509
rect 29089 60469 29101 60503
rect 29135 60500 29147 60503
rect 29822 60500 29828 60512
rect 29135 60472 29828 60500
rect 29135 60469 29147 60472
rect 29089 60463 29147 60469
rect 29822 60460 29828 60472
rect 29880 60460 29886 60512
rect 30006 60460 30012 60512
rect 30064 60460 30070 60512
rect 30576 60500 30604 60540
rect 30653 60537 30665 60571
rect 30699 60568 30711 60571
rect 42242 60568 42248 60580
rect 30699 60540 42248 60568
rect 30699 60537 30711 60540
rect 30653 60531 30711 60537
rect 42242 60528 42248 60540
rect 42300 60528 42306 60580
rect 51046 60568 51074 60608
rect 56686 60596 56692 60608
rect 56744 60596 56750 60648
rect 58158 60568 58164 60580
rect 51046 60540 58164 60568
rect 58158 60528 58164 60540
rect 58216 60528 58222 60580
rect 30926 60500 30932 60512
rect 30576 60472 30932 60500
rect 30926 60460 30932 60472
rect 30984 60460 30990 60512
rect 35710 60460 35716 60512
rect 35768 60500 35774 60512
rect 36449 60503 36507 60509
rect 36449 60500 36461 60503
rect 35768 60472 36461 60500
rect 35768 60460 35774 60472
rect 36449 60469 36461 60472
rect 36495 60469 36507 60503
rect 36449 60463 36507 60469
rect 40954 60460 40960 60512
rect 41012 60500 41018 60512
rect 41601 60503 41659 60509
rect 41601 60500 41613 60503
rect 41012 60472 41613 60500
rect 41012 60460 41018 60472
rect 41601 60469 41613 60472
rect 41647 60469 41659 60503
rect 41601 60463 41659 60469
rect 44174 60460 44180 60512
rect 44232 60500 44238 60512
rect 46753 60503 46811 60509
rect 46753 60500 46765 60503
rect 44232 60472 46765 60500
rect 44232 60460 44238 60472
rect 46753 60469 46765 60472
rect 46799 60469 46811 60503
rect 46753 60463 46811 60469
rect 50430 60460 50436 60512
rect 50488 60460 50494 60512
rect 53098 60460 53104 60512
rect 53156 60460 53162 60512
rect 54846 60460 54852 60512
rect 54904 60460 54910 60512
rect 55582 60460 55588 60512
rect 55640 60460 55646 60512
rect 56318 60460 56324 60512
rect 56376 60460 56382 60512
rect 57054 60460 57060 60512
rect 57112 60460 57118 60512
rect 58250 60460 58256 60512
rect 58308 60460 58314 60512
rect 1104 60410 58880 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 58880 60410
rect 1104 60336 58880 60358
rect 3326 60256 3332 60308
rect 3384 60296 3390 60308
rect 20254 60296 20260 60308
rect 3384 60268 20260 60296
rect 3384 60256 3390 60268
rect 20254 60256 20260 60268
rect 20312 60256 20318 60308
rect 58250 60296 58256 60308
rect 22480 60268 58256 60296
rect 15102 60188 15108 60240
rect 15160 60228 15166 60240
rect 19242 60228 19248 60240
rect 15160 60200 19248 60228
rect 15160 60188 15166 60200
rect 19242 60188 19248 60200
rect 19300 60188 19306 60240
rect 19981 60231 20039 60237
rect 19981 60197 19993 60231
rect 20027 60228 20039 60231
rect 20162 60228 20168 60240
rect 20027 60200 20168 60228
rect 20027 60197 20039 60200
rect 19981 60191 20039 60197
rect 20162 60188 20168 60200
rect 20220 60188 20226 60240
rect 21177 60231 21235 60237
rect 21177 60197 21189 60231
rect 21223 60228 21235 60231
rect 21910 60228 21916 60240
rect 21223 60200 21916 60228
rect 21223 60197 21235 60200
rect 21177 60191 21235 60197
rect 21910 60188 21916 60200
rect 21968 60188 21974 60240
rect 17862 60120 17868 60172
rect 17920 60120 17926 60172
rect 18138 60120 18144 60172
rect 18196 60160 18202 60172
rect 18325 60163 18383 60169
rect 18325 60160 18337 60163
rect 18196 60132 18337 60160
rect 18196 60120 18202 60132
rect 18325 60129 18337 60132
rect 18371 60129 18383 60163
rect 22002 60160 22008 60172
rect 18325 60123 18383 60129
rect 19720 60132 22008 60160
rect 2590 60052 2596 60104
rect 2648 60052 2654 60104
rect 5626 60052 5632 60104
rect 5684 60092 5690 60104
rect 7377 60095 7435 60101
rect 7377 60092 7389 60095
rect 5684 60064 7389 60092
rect 5684 60052 5690 60064
rect 7377 60061 7389 60064
rect 7423 60061 7435 60095
rect 7377 60055 7435 60061
rect 7742 60052 7748 60104
rect 7800 60052 7806 60104
rect 18049 60095 18107 60101
rect 18049 60061 18061 60095
rect 18095 60092 18107 60095
rect 18095 60064 18368 60092
rect 18095 60061 18107 60064
rect 18049 60055 18107 60061
rect 934 59984 940 60036
rect 992 60024 998 60036
rect 1673 60027 1731 60033
rect 1673 60024 1685 60027
rect 992 59996 1685 60024
rect 992 59984 998 59996
rect 1673 59993 1685 59996
rect 1719 59993 1731 60027
rect 1673 59987 1731 59993
rect 2038 59984 2044 60036
rect 2096 59984 2102 60036
rect 7558 59984 7564 60036
rect 7616 59984 7622 60036
rect 7653 60027 7711 60033
rect 7653 59993 7665 60027
rect 7699 60024 7711 60027
rect 8202 60024 8208 60036
rect 7699 59996 8208 60024
rect 7699 59993 7711 59996
rect 7653 59987 7711 59993
rect 8202 59984 8208 59996
rect 8260 59984 8266 60036
rect 2498 59916 2504 59968
rect 2556 59956 2562 59968
rect 2685 59959 2743 59965
rect 2685 59956 2697 59959
rect 2556 59928 2697 59956
rect 2556 59916 2562 59928
rect 2685 59925 2697 59928
rect 2731 59925 2743 59959
rect 2685 59919 2743 59925
rect 7929 59959 7987 59965
rect 7929 59925 7941 59959
rect 7975 59956 7987 59959
rect 8018 59956 8024 59968
rect 7975 59928 8024 59956
rect 7975 59925 7987 59928
rect 7929 59919 7987 59925
rect 8018 59916 8024 59928
rect 8076 59916 8082 59968
rect 17586 59916 17592 59968
rect 17644 59956 17650 59968
rect 17681 59959 17739 59965
rect 17681 59956 17693 59959
rect 17644 59928 17693 59956
rect 17644 59916 17650 59928
rect 17681 59925 17693 59928
rect 17727 59925 17739 59959
rect 18340 59956 18368 60064
rect 18414 60052 18420 60104
rect 18472 60052 18478 60104
rect 18506 60052 18512 60104
rect 18564 60092 18570 60104
rect 19429 60095 19487 60101
rect 19429 60092 19441 60095
rect 18564 60064 19441 60092
rect 18564 60052 18570 60064
rect 19429 60061 19441 60064
rect 19475 60061 19487 60095
rect 19610 60092 19616 60104
rect 19429 60055 19487 60061
rect 19536 60064 19616 60092
rect 19150 59984 19156 60036
rect 19208 60024 19214 60036
rect 19536 60024 19564 60064
rect 19610 60052 19616 60064
rect 19668 60052 19674 60104
rect 19720 60101 19748 60132
rect 22002 60120 22008 60132
rect 22060 60120 22066 60172
rect 19886 60101 19892 60104
rect 19705 60095 19763 60101
rect 19705 60061 19717 60095
rect 19751 60061 19763 60095
rect 19705 60055 19763 60061
rect 19849 60095 19892 60101
rect 19849 60061 19861 60095
rect 19849 60055 19892 60061
rect 19886 60052 19892 60055
rect 19944 60052 19950 60104
rect 19978 60052 19984 60104
rect 20036 60092 20042 60104
rect 20625 60095 20683 60101
rect 20625 60092 20637 60095
rect 20036 60064 20637 60092
rect 20036 60052 20042 60064
rect 20625 60061 20637 60064
rect 20671 60061 20683 60095
rect 20625 60055 20683 60061
rect 21045 60095 21103 60101
rect 21045 60061 21057 60095
rect 21091 60092 21103 60095
rect 22189 60095 22247 60101
rect 22189 60092 22201 60095
rect 21091 60064 22201 60092
rect 21091 60061 21103 60064
rect 21045 60055 21103 60061
rect 22189 60061 22201 60064
rect 22235 60092 22247 60095
rect 22278 60092 22284 60104
rect 22235 60064 22284 60092
rect 22235 60061 22247 60064
rect 22189 60055 22247 60061
rect 22278 60052 22284 60064
rect 22336 60052 22342 60104
rect 22480 60101 22508 60268
rect 58250 60256 58256 60268
rect 58308 60256 58314 60308
rect 23290 60188 23296 60240
rect 23348 60228 23354 60240
rect 30558 60228 30564 60240
rect 23348 60200 30564 60228
rect 23348 60188 23354 60200
rect 30558 60188 30564 60200
rect 30616 60188 30622 60240
rect 30742 60188 30748 60240
rect 30800 60228 30806 60240
rect 41138 60228 41144 60240
rect 30800 60200 41144 60228
rect 30800 60188 30806 60200
rect 41138 60188 41144 60200
rect 41196 60188 41202 60240
rect 41230 60188 41236 60240
rect 41288 60188 41294 60240
rect 41598 60188 41604 60240
rect 41656 60228 41662 60240
rect 41656 60200 42748 60228
rect 41656 60188 41662 60200
rect 42720 60172 42748 60200
rect 24854 60160 24860 60172
rect 22848 60132 24860 60160
rect 22848 60104 22876 60132
rect 24854 60120 24860 60132
rect 24912 60120 24918 60172
rect 29086 60160 29092 60172
rect 28092 60132 29092 60160
rect 22465 60095 22523 60101
rect 22465 60061 22477 60095
rect 22511 60061 22523 60095
rect 22465 60055 22523 60061
rect 22554 60052 22560 60104
rect 22612 60052 22618 60104
rect 22830 60052 22836 60104
rect 22888 60052 22894 60104
rect 23014 60052 23020 60104
rect 23072 60052 23078 60104
rect 23198 60052 23204 60104
rect 23256 60092 23262 60104
rect 28092 60101 28120 60132
rect 29086 60120 29092 60132
rect 29144 60120 29150 60172
rect 29178 60120 29184 60172
rect 29236 60160 29242 60172
rect 29236 60132 30880 60160
rect 29236 60120 29242 60132
rect 23661 60095 23719 60101
rect 23661 60092 23673 60095
rect 23256 60064 23673 60092
rect 23256 60052 23262 60064
rect 23661 60061 23673 60064
rect 23707 60061 23719 60095
rect 23661 60055 23719 60061
rect 27801 60095 27859 60101
rect 27801 60061 27813 60095
rect 27847 60092 27859 60095
rect 28077 60095 28135 60101
rect 28077 60092 28089 60095
rect 27847 60064 28089 60092
rect 27847 60061 27859 60064
rect 27801 60055 27859 60061
rect 28077 60061 28089 60064
rect 28123 60061 28135 60095
rect 28077 60055 28135 60061
rect 28166 60052 28172 60104
rect 28224 60052 28230 60104
rect 28542 60095 28600 60101
rect 28542 60092 28554 60095
rect 28276 60064 28554 60092
rect 20806 60024 20812 60036
rect 19208 59996 19564 60024
rect 19812 59996 20812 60024
rect 19208 59984 19214 59996
rect 19812 59956 19840 59996
rect 20806 59984 20812 59996
rect 20864 59984 20870 60036
rect 20898 59984 20904 60036
rect 20956 59984 20962 60036
rect 28276 60024 28304 60064
rect 28542 60061 28554 60064
rect 28588 60092 28600 60095
rect 30190 60092 30196 60104
rect 28588 60064 30196 60092
rect 28588 60061 28600 60064
rect 28542 60055 28600 60061
rect 30190 60052 30196 60064
rect 30248 60092 30254 60104
rect 30628 60095 30686 60101
rect 30628 60092 30640 60095
rect 30248 60064 30640 60092
rect 30248 60052 30254 60064
rect 30628 60061 30640 60064
rect 30674 60061 30686 60095
rect 30628 60055 30686 60061
rect 30742 60052 30748 60104
rect 30800 60052 30806 60104
rect 23676 59996 28304 60024
rect 28353 60027 28411 60033
rect 23676 59968 23704 59996
rect 28353 59993 28365 60027
rect 28399 59993 28411 60027
rect 28353 59987 28411 59993
rect 28445 60027 28503 60033
rect 28445 59993 28457 60027
rect 28491 60024 28503 60027
rect 28902 60024 28908 60036
rect 28491 59996 28908 60024
rect 28491 59993 28503 59996
rect 28445 59987 28503 59993
rect 18340 59928 19840 59956
rect 17681 59919 17739 59925
rect 19886 59916 19892 59968
rect 19944 59956 19950 59968
rect 19978 59956 19984 59968
rect 19944 59928 19984 59956
rect 19944 59916 19950 59928
rect 19978 59916 19984 59928
rect 20036 59956 20042 59968
rect 21266 59956 21272 59968
rect 20036 59928 21272 59956
rect 20036 59916 20042 59928
rect 21266 59916 21272 59928
rect 21324 59916 21330 59968
rect 21818 59916 21824 59968
rect 21876 59916 21882 59968
rect 22278 59916 22284 59968
rect 22336 59956 22342 59968
rect 23382 59956 23388 59968
rect 22336 59928 23388 59956
rect 22336 59916 22342 59928
rect 23382 59916 23388 59928
rect 23440 59916 23446 59968
rect 23658 59916 23664 59968
rect 23716 59916 23722 59968
rect 23750 59916 23756 59968
rect 23808 59956 23814 59968
rect 23845 59959 23903 59965
rect 23845 59956 23857 59959
rect 23808 59928 23857 59956
rect 23808 59916 23814 59928
rect 23845 59925 23857 59928
rect 23891 59925 23903 59959
rect 28368 59956 28396 59987
rect 28902 59984 28908 59996
rect 28960 59984 28966 60036
rect 30006 59984 30012 60036
rect 30064 60024 30070 60036
rect 30852 60033 30880 60132
rect 40696 60132 42196 60160
rect 30926 60052 30932 60104
rect 30984 60101 30990 60104
rect 30984 60095 31023 60101
rect 31011 60061 31023 60095
rect 30984 60055 31023 60061
rect 30984 60052 30990 60055
rect 31110 60052 31116 60104
rect 31168 60052 31174 60104
rect 31202 60052 31208 60104
rect 31260 60092 31266 60104
rect 32401 60095 32459 60101
rect 32401 60092 32413 60095
rect 31260 60064 32413 60092
rect 31260 60052 31266 60064
rect 32401 60061 32413 60064
rect 32447 60061 32459 60095
rect 32401 60055 32459 60061
rect 32585 60095 32643 60101
rect 32585 60061 32597 60095
rect 32631 60061 32643 60095
rect 32585 60055 32643 60061
rect 30101 60027 30159 60033
rect 30101 60024 30113 60027
rect 30064 59996 30113 60024
rect 30064 59984 30070 59996
rect 30101 59993 30113 59996
rect 30147 60024 30159 60027
rect 30837 60027 30895 60033
rect 30147 59996 30604 60024
rect 30147 59993 30159 59996
rect 30101 59987 30159 59993
rect 28626 59956 28632 59968
rect 28368 59928 28632 59956
rect 23845 59919 23903 59925
rect 28626 59916 28632 59928
rect 28684 59916 28690 59968
rect 28718 59916 28724 59968
rect 28776 59916 28782 59968
rect 29086 59916 29092 59968
rect 29144 59916 29150 59968
rect 30466 59916 30472 59968
rect 30524 59916 30530 59968
rect 30576 59956 30604 59996
rect 30837 59993 30849 60027
rect 30883 59993 30895 60027
rect 30837 59987 30895 59993
rect 31128 59956 31156 60052
rect 30576 59928 31156 59956
rect 31665 59959 31723 59965
rect 31665 59925 31677 59959
rect 31711 59956 31723 59959
rect 32214 59956 32220 59968
rect 31711 59928 32220 59956
rect 31711 59925 31723 59928
rect 31665 59919 31723 59925
rect 32214 59916 32220 59928
rect 32272 59916 32278 59968
rect 32490 59916 32496 59968
rect 32548 59956 32554 59968
rect 32600 59956 32628 60055
rect 32950 60052 32956 60104
rect 33008 60052 33014 60104
rect 33045 60095 33103 60101
rect 33045 60061 33057 60095
rect 33091 60092 33103 60095
rect 34514 60092 34520 60104
rect 33091 60064 34520 60092
rect 33091 60061 33103 60064
rect 33045 60055 33103 60061
rect 34514 60052 34520 60064
rect 34572 60052 34578 60104
rect 40696 60101 40724 60132
rect 40681 60095 40739 60101
rect 40681 60061 40693 60095
rect 40727 60061 40739 60095
rect 40681 60055 40739 60061
rect 40954 60052 40960 60104
rect 41012 60052 41018 60104
rect 41101 60095 41159 60101
rect 41101 60061 41113 60095
rect 41147 60092 41159 60095
rect 41598 60092 41604 60104
rect 41147 60064 41604 60092
rect 41147 60061 41159 60064
rect 41101 60055 41159 60061
rect 41598 60052 41604 60064
rect 41656 60052 41662 60104
rect 40862 59984 40868 60036
rect 40920 59984 40926 60036
rect 41785 60027 41843 60033
rect 41785 59993 41797 60027
rect 41831 60024 41843 60027
rect 42058 60024 42064 60036
rect 41831 59996 42064 60024
rect 41831 59993 41843 59996
rect 41785 59987 41843 59993
rect 42058 59984 42064 59996
rect 42116 59984 42122 60036
rect 42168 60024 42196 60132
rect 42242 60120 42248 60172
rect 42300 60120 42306 60172
rect 42702 60120 42708 60172
rect 42760 60120 42766 60172
rect 50430 60160 50436 60172
rect 42812 60132 50436 60160
rect 42426 60052 42432 60104
rect 42484 60052 42490 60104
rect 42812 60101 42840 60132
rect 50430 60120 50436 60132
rect 50488 60120 50494 60172
rect 56226 60160 56232 60172
rect 55186 60132 56232 60160
rect 42797 60095 42855 60101
rect 42797 60061 42809 60095
rect 42843 60061 42855 60095
rect 42797 60055 42855 60061
rect 42168 59996 51074 60024
rect 33042 59956 33048 59968
rect 32548 59928 33048 59956
rect 32548 59916 32554 59928
rect 33042 59916 33048 59928
rect 33100 59956 33106 59968
rect 42426 59956 42432 59968
rect 33100 59928 42432 59956
rect 33100 59916 33106 59928
rect 42426 59916 42432 59928
rect 42484 59916 42490 59968
rect 51046 59956 51074 59996
rect 55186 59956 55214 60132
rect 56226 60120 56232 60132
rect 56284 60120 56290 60172
rect 58986 60160 58992 60172
rect 57256 60132 58992 60160
rect 56505 60095 56563 60101
rect 56505 60061 56517 60095
rect 56551 60092 56563 60095
rect 56778 60092 56784 60104
rect 56551 60064 56784 60092
rect 56551 60061 56563 60064
rect 56505 60055 56563 60061
rect 56778 60052 56784 60064
rect 56836 60052 56842 60104
rect 57256 60101 57284 60132
rect 58986 60120 58992 60132
rect 59044 60120 59050 60172
rect 57241 60095 57299 60101
rect 57241 60061 57253 60095
rect 57287 60061 57299 60095
rect 57241 60055 57299 60061
rect 57885 60095 57943 60101
rect 57885 60061 57897 60095
rect 57931 60092 57943 60095
rect 57974 60092 57980 60104
rect 57931 60064 57980 60092
rect 57931 60061 57943 60064
rect 57885 60055 57943 60061
rect 57974 60052 57980 60064
rect 58032 60052 58038 60104
rect 56686 59984 56692 60036
rect 56744 59984 56750 60036
rect 58161 60027 58219 60033
rect 58161 59993 58173 60027
rect 58207 60024 58219 60027
rect 59538 60024 59544 60036
rect 58207 59996 59544 60024
rect 58207 59993 58219 59996
rect 58161 59987 58219 59993
rect 59538 59984 59544 59996
rect 59596 59984 59602 60036
rect 51046 59928 55214 59956
rect 57330 59916 57336 59968
rect 57388 59916 57394 59968
rect 1104 59866 58880 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 58880 59866
rect 1104 59792 58880 59814
rect 7742 59712 7748 59764
rect 7800 59752 7806 59764
rect 19978 59752 19984 59764
rect 7800 59724 19984 59752
rect 7800 59712 7806 59724
rect 19978 59712 19984 59724
rect 20036 59712 20042 59764
rect 20898 59712 20904 59764
rect 20956 59752 20962 59764
rect 55582 59752 55588 59764
rect 20956 59724 55588 59752
rect 20956 59712 20962 59724
rect 55582 59712 55588 59724
rect 55640 59712 55646 59764
rect 56226 59712 56232 59764
rect 56284 59752 56290 59764
rect 57425 59755 57483 59761
rect 57425 59752 57437 59755
rect 56284 59724 57437 59752
rect 56284 59712 56290 59724
rect 57425 59721 57437 59724
rect 57471 59721 57483 59755
rect 57425 59715 57483 59721
rect 58158 59712 58164 59764
rect 58216 59752 58222 59764
rect 58253 59755 58311 59761
rect 58253 59752 58265 59755
rect 58216 59724 58265 59752
rect 58216 59712 58222 59724
rect 58253 59721 58265 59724
rect 58299 59721 58311 59755
rect 58253 59715 58311 59721
rect 1578 59644 1584 59696
rect 1636 59684 1642 59696
rect 2593 59687 2651 59693
rect 2593 59684 2605 59687
rect 1636 59656 2605 59684
rect 1636 59644 1642 59656
rect 2593 59653 2605 59656
rect 2639 59653 2651 59687
rect 2593 59647 2651 59653
rect 7558 59644 7564 59696
rect 7616 59684 7622 59696
rect 19150 59684 19156 59696
rect 7616 59656 19156 59684
rect 7616 59644 7622 59656
rect 19150 59644 19156 59656
rect 19208 59644 19214 59696
rect 21085 59687 21143 59693
rect 21085 59653 21097 59687
rect 21131 59684 21143 59687
rect 21358 59684 21364 59696
rect 21131 59656 21364 59684
rect 21131 59653 21143 59656
rect 21085 59647 21143 59653
rect 21358 59644 21364 59656
rect 21416 59644 21422 59696
rect 22281 59687 22339 59693
rect 22281 59653 22293 59687
rect 22327 59684 22339 59687
rect 22830 59684 22836 59696
rect 22327 59656 22836 59684
rect 22327 59653 22339 59656
rect 22281 59647 22339 59653
rect 934 59576 940 59628
rect 992 59616 998 59628
rect 1673 59619 1731 59625
rect 1673 59616 1685 59619
rect 992 59588 1685 59616
rect 992 59576 998 59588
rect 1673 59585 1685 59588
rect 1719 59585 1731 59619
rect 1673 59579 1731 59585
rect 18046 59576 18052 59628
rect 18104 59616 18110 59628
rect 20901 59619 20959 59625
rect 20901 59616 20913 59619
rect 18104 59588 20913 59616
rect 18104 59576 18110 59588
rect 20901 59585 20913 59588
rect 20947 59585 20959 59619
rect 20901 59579 20959 59585
rect 21174 59576 21180 59628
rect 21232 59576 21238 59628
rect 21266 59576 21272 59628
rect 21324 59576 21330 59628
rect 22094 59576 22100 59628
rect 22152 59576 22158 59628
rect 20806 59508 20812 59560
rect 20864 59548 20870 59560
rect 22296 59548 22324 59647
rect 22830 59644 22836 59656
rect 22888 59644 22894 59696
rect 29454 59684 29460 59696
rect 23124 59656 29460 59684
rect 22373 59619 22431 59625
rect 22373 59585 22385 59619
rect 22419 59585 22431 59619
rect 22373 59579 22431 59585
rect 22517 59619 22575 59625
rect 22517 59585 22529 59619
rect 22563 59616 22575 59619
rect 23124 59616 23152 59656
rect 29454 59644 29460 59656
rect 29512 59644 29518 59696
rect 29564 59656 30052 59684
rect 22563 59588 23152 59616
rect 23201 59619 23259 59625
rect 22563 59585 22575 59588
rect 22517 59579 22575 59585
rect 23201 59585 23213 59619
rect 23247 59616 23259 59619
rect 23290 59616 23296 59628
rect 23247 59588 23296 59616
rect 23247 59585 23259 59588
rect 23201 59579 23259 59585
rect 20864 59520 22324 59548
rect 22388 59548 22416 59579
rect 23290 59576 23296 59588
rect 23348 59576 23354 59628
rect 23382 59576 23388 59628
rect 23440 59576 23446 59628
rect 23474 59576 23480 59628
rect 23532 59576 23538 59628
rect 23566 59576 23572 59628
rect 23624 59625 23630 59628
rect 23624 59579 23632 59625
rect 23624 59576 23630 59579
rect 28350 59576 28356 59628
rect 28408 59576 28414 59628
rect 28626 59576 28632 59628
rect 28684 59616 28690 59628
rect 29564 59616 29592 59656
rect 30024 59628 30052 59656
rect 30098 59644 30104 59696
rect 30156 59644 30162 59696
rect 30282 59644 30288 59696
rect 30340 59684 30346 59696
rect 30340 59656 41414 59684
rect 30340 59644 30346 59656
rect 28684 59588 29592 59616
rect 28684 59576 28690 59588
rect 29730 59576 29736 59628
rect 29788 59576 29794 59628
rect 29822 59576 29828 59628
rect 29880 59616 29886 59628
rect 29880 59588 29925 59616
rect 29880 59576 29886 59588
rect 30006 59576 30012 59628
rect 30064 59576 30070 59628
rect 30190 59576 30196 59628
rect 30248 59625 30254 59628
rect 30248 59616 30256 59625
rect 34514 59616 34520 59628
rect 30248 59588 34520 59616
rect 30248 59579 30256 59588
rect 30248 59576 30254 59579
rect 34514 59576 34520 59588
rect 34572 59576 34578 59628
rect 22388 59520 29592 59548
rect 20864 59508 20870 59520
rect 21453 59483 21511 59489
rect 21453 59449 21465 59483
rect 21499 59480 21511 59483
rect 22554 59480 22560 59492
rect 21499 59452 22560 59480
rect 21499 59449 21511 59452
rect 21453 59443 21511 59449
rect 22554 59440 22560 59452
rect 22612 59440 22618 59492
rect 23382 59440 23388 59492
rect 23440 59480 23446 59492
rect 24854 59480 24860 59492
rect 23440 59452 24860 59480
rect 23440 59440 23446 59452
rect 24854 59440 24860 59452
rect 24912 59440 24918 59492
rect 29564 59480 29592 59520
rect 29638 59508 29644 59560
rect 29696 59548 29702 59560
rect 29696 59520 31754 59548
rect 29696 59508 29702 59520
rect 30282 59480 30288 59492
rect 29564 59452 30288 59480
rect 30282 59440 30288 59452
rect 30340 59440 30346 59492
rect 30374 59440 30380 59492
rect 30432 59440 30438 59492
rect 31726 59480 31754 59520
rect 40862 59480 40868 59492
rect 30484 59452 30788 59480
rect 31726 59452 40868 59480
rect 1946 59372 1952 59424
rect 2004 59372 2010 59424
rect 2314 59372 2320 59424
rect 2372 59412 2378 59424
rect 2685 59415 2743 59421
rect 2685 59412 2697 59415
rect 2372 59384 2697 59412
rect 2372 59372 2378 59384
rect 2685 59381 2697 59384
rect 2731 59381 2743 59415
rect 2685 59375 2743 59381
rect 19242 59372 19248 59424
rect 19300 59412 19306 59424
rect 22462 59412 22468 59424
rect 19300 59384 22468 59412
rect 19300 59372 19306 59384
rect 22462 59372 22468 59384
rect 22520 59372 22526 59424
rect 22649 59415 22707 59421
rect 22649 59381 22661 59415
rect 22695 59412 22707 59415
rect 22922 59412 22928 59424
rect 22695 59384 22928 59412
rect 22695 59381 22707 59384
rect 22649 59375 22707 59381
rect 22922 59372 22928 59384
rect 22980 59372 22986 59424
rect 23753 59415 23811 59421
rect 23753 59381 23765 59415
rect 23799 59412 23811 59415
rect 24486 59412 24492 59424
rect 23799 59384 24492 59412
rect 23799 59381 23811 59384
rect 23753 59375 23811 59381
rect 24486 59372 24492 59384
rect 24544 59372 24550 59424
rect 29457 59415 29515 59421
rect 29457 59381 29469 59415
rect 29503 59412 29515 59415
rect 29730 59412 29736 59424
rect 29503 59384 29736 59412
rect 29503 59381 29515 59384
rect 29457 59375 29515 59381
rect 29730 59372 29736 59384
rect 29788 59372 29794 59424
rect 30006 59372 30012 59424
rect 30064 59412 30070 59424
rect 30484 59412 30512 59452
rect 30064 59384 30512 59412
rect 30064 59372 30070 59384
rect 30650 59372 30656 59424
rect 30708 59372 30714 59424
rect 30760 59412 30788 59452
rect 40862 59440 40868 59452
rect 40920 59440 40926 59492
rect 41386 59480 41414 59656
rect 42426 59644 42432 59696
rect 42484 59684 42490 59696
rect 57333 59687 57391 59693
rect 42484 59656 43300 59684
rect 42484 59644 42490 59656
rect 41782 59576 41788 59628
rect 41840 59616 41846 59628
rect 43272 59625 43300 59656
rect 57333 59653 57345 59687
rect 57379 59684 57391 59687
rect 58802 59684 58808 59696
rect 57379 59656 58808 59684
rect 57379 59653 57391 59656
rect 57333 59647 57391 59653
rect 58802 59644 58808 59656
rect 58860 59644 58866 59696
rect 43073 59619 43131 59625
rect 43073 59616 43085 59619
rect 41840 59588 43085 59616
rect 41840 59576 41846 59588
rect 43073 59585 43085 59588
rect 43119 59585 43131 59619
rect 43073 59579 43131 59585
rect 43257 59619 43315 59625
rect 43257 59585 43269 59619
rect 43303 59585 43315 59619
rect 43257 59579 43315 59585
rect 43625 59619 43683 59625
rect 43625 59585 43637 59619
rect 43671 59616 43683 59619
rect 53098 59616 53104 59628
rect 43671 59588 53104 59616
rect 43671 59585 43683 59588
rect 43625 59579 43683 59585
rect 53098 59576 53104 59588
rect 53156 59576 53162 59628
rect 58066 59576 58072 59628
rect 58124 59576 58130 59628
rect 42702 59508 42708 59560
rect 42760 59508 42766 59560
rect 42794 59508 42800 59560
rect 42852 59548 42858 59560
rect 43533 59551 43591 59557
rect 43533 59548 43545 59551
rect 42852 59520 43545 59548
rect 42852 59508 42858 59520
rect 43533 59517 43545 59520
rect 43579 59517 43591 59551
rect 56318 59548 56324 59560
rect 43533 59511 43591 59517
rect 51046 59520 56324 59548
rect 51046 59480 51074 59520
rect 56318 59508 56324 59520
rect 56376 59508 56382 59560
rect 41386 59452 51074 59480
rect 57146 59440 57152 59492
rect 57204 59480 57210 59492
rect 58710 59480 58716 59492
rect 57204 59452 58716 59480
rect 57204 59440 57210 59452
rect 58710 59440 58716 59452
rect 58768 59440 58774 59492
rect 32490 59412 32496 59424
rect 30760 59384 32496 59412
rect 32490 59372 32496 59384
rect 32548 59372 32554 59424
rect 1104 59322 58880 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 58880 59322
rect 1104 59248 58880 59270
rect 57333 59211 57391 59217
rect 57333 59208 57345 59211
rect 19444 59180 57345 59208
rect 1946 59032 1952 59084
rect 2004 59072 2010 59084
rect 2004 59044 6914 59072
rect 2004 59032 2010 59044
rect 842 58964 848 59016
rect 900 59004 906 59016
rect 1673 59007 1731 59013
rect 1673 59004 1685 59007
rect 900 58976 1685 59004
rect 900 58964 906 58976
rect 1673 58973 1685 58976
rect 1719 58973 1731 59007
rect 1673 58967 1731 58973
rect 6886 58936 6914 59044
rect 19444 59013 19472 59180
rect 57333 59177 57345 59180
rect 57379 59177 57391 59211
rect 57333 59171 57391 59177
rect 19518 59100 19524 59152
rect 19576 59140 19582 59152
rect 19981 59143 20039 59149
rect 19981 59140 19993 59143
rect 19576 59112 19993 59140
rect 19576 59100 19582 59112
rect 19981 59109 19993 59112
rect 20027 59109 20039 59143
rect 19981 59103 20039 59109
rect 38838 59100 38844 59152
rect 38896 59140 38902 59152
rect 58342 59140 58348 59152
rect 38896 59112 58348 59140
rect 38896 59100 38902 59112
rect 58342 59100 58348 59112
rect 58400 59100 58406 59152
rect 41325 59075 41383 59081
rect 41325 59072 41337 59075
rect 19536 59044 41337 59072
rect 19429 59007 19487 59013
rect 19429 58973 19441 59007
rect 19475 58973 19487 59007
rect 19429 58967 19487 58973
rect 19536 58936 19564 59044
rect 41325 59041 41337 59044
rect 41371 59041 41383 59075
rect 41325 59035 41383 59041
rect 41598 59032 41604 59084
rect 41656 59072 41662 59084
rect 41785 59075 41843 59081
rect 41785 59072 41797 59075
rect 41656 59044 41797 59072
rect 41656 59032 41662 59044
rect 41785 59041 41797 59044
rect 41831 59041 41843 59075
rect 50614 59072 50620 59084
rect 41785 59035 41843 59041
rect 41892 59044 50620 59072
rect 19702 58964 19708 59016
rect 19760 58964 19766 59016
rect 19849 59007 19907 59013
rect 19849 58973 19861 59007
rect 19895 59004 19907 59007
rect 21358 59004 21364 59016
rect 19895 58976 21364 59004
rect 19895 58973 19907 58976
rect 19849 58967 19907 58973
rect 21358 58964 21364 58976
rect 21416 59004 21422 59016
rect 23566 59004 23572 59016
rect 21416 58976 23572 59004
rect 21416 58964 21422 58976
rect 23566 58964 23572 58976
rect 23624 58964 23630 59016
rect 41506 58964 41512 59016
rect 41564 58964 41570 59016
rect 41892 59013 41920 59044
rect 50614 59032 50620 59044
rect 50672 59032 50678 59084
rect 41877 59007 41935 59013
rect 41877 58973 41889 59007
rect 41923 58973 41935 59007
rect 41877 58967 41935 58973
rect 57146 58964 57152 59016
rect 57204 58964 57210 59016
rect 57885 59007 57943 59013
rect 57885 58973 57897 59007
rect 57931 59004 57943 59007
rect 58986 59004 58992 59016
rect 57931 58976 58992 59004
rect 57931 58973 57943 58976
rect 57885 58967 57943 58973
rect 58986 58964 58992 58976
rect 59044 58964 59050 59016
rect 6886 58908 19564 58936
rect 19613 58939 19671 58945
rect 19613 58905 19625 58939
rect 19659 58905 19671 58939
rect 19613 58899 19671 58905
rect 58161 58939 58219 58945
rect 58161 58905 58173 58939
rect 58207 58936 58219 58939
rect 58894 58936 58900 58948
rect 58207 58908 58900 58936
rect 58207 58905 58219 58908
rect 58161 58899 58219 58905
rect 1765 58871 1823 58877
rect 1765 58837 1777 58871
rect 1811 58868 1823 58871
rect 18506 58868 18512 58880
rect 1811 58840 18512 58868
rect 1811 58837 1823 58840
rect 1765 58831 1823 58837
rect 18506 58828 18512 58840
rect 18564 58828 18570 58880
rect 19628 58868 19656 58899
rect 58894 58896 58900 58908
rect 58952 58896 58958 58948
rect 20070 58868 20076 58880
rect 19628 58840 20076 58868
rect 20070 58828 20076 58840
rect 20128 58828 20134 58880
rect 41138 58828 41144 58880
rect 41196 58828 41202 58880
rect 1104 58778 58880 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 58880 58778
rect 1104 58704 58880 58726
rect 2038 58624 2044 58676
rect 2096 58664 2102 58676
rect 2096 58636 41368 58664
rect 2096 58624 2102 58636
rect 934 58488 940 58540
rect 992 58528 998 58540
rect 1581 58531 1639 58537
rect 1581 58528 1593 58531
rect 992 58500 1593 58528
rect 992 58488 998 58500
rect 1581 58497 1593 58500
rect 1627 58497 1639 58531
rect 1581 58491 1639 58497
rect 34514 58488 34520 58540
rect 34572 58528 34578 58540
rect 35713 58531 35771 58537
rect 35713 58528 35725 58531
rect 34572 58500 35725 58528
rect 34572 58488 34578 58500
rect 35713 58497 35725 58500
rect 35759 58497 35771 58531
rect 37918 58528 37924 58540
rect 35713 58491 35771 58497
rect 36004 58500 37924 58528
rect 1857 58463 1915 58469
rect 1857 58429 1869 58463
rect 1903 58460 1915 58463
rect 3418 58460 3424 58472
rect 1903 58432 3424 58460
rect 1903 58429 1915 58432
rect 1857 58423 1915 58429
rect 3418 58420 3424 58432
rect 3476 58420 3482 58472
rect 35802 58420 35808 58472
rect 35860 58460 35866 58472
rect 36004 58469 36032 58500
rect 37918 58488 37924 58500
rect 37976 58488 37982 58540
rect 38194 58488 38200 58540
rect 38252 58488 38258 58540
rect 38286 58488 38292 58540
rect 38344 58488 38350 58540
rect 38470 58488 38476 58540
rect 38528 58528 38534 58540
rect 38565 58531 38623 58537
rect 38565 58528 38577 58531
rect 38528 58500 38577 58528
rect 38528 58488 38534 58500
rect 38565 58497 38577 58500
rect 38611 58497 38623 58531
rect 38565 58491 38623 58497
rect 38838 58488 38844 58540
rect 38896 58488 38902 58540
rect 41340 58537 41368 58636
rect 58158 58556 58164 58608
rect 58216 58556 58222 58608
rect 41325 58531 41383 58537
rect 41325 58497 41337 58531
rect 41371 58497 41383 58531
rect 41325 58491 41383 58497
rect 41509 58531 41567 58537
rect 41509 58497 41521 58531
rect 41555 58497 41567 58531
rect 41509 58491 41567 58497
rect 41877 58531 41935 58537
rect 41877 58497 41889 58531
rect 41923 58528 41935 58531
rect 49694 58528 49700 58540
rect 41923 58500 49700 58528
rect 41923 58497 41935 58500
rect 41877 58491 41935 58497
rect 35989 58463 36047 58469
rect 35989 58460 36001 58463
rect 35860 58432 36001 58460
rect 35860 58420 35866 58432
rect 35989 58429 36001 58432
rect 36035 58429 36047 58463
rect 35989 58423 36047 58429
rect 40034 58420 40040 58472
rect 40092 58460 40098 58472
rect 41524 58460 41552 58491
rect 49694 58488 49700 58500
rect 49752 58488 49758 58540
rect 40092 58432 41552 58460
rect 41785 58463 41843 58469
rect 40092 58420 40098 58432
rect 41785 58429 41797 58463
rect 41831 58429 41843 58463
rect 41785 58423 41843 58429
rect 36906 58352 36912 58404
rect 36964 58392 36970 58404
rect 38286 58392 38292 58404
rect 36964 58364 38292 58392
rect 36964 58352 36970 58364
rect 38286 58352 38292 58364
rect 38344 58352 38350 58404
rect 41598 58392 41604 58404
rect 38626 58364 41604 58392
rect 37550 58284 37556 58336
rect 37608 58284 37614 58336
rect 37918 58284 37924 58336
rect 37976 58324 37982 58336
rect 38626 58324 38654 58364
rect 41598 58352 41604 58364
rect 41656 58392 41662 58404
rect 41800 58392 41828 58423
rect 41656 58364 41828 58392
rect 41656 58352 41662 58364
rect 37976 58296 38654 58324
rect 41141 58327 41199 58333
rect 37976 58284 37982 58296
rect 41141 58293 41153 58327
rect 41187 58324 41199 58327
rect 42610 58324 42616 58336
rect 41187 58296 42616 58324
rect 41187 58293 41199 58296
rect 41141 58287 41199 58293
rect 42610 58284 42616 58296
rect 42668 58284 42674 58336
rect 58250 58284 58256 58336
rect 58308 58284 58314 58336
rect 1104 58234 58880 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 58880 58234
rect 1104 58160 58880 58182
rect 35802 57984 35808 57996
rect 35636 57956 35808 57984
rect 934 57876 940 57928
rect 992 57916 998 57928
rect 35636 57925 35664 57956
rect 35802 57944 35808 57956
rect 35860 57944 35866 57996
rect 1581 57919 1639 57925
rect 1581 57916 1593 57919
rect 992 57888 1593 57916
rect 992 57876 998 57888
rect 1581 57885 1593 57888
rect 1627 57885 1639 57919
rect 1581 57879 1639 57885
rect 35621 57919 35679 57925
rect 35621 57885 35633 57919
rect 35667 57885 35679 57919
rect 35621 57879 35679 57885
rect 35710 57876 35716 57928
rect 35768 57876 35774 57928
rect 35989 57919 36047 57925
rect 35989 57885 36001 57919
rect 36035 57885 36047 57919
rect 35989 57879 36047 57885
rect 1857 57851 1915 57857
rect 1857 57817 1869 57851
rect 1903 57848 1915 57851
rect 5994 57848 6000 57860
rect 1903 57820 6000 57848
rect 1903 57817 1915 57820
rect 1857 57811 1915 57817
rect 5994 57808 6000 57820
rect 6052 57808 6058 57860
rect 34790 57808 34796 57860
rect 34848 57848 34854 57860
rect 35161 57851 35219 57857
rect 35161 57848 35173 57851
rect 34848 57820 35173 57848
rect 34848 57808 34854 57820
rect 35161 57817 35173 57820
rect 35207 57817 35219 57851
rect 35161 57811 35219 57817
rect 35434 57740 35440 57792
rect 35492 57780 35498 57792
rect 36004 57780 36032 57879
rect 36262 57876 36268 57928
rect 36320 57876 36326 57928
rect 36541 57919 36599 57925
rect 36541 57885 36553 57919
rect 36587 57916 36599 57919
rect 58250 57916 58256 57928
rect 36587 57888 58256 57916
rect 36587 57885 36599 57888
rect 36541 57879 36599 57885
rect 58250 57876 58256 57888
rect 58308 57876 58314 57928
rect 57974 57808 57980 57860
rect 58032 57808 58038 57860
rect 35492 57752 36032 57780
rect 35492 57740 35498 57752
rect 58066 57740 58072 57792
rect 58124 57740 58130 57792
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 934 57400 940 57452
rect 992 57440 998 57452
rect 1581 57443 1639 57449
rect 1581 57440 1593 57443
rect 992 57412 1593 57440
rect 992 57400 998 57412
rect 1581 57409 1593 57412
rect 1627 57409 1639 57443
rect 1581 57403 1639 57409
rect 1762 57196 1768 57248
rect 1820 57196 1826 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 33410 56992 33416 57044
rect 33468 57032 33474 57044
rect 33468 57004 38654 57032
rect 33468 56992 33474 57004
rect 24854 56924 24860 56976
rect 24912 56964 24918 56976
rect 36262 56964 36268 56976
rect 24912 56936 36268 56964
rect 24912 56924 24918 56936
rect 33336 56905 33364 56936
rect 36262 56924 36268 56936
rect 36320 56924 36326 56976
rect 33321 56899 33379 56905
rect 33321 56865 33333 56899
rect 33367 56865 33379 56899
rect 38626 56896 38654 57004
rect 41138 56992 41144 57044
rect 41196 57032 41202 57044
rect 43254 57032 43260 57044
rect 41196 57004 43260 57032
rect 41196 56992 41202 57004
rect 43254 56992 43260 57004
rect 43312 56992 43318 57044
rect 56502 56964 56508 56976
rect 41386 56936 56508 56964
rect 41386 56896 41414 56936
rect 56502 56924 56508 56936
rect 56560 56924 56566 56976
rect 38626 56868 41414 56896
rect 33321 56859 33379 56865
rect 22462 56788 22468 56840
rect 22520 56828 22526 56840
rect 32861 56831 32919 56837
rect 32861 56828 32873 56831
rect 22520 56800 32873 56828
rect 22520 56788 22526 56800
rect 32861 56797 32873 56800
rect 32907 56797 32919 56831
rect 32861 56791 32919 56797
rect 33042 56788 33048 56840
rect 33100 56788 33106 56840
rect 33410 56788 33416 56840
rect 33468 56788 33474 56840
rect 57885 56831 57943 56837
rect 57885 56797 57897 56831
rect 57931 56828 57943 56831
rect 58986 56828 58992 56840
rect 57931 56800 58992 56828
rect 57931 56797 57943 56800
rect 57885 56791 57943 56797
rect 58986 56788 58992 56800
rect 59044 56788 59050 56840
rect 934 56720 940 56772
rect 992 56760 998 56772
rect 1673 56763 1731 56769
rect 1673 56760 1685 56763
rect 992 56732 1685 56760
rect 992 56720 998 56732
rect 1673 56729 1685 56732
rect 1719 56729 1731 56763
rect 41414 56760 41420 56772
rect 1673 56723 1731 56729
rect 22066 56732 41420 56760
rect 1949 56695 2007 56701
rect 1949 56661 1961 56695
rect 1995 56692 2007 56695
rect 22066 56692 22094 56732
rect 41414 56720 41420 56732
rect 41472 56720 41478 56772
rect 55858 56720 55864 56772
rect 55916 56760 55922 56772
rect 58161 56763 58219 56769
rect 58161 56760 58173 56763
rect 55916 56732 58173 56760
rect 55916 56720 55922 56732
rect 58161 56729 58173 56732
rect 58207 56729 58219 56763
rect 58161 56723 58219 56729
rect 1995 56664 22094 56692
rect 1995 56661 2007 56664
rect 1949 56655 2007 56661
rect 32674 56652 32680 56704
rect 32732 56652 32738 56704
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 56502 56448 56508 56500
rect 56560 56488 56566 56500
rect 58253 56491 58311 56497
rect 58253 56488 58265 56491
rect 56560 56460 58265 56488
rect 56560 56448 56566 56460
rect 58253 56457 58265 56460
rect 58299 56457 58311 56491
rect 58253 56451 58311 56457
rect 58161 56423 58219 56429
rect 58161 56389 58173 56423
rect 58207 56420 58219 56423
rect 58986 56420 58992 56432
rect 58207 56392 58992 56420
rect 58207 56389 58219 56392
rect 58161 56383 58219 56389
rect 58986 56380 58992 56392
rect 59044 56380 59050 56432
rect 41506 56312 41512 56364
rect 41564 56312 41570 56364
rect 41877 56355 41935 56361
rect 41877 56321 41889 56355
rect 41923 56352 41935 56355
rect 46842 56352 46848 56364
rect 41923 56324 46848 56352
rect 41923 56321 41935 56324
rect 41877 56315 41935 56321
rect 46842 56312 46848 56324
rect 46900 56312 46906 56364
rect 41414 56244 41420 56296
rect 41472 56244 41478 56296
rect 41785 56287 41843 56293
rect 41785 56253 41797 56287
rect 41831 56253 41843 56287
rect 41785 56247 41843 56253
rect 41230 56176 41236 56228
rect 41288 56216 41294 56228
rect 41598 56216 41604 56228
rect 41288 56188 41604 56216
rect 41288 56176 41294 56188
rect 41598 56176 41604 56188
rect 41656 56216 41662 56228
rect 41800 56216 41828 56247
rect 41656 56188 41828 56216
rect 41656 56176 41662 56188
rect 41141 56151 41199 56157
rect 41141 56117 41153 56151
rect 41187 56148 41199 56151
rect 41322 56148 41328 56160
rect 41187 56120 41328 56148
rect 41187 56117 41199 56120
rect 41141 56111 41199 56117
rect 41322 56108 41328 56120
rect 41380 56108 41386 56160
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 23566 55904 23572 55956
rect 23624 55944 23630 55956
rect 30466 55944 30472 55956
rect 23624 55916 30472 55944
rect 23624 55904 23630 55916
rect 30466 55904 30472 55916
rect 30524 55904 30530 55956
rect 58342 55904 58348 55956
rect 58400 55904 58406 55956
rect 1762 55836 1768 55888
rect 1820 55876 1826 55888
rect 1820 55848 30788 55876
rect 1820 55836 1826 55848
rect 24118 55768 24124 55820
rect 24176 55808 24182 55820
rect 25133 55811 25191 55817
rect 25133 55808 25145 55811
rect 24176 55780 25145 55808
rect 24176 55768 24182 55780
rect 25133 55777 25145 55780
rect 25179 55777 25191 55811
rect 30558 55808 30564 55820
rect 25133 55771 25191 55777
rect 25240 55780 30564 55808
rect 25240 55749 25268 55780
rect 30558 55768 30564 55780
rect 30616 55768 30622 55820
rect 25225 55743 25283 55749
rect 25225 55709 25237 55743
rect 25271 55709 25283 55743
rect 25225 55703 25283 55709
rect 25593 55743 25651 55749
rect 25593 55709 25605 55743
rect 25639 55709 25651 55743
rect 25593 55703 25651 55709
rect 934 55632 940 55684
rect 992 55672 998 55684
rect 1673 55675 1731 55681
rect 1673 55672 1685 55675
rect 992 55644 1685 55672
rect 992 55632 998 55644
rect 1673 55641 1685 55644
rect 1719 55641 1731 55675
rect 1673 55635 1731 55641
rect 24578 55632 24584 55684
rect 24636 55632 24642 55684
rect 1765 55607 1823 55613
rect 1765 55573 1777 55607
rect 1811 55604 1823 55607
rect 25608 55604 25636 55703
rect 25682 55700 25688 55752
rect 25740 55740 25746 55752
rect 25740 55712 30328 55740
rect 25740 55700 25746 55712
rect 29730 55632 29736 55684
rect 29788 55632 29794 55684
rect 30300 55672 30328 55712
rect 30374 55700 30380 55752
rect 30432 55700 30438 55752
rect 30466 55700 30472 55752
rect 30524 55700 30530 55752
rect 30760 55749 30788 55848
rect 30745 55743 30803 55749
rect 30745 55709 30757 55743
rect 30791 55709 30803 55743
rect 30745 55703 30803 55709
rect 30837 55743 30895 55749
rect 30837 55709 30849 55743
rect 30883 55740 30895 55743
rect 40034 55740 40040 55752
rect 30883 55712 40040 55740
rect 30883 55709 30895 55712
rect 30837 55703 30895 55709
rect 30852 55672 30880 55703
rect 40034 55700 40040 55712
rect 40092 55700 40098 55752
rect 30300 55644 30880 55672
rect 1811 55576 25636 55604
rect 1811 55573 1823 55576
rect 1765 55567 1823 55573
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 1765 55403 1823 55409
rect 1765 55369 1777 55403
rect 1811 55400 1823 55403
rect 1811 55372 6914 55400
rect 1811 55369 1823 55372
rect 1765 55363 1823 55369
rect 6886 55332 6914 55372
rect 24302 55360 24308 55412
rect 24360 55400 24366 55412
rect 25682 55400 25688 55412
rect 24360 55372 25688 55400
rect 24360 55360 24366 55372
rect 25682 55360 25688 55372
rect 25740 55360 25746 55412
rect 41506 55400 41512 55412
rect 41064 55372 41512 55400
rect 6886 55304 31754 55332
rect 934 55224 940 55276
rect 992 55264 998 55276
rect 1581 55267 1639 55273
rect 1581 55264 1593 55267
rect 992 55236 1593 55264
rect 992 55224 998 55236
rect 1581 55233 1593 55236
rect 1627 55233 1639 55267
rect 1581 55227 1639 55233
rect 23753 55267 23811 55273
rect 23753 55233 23765 55267
rect 23799 55264 23811 55267
rect 23934 55264 23940 55276
rect 23799 55236 23940 55264
rect 23799 55233 23811 55236
rect 23753 55227 23811 55233
rect 23934 55224 23940 55236
rect 23992 55224 23998 55276
rect 24026 55224 24032 55276
rect 24084 55264 24090 55276
rect 24084 55236 24348 55264
rect 24084 55224 24090 55236
rect 24320 55205 24348 55236
rect 24394 55224 24400 55276
rect 24452 55224 24458 55276
rect 24762 55224 24768 55276
rect 24820 55224 24826 55276
rect 24946 55224 24952 55276
rect 25004 55264 25010 55276
rect 25314 55264 25320 55276
rect 25004 55236 25320 55264
rect 25004 55224 25010 55236
rect 25314 55224 25320 55236
rect 25372 55224 25378 55276
rect 31726 55264 31754 55304
rect 41064 55276 41092 55372
rect 41506 55360 41512 55372
rect 41564 55360 41570 55412
rect 41141 55335 41199 55341
rect 41141 55301 41153 55335
rect 41187 55332 41199 55335
rect 44174 55332 44180 55344
rect 41187 55304 44180 55332
rect 41187 55301 41199 55304
rect 41141 55295 41199 55301
rect 44174 55292 44180 55304
rect 44232 55292 44238 55344
rect 40865 55267 40923 55273
rect 40865 55264 40877 55267
rect 31726 55236 40877 55264
rect 40865 55233 40877 55236
rect 40911 55233 40923 55267
rect 40865 55227 40923 55233
rect 41046 55224 41052 55276
rect 41104 55224 41110 55276
rect 41230 55224 41236 55276
rect 41288 55273 41294 55276
rect 41288 55264 41296 55273
rect 41434 55267 41492 55273
rect 41288 55236 41333 55264
rect 41288 55227 41296 55236
rect 41434 55233 41446 55267
rect 41480 55264 41492 55267
rect 42058 55264 42064 55276
rect 41480 55236 42064 55264
rect 41480 55233 41492 55236
rect 41434 55227 41492 55233
rect 41288 55224 41294 55227
rect 42058 55224 42064 55236
rect 42116 55224 42122 55276
rect 24305 55199 24363 55205
rect 24305 55165 24317 55199
rect 24351 55165 24363 55199
rect 24305 55159 24363 55165
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 28718 54720 28724 54732
rect 23492 54692 28724 54720
rect 23492 54661 23520 54692
rect 28718 54680 28724 54692
rect 28776 54680 28782 54732
rect 23477 54655 23535 54661
rect 23477 54621 23489 54655
rect 23523 54621 23535 54655
rect 23477 54615 23535 54621
rect 23566 54612 23572 54664
rect 23624 54612 23630 54664
rect 23845 54655 23903 54661
rect 23845 54621 23857 54655
rect 23891 54621 23903 54655
rect 23845 54615 23903 54621
rect 24029 54655 24087 54661
rect 24029 54621 24041 54655
rect 24075 54652 24087 54655
rect 24302 54652 24308 54664
rect 24075 54624 24308 54652
rect 24075 54621 24087 54624
rect 24029 54615 24087 54621
rect 934 54544 940 54596
rect 992 54584 998 54596
rect 1673 54587 1731 54593
rect 1673 54584 1685 54587
rect 992 54556 1685 54584
rect 992 54544 998 54556
rect 1673 54553 1685 54556
rect 1719 54553 1731 54587
rect 1673 54547 1731 54553
rect 22094 54544 22100 54596
rect 22152 54584 22158 54596
rect 22833 54587 22891 54593
rect 22833 54584 22845 54587
rect 22152 54556 22845 54584
rect 22152 54544 22158 54556
rect 22833 54553 22845 54556
rect 22879 54553 22891 54587
rect 22833 54547 22891 54553
rect 1765 54519 1823 54525
rect 1765 54485 1777 54519
rect 1811 54516 1823 54519
rect 23860 54516 23888 54615
rect 24302 54612 24308 54624
rect 24360 54612 24366 54664
rect 58342 54612 58348 54664
rect 58400 54612 58406 54664
rect 1811 54488 23888 54516
rect 1811 54485 1823 54488
rect 1765 54479 1823 54485
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 934 54136 940 54188
rect 992 54176 998 54188
rect 1581 54179 1639 54185
rect 1581 54176 1593 54179
rect 992 54148 1593 54176
rect 992 54136 998 54148
rect 1581 54145 1593 54148
rect 1627 54145 1639 54179
rect 1581 54139 1639 54145
rect 1762 53932 1768 53984
rect 1820 53932 1826 53984
rect 23566 53932 23572 53984
rect 23624 53972 23630 53984
rect 24210 53972 24216 53984
rect 23624 53944 24216 53972
rect 23624 53932 23630 53944
rect 24210 53932 24216 53944
rect 24268 53932 24274 53984
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 40126 53660 40132 53712
rect 40184 53700 40190 53712
rect 40957 53703 41015 53709
rect 40957 53700 40969 53703
rect 40184 53672 40969 53700
rect 40184 53660 40190 53672
rect 40957 53669 40969 53672
rect 41003 53669 41015 53703
rect 40957 53663 41015 53669
rect 24946 53592 24952 53644
rect 25004 53632 25010 53644
rect 41046 53632 41052 53644
rect 25004 53604 41052 53632
rect 25004 53592 25010 53604
rect 40604 53573 40632 53604
rect 41046 53592 41052 53604
rect 41104 53592 41110 53644
rect 40405 53567 40463 53573
rect 40405 53564 40417 53567
rect 40052 53536 40417 53564
rect 21266 53456 21272 53508
rect 21324 53496 21330 53508
rect 24394 53496 24400 53508
rect 21324 53468 24400 53496
rect 21324 53456 21330 53468
rect 24394 53456 24400 53468
rect 24452 53456 24458 53508
rect 1762 53388 1768 53440
rect 1820 53428 1826 53440
rect 40052 53437 40080 53536
rect 40405 53533 40417 53536
rect 40451 53533 40463 53567
rect 40405 53527 40463 53533
rect 40589 53567 40647 53573
rect 40589 53533 40601 53567
rect 40635 53533 40647 53567
rect 40589 53527 40647 53533
rect 40825 53567 40883 53573
rect 40825 53533 40837 53567
rect 40871 53564 40883 53567
rect 41230 53564 41236 53576
rect 40871 53536 41236 53564
rect 40871 53533 40883 53536
rect 40825 53527 40883 53533
rect 41230 53524 41236 53536
rect 41288 53524 41294 53576
rect 40681 53499 40739 53505
rect 40681 53465 40693 53499
rect 40727 53496 40739 53499
rect 44818 53496 44824 53508
rect 40727 53468 44824 53496
rect 40727 53465 40739 53468
rect 40681 53459 40739 53465
rect 44818 53456 44824 53468
rect 44876 53456 44882 53508
rect 40037 53431 40095 53437
rect 40037 53428 40049 53431
rect 1820 53400 40049 53428
rect 1820 53388 1826 53400
rect 40037 53397 40049 53400
rect 40083 53397 40095 53431
rect 40037 53391 40095 53397
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 24946 53224 24952 53236
rect 23768 53196 24952 53224
rect 23768 53165 23796 53196
rect 24946 53184 24952 53196
rect 25004 53184 25010 53236
rect 23753 53159 23811 53165
rect 23753 53125 23765 53159
rect 23799 53125 23811 53159
rect 23753 53119 23811 53125
rect 23845 53159 23903 53165
rect 23845 53125 23857 53159
rect 23891 53156 23903 53159
rect 23891 53128 31754 53156
rect 23891 53125 23903 53128
rect 23845 53119 23903 53125
rect 934 53048 940 53100
rect 992 53088 998 53100
rect 1673 53091 1731 53097
rect 1673 53088 1685 53091
rect 992 53060 1685 53088
rect 992 53048 998 53060
rect 1673 53057 1685 53060
rect 1719 53057 1731 53091
rect 23569 53091 23627 53097
rect 23569 53088 23581 53091
rect 1673 53051 1731 53057
rect 6886 53060 23581 53088
rect 1765 52887 1823 52893
rect 1765 52853 1777 52887
rect 1811 52884 1823 52887
rect 6886 52884 6914 53060
rect 23569 53057 23581 53060
rect 23615 53057 23627 53091
rect 23569 53051 23627 53057
rect 23658 53048 23664 53100
rect 23716 53088 23722 53100
rect 23937 53091 23995 53097
rect 23937 53088 23949 53091
rect 23716 53060 23949 53088
rect 23716 53048 23722 53060
rect 23937 53057 23949 53060
rect 23983 53057 23995 53091
rect 23937 53051 23995 53057
rect 23952 53020 23980 53051
rect 24394 53048 24400 53100
rect 24452 53088 24458 53100
rect 24581 53091 24639 53097
rect 24581 53088 24593 53091
rect 24452 53060 24593 53088
rect 24452 53048 24458 53060
rect 24581 53057 24593 53060
rect 24627 53057 24639 53091
rect 31726 53088 31754 53128
rect 45370 53088 45376 53100
rect 31726 53060 45376 53088
rect 24581 53051 24639 53057
rect 45370 53048 45376 53060
rect 45428 53048 45434 53100
rect 24765 53023 24823 53029
rect 24765 53020 24777 53023
rect 23952 52992 24777 53020
rect 24765 52989 24777 52992
rect 24811 52989 24823 53023
rect 24765 52983 24823 52989
rect 1811 52856 6914 52884
rect 1811 52853 1823 52856
rect 1765 52847 1823 52853
rect 23842 52844 23848 52896
rect 23900 52884 23906 52896
rect 24121 52887 24179 52893
rect 24121 52884 24133 52887
rect 23900 52856 24133 52884
rect 23900 52844 23906 52856
rect 24121 52853 24133 52856
rect 24167 52853 24179 52887
rect 24121 52847 24179 52853
rect 58342 52844 58348 52896
rect 58400 52844 58406 52896
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 24946 52640 24952 52692
rect 25004 52640 25010 52692
rect 2038 52436 2044 52488
rect 2096 52436 2102 52488
rect 934 52368 940 52420
rect 992 52408 998 52420
rect 1673 52411 1731 52417
rect 1673 52408 1685 52411
rect 992 52380 1685 52408
rect 992 52368 998 52380
rect 1673 52377 1685 52380
rect 1719 52377 1731 52411
rect 1673 52371 1731 52377
rect 21450 52368 21456 52420
rect 21508 52408 21514 52420
rect 24673 52411 24731 52417
rect 24673 52408 24685 52411
rect 21508 52380 24685 52408
rect 21508 52368 21514 52380
rect 24673 52377 24685 52380
rect 24719 52377 24731 52411
rect 24673 52371 24731 52377
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 20254 52096 20260 52148
rect 20312 52136 20318 52148
rect 21177 52139 21235 52145
rect 21177 52136 21189 52139
rect 20312 52108 21189 52136
rect 20312 52096 20318 52108
rect 21177 52105 21189 52108
rect 21223 52105 21235 52139
rect 21177 52099 21235 52105
rect 1857 52071 1915 52077
rect 1857 52037 1869 52071
rect 1903 52068 1915 52071
rect 8205 52071 8263 52077
rect 8205 52068 8217 52071
rect 1903 52040 8217 52068
rect 1903 52037 1915 52040
rect 1857 52031 1915 52037
rect 8205 52037 8217 52040
rect 8251 52037 8263 52071
rect 8205 52031 8263 52037
rect 934 51960 940 52012
rect 992 52000 998 52012
rect 1673 52003 1731 52009
rect 1673 52000 1685 52003
rect 992 51972 1685 52000
rect 992 51960 998 51972
rect 1673 51969 1685 51972
rect 1719 51969 1731 52003
rect 1673 51963 1731 51969
rect 8018 51960 8024 52012
rect 8076 51960 8082 52012
rect 8294 51960 8300 52012
rect 8352 51960 8358 52012
rect 21269 52003 21327 52009
rect 21269 51969 21281 52003
rect 21315 52000 21327 52003
rect 22186 52000 22192 52012
rect 21315 51972 22192 52000
rect 21315 51969 21327 51972
rect 21269 51963 21327 51969
rect 22186 51960 22192 51972
rect 22244 52000 22250 52012
rect 22830 52000 22836 52012
rect 22244 51972 22836 52000
rect 22244 51960 22250 51972
rect 22830 51960 22836 51972
rect 22888 51960 22894 52012
rect 17862 51892 17868 51944
rect 17920 51932 17926 51944
rect 20993 51935 21051 51941
rect 20993 51932 21005 51935
rect 17920 51904 21005 51932
rect 17920 51892 17926 51904
rect 20993 51901 21005 51904
rect 21039 51901 21051 51935
rect 20993 51895 21051 51901
rect 20901 51867 20959 51873
rect 20901 51833 20913 51867
rect 20947 51864 20959 51867
rect 20947 51836 31754 51864
rect 20947 51833 20959 51836
rect 20901 51827 20959 51833
rect 7834 51756 7840 51808
rect 7892 51756 7898 51808
rect 20530 51756 20536 51808
rect 20588 51756 20594 51808
rect 20809 51799 20867 51805
rect 20809 51765 20821 51799
rect 20855 51796 20867 51799
rect 24210 51796 24216 51808
rect 20855 51768 24216 51796
rect 20855 51765 20867 51768
rect 20809 51759 20867 51765
rect 24210 51756 24216 51768
rect 24268 51756 24274 51808
rect 31726 51796 31754 51836
rect 41138 51796 41144 51808
rect 31726 51768 41144 51796
rect 41138 51756 41144 51768
rect 41196 51756 41202 51808
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 58342 51348 58348 51400
rect 58400 51348 58406 51400
rect 934 51280 940 51332
rect 992 51320 998 51332
rect 1673 51323 1731 51329
rect 1673 51320 1685 51323
rect 992 51292 1685 51320
rect 992 51280 998 51292
rect 1673 51289 1685 51292
rect 1719 51289 1731 51323
rect 1673 51283 1731 51289
rect 1857 51323 1915 51329
rect 1857 51289 1869 51323
rect 1903 51320 1915 51323
rect 3970 51320 3976 51332
rect 1903 51292 3976 51320
rect 1903 51289 1915 51292
rect 1857 51283 1915 51289
rect 3970 51280 3976 51292
rect 4028 51280 4034 51332
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 2682 50940 2688 50992
rect 2740 50980 2746 50992
rect 3881 50983 3939 50989
rect 3881 50980 3893 50983
rect 2740 50952 3893 50980
rect 2740 50940 2746 50952
rect 3881 50949 3893 50952
rect 3927 50949 3939 50983
rect 3881 50943 3939 50949
rect 3970 50940 3976 50992
rect 4028 50940 4034 50992
rect 3697 50915 3755 50921
rect 3697 50881 3709 50915
rect 3743 50881 3755 50915
rect 3697 50875 3755 50881
rect 3712 50844 3740 50875
rect 4062 50872 4068 50924
rect 4120 50921 4126 50924
rect 4120 50912 4128 50921
rect 4120 50884 4165 50912
rect 4120 50875 4128 50884
rect 4120 50872 4126 50875
rect 4614 50844 4620 50856
rect 3712 50816 4620 50844
rect 4614 50804 4620 50816
rect 4672 50804 4678 50856
rect 4249 50711 4307 50717
rect 4249 50677 4261 50711
rect 4295 50708 4307 50711
rect 6270 50708 6276 50720
rect 4295 50680 6276 50708
rect 4295 50677 4307 50680
rect 4249 50671 4307 50677
rect 6270 50668 6276 50680
rect 6328 50668 6334 50720
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 27338 50396 27344 50448
rect 27396 50436 27402 50448
rect 40770 50436 40776 50448
rect 27396 50408 40776 50436
rect 27396 50396 27402 50408
rect 40770 50396 40776 50408
rect 40828 50396 40834 50448
rect 5994 50328 6000 50380
rect 6052 50368 6058 50380
rect 29546 50368 29552 50380
rect 6052 50340 29552 50368
rect 6052 50328 6058 50340
rect 29546 50328 29552 50340
rect 29604 50328 29610 50380
rect 32674 50328 32680 50380
rect 32732 50368 32738 50380
rect 33226 50368 33232 50380
rect 32732 50340 33232 50368
rect 32732 50328 32738 50340
rect 33226 50328 33232 50340
rect 33284 50328 33290 50380
rect 36538 50328 36544 50380
rect 36596 50368 36602 50380
rect 56594 50368 56600 50380
rect 36596 50340 56600 50368
rect 36596 50328 36602 50340
rect 56594 50328 56600 50340
rect 56652 50328 56658 50380
rect 57514 50260 57520 50312
rect 57572 50300 57578 50312
rect 57885 50303 57943 50309
rect 57885 50300 57897 50303
rect 57572 50272 57897 50300
rect 57572 50260 57578 50272
rect 57885 50269 57897 50272
rect 57931 50269 57943 50303
rect 57885 50263 57943 50269
rect 934 50192 940 50244
rect 992 50232 998 50244
rect 1673 50235 1731 50241
rect 1673 50232 1685 50235
rect 992 50204 1685 50232
rect 992 50192 998 50204
rect 1673 50201 1685 50204
rect 1719 50201 1731 50235
rect 1673 50195 1731 50201
rect 1857 50235 1915 50241
rect 1857 50201 1869 50235
rect 1903 50232 1915 50235
rect 2038 50232 2044 50244
rect 1903 50204 2044 50232
rect 1903 50201 1915 50204
rect 1857 50195 1915 50201
rect 2038 50192 2044 50204
rect 2096 50192 2102 50244
rect 58161 50235 58219 50241
rect 58161 50201 58173 50235
rect 58207 50232 58219 50235
rect 58986 50232 58992 50244
rect 58207 50204 58992 50232
rect 58207 50201 58219 50204
rect 58161 50195 58219 50201
rect 58986 50192 58992 50204
rect 59044 50192 59050 50244
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 934 49784 940 49836
rect 992 49824 998 49836
rect 1581 49827 1639 49833
rect 1581 49824 1593 49827
rect 992 49796 1593 49824
rect 992 49784 998 49796
rect 1581 49793 1593 49796
rect 1627 49793 1639 49827
rect 1581 49787 1639 49793
rect 4062 49784 4068 49836
rect 4120 49824 4126 49836
rect 6822 49824 6828 49836
rect 4120 49796 6828 49824
rect 4120 49784 4126 49796
rect 6822 49784 6828 49796
rect 6880 49824 6886 49836
rect 8294 49824 8300 49836
rect 6880 49796 8300 49824
rect 6880 49784 6886 49796
rect 8294 49784 8300 49796
rect 8352 49784 8358 49836
rect 13078 49756 13084 49768
rect 1780 49728 13084 49756
rect 1780 49697 1808 49728
rect 13078 49716 13084 49728
rect 13136 49716 13142 49768
rect 1765 49691 1823 49697
rect 1765 49657 1777 49691
rect 1811 49657 1823 49691
rect 1765 49651 1823 49657
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 934 49172 940 49224
rect 992 49212 998 49224
rect 1581 49215 1639 49221
rect 1581 49212 1593 49215
rect 992 49184 1593 49212
rect 992 49172 998 49184
rect 1581 49181 1593 49184
rect 1627 49181 1639 49215
rect 1581 49175 1639 49181
rect 57974 49104 57980 49156
rect 58032 49104 58038 49156
rect 58345 49147 58403 49153
rect 58345 49113 58357 49147
rect 58391 49144 58403 49147
rect 59446 49144 59452 49156
rect 58391 49116 59452 49144
rect 58391 49113 58403 49116
rect 58345 49107 58403 49113
rect 59446 49104 59452 49116
rect 59504 49104 59510 49156
rect 1765 49079 1823 49085
rect 1765 49045 1777 49079
rect 1811 49076 1823 49079
rect 6454 49076 6460 49088
rect 1811 49048 6460 49076
rect 1811 49045 1823 49048
rect 1765 49039 1823 49045
rect 6454 49036 6460 49048
rect 6512 49036 6518 49088
rect 25406 49036 25412 49088
rect 25464 49076 25470 49088
rect 43070 49076 43076 49088
rect 25464 49048 43076 49076
rect 25464 49036 25470 49048
rect 43070 49036 43076 49048
rect 43128 49036 43134 49088
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 934 48696 940 48748
rect 992 48736 998 48748
rect 1673 48739 1731 48745
rect 1673 48736 1685 48739
rect 992 48708 1685 48736
rect 992 48696 998 48708
rect 1673 48705 1685 48708
rect 1719 48705 1731 48739
rect 1673 48699 1731 48705
rect 1857 48603 1915 48609
rect 1857 48569 1869 48603
rect 1903 48600 1915 48603
rect 1946 48600 1952 48612
rect 1903 48572 1952 48600
rect 1903 48569 1915 48572
rect 1857 48563 1915 48569
rect 1946 48560 1952 48572
rect 2004 48560 2010 48612
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 2593 48263 2651 48269
rect 2593 48229 2605 48263
rect 2639 48260 2651 48263
rect 17862 48260 17868 48272
rect 2639 48232 17868 48260
rect 2639 48229 2651 48232
rect 2593 48223 2651 48229
rect 17862 48220 17868 48232
rect 17920 48220 17926 48272
rect 55950 48220 55956 48272
rect 56008 48260 56014 48272
rect 58066 48260 58072 48272
rect 56008 48232 58072 48260
rect 56008 48220 56014 48232
rect 58066 48220 58072 48232
rect 58124 48220 58130 48272
rect 4062 48192 4068 48204
rect 2240 48164 4068 48192
rect 2038 48084 2044 48136
rect 2096 48084 2102 48136
rect 2240 48133 2268 48164
rect 4062 48152 4068 48164
rect 4120 48152 4126 48204
rect 6822 48152 6828 48204
rect 6880 48192 6886 48204
rect 9030 48192 9036 48204
rect 6880 48164 9036 48192
rect 6880 48152 6886 48164
rect 9030 48152 9036 48164
rect 9088 48152 9094 48204
rect 2225 48127 2283 48133
rect 2225 48093 2237 48127
rect 2271 48093 2283 48127
rect 2225 48087 2283 48093
rect 2406 48084 2412 48136
rect 2464 48133 2470 48136
rect 2464 48087 2472 48133
rect 2464 48084 2470 48087
rect 57790 48084 57796 48136
rect 57848 48124 57854 48136
rect 57885 48127 57943 48133
rect 57885 48124 57897 48127
rect 57848 48096 57897 48124
rect 57848 48084 57854 48096
rect 57885 48093 57897 48096
rect 57931 48093 57943 48127
rect 57885 48087 57943 48093
rect 2317 48059 2375 48065
rect 2317 48025 2329 48059
rect 2363 48025 2375 48059
rect 2317 48019 2375 48025
rect 1578 47948 1584 48000
rect 1636 47988 1642 48000
rect 2332 47988 2360 48019
rect 58158 48016 58164 48068
rect 58216 48016 58222 48068
rect 1636 47960 2360 47988
rect 1636 47948 1642 47960
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 31294 47744 31300 47796
rect 31352 47784 31358 47796
rect 40402 47784 40408 47796
rect 31352 47756 40408 47784
rect 31352 47744 31358 47756
rect 40402 47744 40408 47756
rect 40460 47744 40466 47796
rect 30650 47676 30656 47728
rect 30708 47716 30714 47728
rect 44082 47716 44088 47728
rect 30708 47688 44088 47716
rect 30708 47676 30714 47688
rect 44082 47676 44088 47688
rect 44140 47676 44146 47728
rect 934 47608 940 47660
rect 992 47648 998 47660
rect 1673 47651 1731 47657
rect 1673 47648 1685 47651
rect 992 47620 1685 47648
rect 992 47608 998 47620
rect 1673 47617 1685 47620
rect 1719 47617 1731 47651
rect 1673 47611 1731 47617
rect 9122 47608 9128 47660
rect 9180 47648 9186 47660
rect 34514 47648 34520 47660
rect 9180 47620 34520 47648
rect 9180 47608 9186 47620
rect 34514 47608 34520 47620
rect 34572 47608 34578 47660
rect 58066 47608 58072 47660
rect 58124 47608 58130 47660
rect 3418 47540 3424 47592
rect 3476 47580 3482 47592
rect 32214 47580 32220 47592
rect 3476 47552 32220 47580
rect 3476 47540 3482 47552
rect 32214 47540 32220 47552
rect 32272 47540 32278 47592
rect 1762 47404 1768 47456
rect 1820 47404 1826 47456
rect 58253 47447 58311 47453
rect 58253 47413 58265 47447
rect 58299 47444 58311 47447
rect 58802 47444 58808 47456
rect 58299 47416 58808 47444
rect 58299 47413 58311 47416
rect 58253 47407 58311 47413
rect 58802 47404 58808 47416
rect 58860 47404 58866 47456
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 1765 47175 1823 47181
rect 1765 47141 1777 47175
rect 1811 47172 1823 47175
rect 8938 47172 8944 47184
rect 1811 47144 8944 47172
rect 1811 47141 1823 47144
rect 1765 47135 1823 47141
rect 8938 47132 8944 47144
rect 8996 47132 9002 47184
rect 934 46996 940 47048
rect 992 47036 998 47048
rect 1581 47039 1639 47045
rect 1581 47036 1593 47039
rect 992 47008 1593 47036
rect 992 46996 998 47008
rect 1581 47005 1593 47008
rect 1627 47005 1639 47039
rect 1581 46999 1639 47005
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 934 46520 940 46572
rect 992 46560 998 46572
rect 1581 46563 1639 46569
rect 1581 46560 1593 46563
rect 992 46532 1593 46560
rect 992 46520 998 46532
rect 1581 46529 1593 46532
rect 1627 46529 1639 46563
rect 1581 46523 1639 46529
rect 1765 46359 1823 46365
rect 1765 46325 1777 46359
rect 1811 46356 1823 46359
rect 36354 46356 36360 46368
rect 1811 46328 36360 46356
rect 1811 46325 1823 46328
rect 1765 46319 1823 46325
rect 36354 46316 36360 46328
rect 36412 46316 36418 46368
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 58158 45976 58164 46028
rect 58216 45976 58222 46028
rect 57698 45908 57704 45960
rect 57756 45948 57762 45960
rect 57885 45951 57943 45957
rect 57885 45948 57897 45951
rect 57756 45920 57897 45948
rect 57756 45908 57762 45920
rect 57885 45917 57897 45920
rect 57931 45917 57943 45951
rect 57885 45911 57943 45917
rect 934 45840 940 45892
rect 992 45880 998 45892
rect 1673 45883 1731 45889
rect 1673 45880 1685 45883
rect 992 45852 1685 45880
rect 992 45840 998 45852
rect 1673 45849 1685 45852
rect 1719 45849 1731 45883
rect 1673 45843 1731 45849
rect 1765 45815 1823 45821
rect 1765 45781 1777 45815
rect 1811 45812 1823 45815
rect 15194 45812 15200 45824
rect 1811 45784 15200 45812
rect 1811 45781 1823 45784
rect 1765 45775 1823 45781
rect 15194 45772 15200 45784
rect 15252 45772 15258 45824
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 17420 45580 17632 45608
rect 15194 45500 15200 45552
rect 15252 45540 15258 45552
rect 17420 45540 17448 45580
rect 15252 45512 17264 45540
rect 15252 45500 15258 45512
rect 17236 45481 17264 45512
rect 17328 45512 17448 45540
rect 17129 45475 17187 45481
rect 17129 45441 17141 45475
rect 17175 45441 17187 45475
rect 17129 45435 17187 45441
rect 17222 45475 17280 45481
rect 17222 45441 17234 45475
rect 17268 45441 17280 45475
rect 17222 45435 17280 45441
rect 17144 45404 17172 45435
rect 17328 45404 17356 45512
rect 17494 45500 17500 45552
rect 17552 45500 17558 45552
rect 17604 45540 17632 45580
rect 17604 45512 26234 45540
rect 17405 45475 17463 45481
rect 17405 45441 17417 45475
rect 17451 45441 17463 45475
rect 17405 45435 17463 45441
rect 17635 45475 17693 45481
rect 17635 45441 17647 45475
rect 17681 45472 17693 45475
rect 21082 45472 21088 45484
rect 17681 45444 21088 45472
rect 17681 45441 17693 45444
rect 17635 45435 17693 45441
rect 17144 45376 17356 45404
rect 17420 45404 17448 45435
rect 21082 45432 21088 45444
rect 21140 45432 21146 45484
rect 21450 45404 21456 45416
rect 17420 45376 21456 45404
rect 9030 45296 9036 45348
rect 9088 45336 9094 45348
rect 17420 45336 17448 45376
rect 21450 45364 21456 45376
rect 21508 45364 21514 45416
rect 26206 45404 26234 45512
rect 33778 45500 33784 45552
rect 33836 45540 33842 45552
rect 36541 45543 36599 45549
rect 36541 45540 36553 45543
rect 33836 45512 36553 45540
rect 33836 45500 33842 45512
rect 36541 45509 36553 45512
rect 36587 45509 36599 45543
rect 38197 45543 38255 45549
rect 38197 45540 38209 45543
rect 36541 45503 36599 45509
rect 37384 45512 38209 45540
rect 37384 45484 37412 45512
rect 38197 45509 38209 45512
rect 38243 45509 38255 45543
rect 38197 45503 38255 45509
rect 38289 45543 38347 45549
rect 38289 45509 38301 45543
rect 38335 45540 38347 45543
rect 57054 45540 57060 45552
rect 38335 45512 57060 45540
rect 38335 45509 38347 45512
rect 38289 45503 38347 45509
rect 57054 45500 57060 45512
rect 57112 45500 57118 45552
rect 36354 45432 36360 45484
rect 36412 45432 36418 45484
rect 36630 45432 36636 45484
rect 36688 45432 36694 45484
rect 36725 45475 36783 45481
rect 36725 45441 36737 45475
rect 36771 45472 36783 45475
rect 37366 45472 37372 45484
rect 36771 45444 37372 45472
rect 36771 45441 36783 45444
rect 36725 45435 36783 45441
rect 37366 45432 37372 45444
rect 37424 45432 37430 45484
rect 38010 45432 38016 45484
rect 38068 45432 38074 45484
rect 38470 45481 38476 45484
rect 38433 45475 38476 45481
rect 38433 45441 38445 45475
rect 38433 45435 38476 45441
rect 38470 45432 38476 45435
rect 38528 45432 38534 45484
rect 58069 45475 58127 45481
rect 58069 45441 58081 45475
rect 58115 45472 58127 45475
rect 58986 45472 58992 45484
rect 58115 45444 58992 45472
rect 58115 45441 58127 45444
rect 58069 45435 58127 45441
rect 58986 45432 58992 45444
rect 59044 45432 59050 45484
rect 26206 45376 38608 45404
rect 9088 45308 17448 45336
rect 9088 45296 9094 45308
rect 36906 45296 36912 45348
rect 36964 45296 36970 45348
rect 38580 45345 38608 45376
rect 38565 45339 38623 45345
rect 38565 45305 38577 45339
rect 38611 45305 38623 45339
rect 38565 45299 38623 45305
rect 17770 45228 17776 45280
rect 17828 45228 17834 45280
rect 58253 45271 58311 45277
rect 58253 45237 58265 45271
rect 58299 45268 58311 45271
rect 58434 45268 58440 45280
rect 58299 45240 58440 45268
rect 58299 45237 58311 45240
rect 58253 45231 58311 45237
rect 58434 45228 58440 45240
rect 58492 45228 58498 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 35434 45024 35440 45076
rect 35492 45024 35498 45076
rect 35250 44996 35256 45008
rect 26206 44968 35256 44996
rect 21266 44888 21272 44940
rect 21324 44928 21330 44940
rect 26206 44928 26234 44968
rect 35250 44956 35256 44968
rect 35308 44956 35314 45008
rect 21324 44900 26234 44928
rect 34900 44900 35388 44928
rect 21324 44888 21330 44900
rect 934 44820 940 44872
rect 992 44860 998 44872
rect 1581 44863 1639 44869
rect 1581 44860 1593 44863
rect 992 44832 1593 44860
rect 992 44820 998 44832
rect 1581 44829 1593 44832
rect 1627 44829 1639 44863
rect 1581 44823 1639 44829
rect 1854 44820 1860 44872
rect 1912 44820 1918 44872
rect 34900 44869 34928 44900
rect 34885 44863 34943 44869
rect 34885 44829 34897 44863
rect 34931 44829 34943 44863
rect 34885 44823 34943 44829
rect 35066 44820 35072 44872
rect 35124 44820 35130 44872
rect 35250 44820 35256 44872
rect 35308 44869 35314 44872
rect 35308 44823 35316 44869
rect 35360 44860 35388 44900
rect 45738 44860 45744 44872
rect 35360 44832 45744 44860
rect 35308 44820 35314 44823
rect 45738 44820 45744 44832
rect 45796 44820 45802 44872
rect 56962 44820 56968 44872
rect 57020 44820 57026 44872
rect 57241 44863 57299 44869
rect 57241 44829 57253 44863
rect 57287 44860 57299 44863
rect 58986 44860 58992 44872
rect 57287 44832 58992 44860
rect 57287 44829 57299 44832
rect 57241 44823 57299 44829
rect 58986 44820 58992 44832
rect 59044 44820 59050 44872
rect 9214 44752 9220 44804
rect 9272 44792 9278 44804
rect 35161 44795 35219 44801
rect 35161 44792 35173 44795
rect 9272 44764 35173 44792
rect 9272 44752 9278 44764
rect 35161 44761 35173 44764
rect 35207 44761 35219 44795
rect 35161 44755 35219 44761
rect 57977 44795 58035 44801
rect 57977 44761 57989 44795
rect 58023 44792 58035 44795
rect 58710 44792 58716 44804
rect 58023 44764 58716 44792
rect 58023 44761 58035 44764
rect 57977 44755 58035 44761
rect 58710 44752 58716 44764
rect 58768 44752 58774 44804
rect 58253 44727 58311 44733
rect 58253 44693 58265 44727
rect 58299 44724 58311 44727
rect 58342 44724 58348 44736
rect 58299 44696 58348 44724
rect 58299 44693 58311 44696
rect 58253 44687 58311 44693
rect 58342 44684 58348 44696
rect 58400 44684 58406 44736
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 934 44344 940 44396
rect 992 44384 998 44396
rect 1673 44387 1731 44393
rect 1673 44384 1685 44387
rect 992 44356 1685 44384
rect 992 44344 998 44356
rect 1673 44353 1685 44356
rect 1719 44353 1731 44387
rect 1673 44347 1731 44353
rect 1857 44251 1915 44257
rect 1857 44217 1869 44251
rect 1903 44248 1915 44251
rect 9582 44248 9588 44260
rect 1903 44220 9588 44248
rect 1903 44217 1915 44220
rect 1857 44211 1915 44217
rect 9582 44208 9588 44220
rect 9640 44208 9646 44260
rect 34698 44140 34704 44192
rect 34756 44180 34762 44192
rect 35066 44180 35072 44192
rect 34756 44152 35072 44180
rect 34756 44140 34762 44152
rect 35066 44140 35072 44152
rect 35124 44140 35130 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 34238 43868 34244 43920
rect 34296 43868 34302 43920
rect 9582 43732 9588 43784
rect 9640 43772 9646 43784
rect 33689 43775 33747 43781
rect 33689 43772 33701 43775
rect 9640 43744 33701 43772
rect 9640 43732 9646 43744
rect 33689 43741 33701 43744
rect 33735 43741 33747 43775
rect 33689 43735 33747 43741
rect 34054 43732 34060 43784
rect 34112 43781 34118 43784
rect 34112 43772 34120 43781
rect 34112 43744 34157 43772
rect 34112 43735 34120 43744
rect 34112 43732 34118 43735
rect 53834 43732 53840 43784
rect 53892 43772 53898 43784
rect 57885 43775 57943 43781
rect 57885 43772 57897 43775
rect 53892 43744 57897 43772
rect 53892 43732 53898 43744
rect 57885 43741 57897 43744
rect 57931 43741 57943 43775
rect 57885 43735 57943 43741
rect 934 43664 940 43716
rect 992 43704 998 43716
rect 1673 43707 1731 43713
rect 1673 43704 1685 43707
rect 992 43676 1685 43704
rect 992 43664 998 43676
rect 1673 43673 1685 43676
rect 1719 43673 1731 43707
rect 1673 43667 1731 43673
rect 33778 43664 33784 43716
rect 33836 43704 33842 43716
rect 33873 43707 33931 43713
rect 33873 43704 33885 43707
rect 33836 43676 33885 43704
rect 33836 43664 33842 43676
rect 33873 43673 33885 43676
rect 33919 43673 33931 43707
rect 33873 43667 33931 43673
rect 33965 43707 34023 43713
rect 33965 43673 33977 43707
rect 34011 43704 34023 43707
rect 35894 43704 35900 43716
rect 34011 43676 35900 43704
rect 34011 43673 34023 43676
rect 33965 43667 34023 43673
rect 35894 43664 35900 43676
rect 35952 43664 35958 43716
rect 58158 43664 58164 43716
rect 58216 43664 58222 43716
rect 1765 43639 1823 43645
rect 1765 43605 1777 43639
rect 1811 43636 1823 43639
rect 32306 43636 32312 43648
rect 1811 43608 32312 43636
rect 1811 43605 1823 43608
rect 1765 43599 1823 43605
rect 32306 43596 32312 43608
rect 32364 43596 32370 43648
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 32585 43367 32643 43373
rect 32585 43333 32597 43367
rect 32631 43364 32643 43367
rect 32631 43336 35894 43364
rect 32631 43333 32643 43336
rect 32585 43327 32643 43333
rect 934 43256 940 43308
rect 992 43296 998 43308
rect 1581 43299 1639 43305
rect 1581 43296 1593 43299
rect 992 43268 1593 43296
rect 992 43256 998 43268
rect 1581 43265 1593 43268
rect 1627 43265 1639 43299
rect 1581 43259 1639 43265
rect 32306 43256 32312 43308
rect 32364 43256 32370 43308
rect 32490 43256 32496 43308
rect 32548 43256 32554 43308
rect 32674 43256 32680 43308
rect 32732 43305 32738 43308
rect 32732 43296 32740 43305
rect 35866 43296 35894 43336
rect 54846 43296 54852 43308
rect 32732 43268 32777 43296
rect 35866 43268 54852 43296
rect 32732 43259 32740 43268
rect 32732 43256 32738 43259
rect 54846 43256 54852 43268
rect 54904 43256 54910 43308
rect 1762 43052 1768 43104
rect 1820 43052 1826 43104
rect 31754 43052 31760 43104
rect 31812 43092 31818 43104
rect 32861 43095 32919 43101
rect 32861 43092 32873 43095
rect 31812 43064 32873 43092
rect 31812 43052 31818 43064
rect 32861 43061 32873 43064
rect 32907 43061 32919 43095
rect 32861 43055 32919 43061
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 32674 42780 32680 42832
rect 32732 42820 32738 42832
rect 32732 42792 33916 42820
rect 32732 42780 32738 42792
rect 24302 42712 24308 42764
rect 24360 42752 24366 42764
rect 32490 42752 32496 42764
rect 24360 42724 32496 42752
rect 24360 42712 24366 42724
rect 32490 42712 32496 42724
rect 32548 42752 32554 42764
rect 33778 42752 33784 42764
rect 32548 42724 33784 42752
rect 32548 42712 32554 42724
rect 33042 42684 33048 42696
rect 26206 42656 33048 42684
rect 22186 42576 22192 42628
rect 22244 42616 22250 42628
rect 24394 42616 24400 42628
rect 22244 42588 24400 42616
rect 22244 42576 22250 42588
rect 24394 42576 24400 42588
rect 24452 42616 24458 42628
rect 26206 42616 26234 42656
rect 33042 42644 33048 42656
rect 33100 42644 33106 42696
rect 33134 42644 33140 42696
rect 33192 42644 33198 42696
rect 33704 42693 33732 42724
rect 33778 42712 33784 42724
rect 33836 42712 33842 42764
rect 33888 42752 33916 42792
rect 33888 42724 37688 42752
rect 33413 42687 33471 42693
rect 33413 42653 33425 42687
rect 33459 42653 33471 42687
rect 33413 42647 33471 42653
rect 33689 42687 33747 42693
rect 33689 42653 33701 42687
rect 33735 42653 33747 42687
rect 33689 42647 33747 42653
rect 24452 42588 26234 42616
rect 24452 42576 24458 42588
rect 32030 42576 32036 42628
rect 32088 42616 32094 42628
rect 32585 42619 32643 42625
rect 32585 42616 32597 42619
rect 32088 42588 32597 42616
rect 32088 42576 32094 42588
rect 32585 42585 32597 42588
rect 32631 42585 32643 42619
rect 32585 42579 32643 42585
rect 33428 42548 33456 42647
rect 33870 42644 33876 42696
rect 33928 42644 33934 42696
rect 37274 42644 37280 42696
rect 37332 42644 37338 42696
rect 37660 42693 37688 42724
rect 37645 42687 37703 42693
rect 37645 42653 37657 42687
rect 37691 42653 37703 42687
rect 37645 42647 37703 42653
rect 57057 42687 57115 42693
rect 57057 42653 57069 42687
rect 57103 42684 57115 42687
rect 58986 42684 58992 42696
rect 57103 42656 58992 42684
rect 57103 42653 57115 42656
rect 57057 42647 57115 42653
rect 58986 42644 58992 42656
rect 59044 42644 59050 42696
rect 37366 42576 37372 42628
rect 37424 42616 37430 42628
rect 37461 42619 37519 42625
rect 37461 42616 37473 42619
rect 37424 42588 37473 42616
rect 37424 42576 37430 42588
rect 37461 42585 37473 42588
rect 37507 42585 37519 42619
rect 37461 42579 37519 42585
rect 37553 42619 37611 42625
rect 37553 42585 37565 42619
rect 37599 42616 37611 42619
rect 54294 42616 54300 42628
rect 37599 42588 54300 42616
rect 37599 42585 37611 42588
rect 37553 42579 37611 42585
rect 54294 42576 54300 42588
rect 54352 42576 54358 42628
rect 57974 42576 57980 42628
rect 58032 42576 58038 42628
rect 58345 42619 58403 42625
rect 58345 42585 58357 42619
rect 58391 42616 58403 42619
rect 58526 42616 58532 42628
rect 58391 42588 58532 42616
rect 58391 42585 58403 42588
rect 58345 42579 58403 42585
rect 58526 42576 58532 42588
rect 58584 42576 58590 42628
rect 37829 42551 37887 42557
rect 37829 42548 37841 42551
rect 33428 42520 37841 42548
rect 37829 42517 37841 42520
rect 37875 42517 37887 42551
rect 37829 42511 37887 42517
rect 39298 42508 39304 42560
rect 39356 42548 39362 42560
rect 57149 42551 57207 42557
rect 57149 42548 57161 42551
rect 39356 42520 57161 42548
rect 39356 42508 39362 42520
rect 57149 42517 57161 42520
rect 57195 42517 57207 42551
rect 57149 42511 57207 42517
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 37274 42304 37280 42356
rect 37332 42344 37338 42356
rect 39390 42344 39396 42356
rect 37332 42316 39396 42344
rect 37332 42304 37338 42316
rect 39390 42304 39396 42316
rect 39448 42304 39454 42356
rect 934 42168 940 42220
rect 992 42208 998 42220
rect 1581 42211 1639 42217
rect 1581 42208 1593 42211
rect 992 42180 1593 42208
rect 992 42168 998 42180
rect 1581 42177 1593 42180
rect 1627 42177 1639 42211
rect 1581 42171 1639 42177
rect 1762 42168 1768 42220
rect 1820 42208 1826 42220
rect 33870 42208 33876 42220
rect 1820 42180 33876 42208
rect 1820 42168 1826 42180
rect 33870 42168 33876 42180
rect 33928 42168 33934 42220
rect 13078 42100 13084 42152
rect 13136 42140 13142 42152
rect 23658 42140 23664 42152
rect 13136 42112 23664 42140
rect 13136 42100 13142 42112
rect 23658 42100 23664 42112
rect 23716 42100 23722 42152
rect 33134 42100 33140 42152
rect 33192 42140 33198 42152
rect 33778 42140 33784 42152
rect 33192 42112 33784 42140
rect 33192 42100 33198 42112
rect 33778 42100 33784 42112
rect 33836 42140 33842 42152
rect 34054 42140 34060 42152
rect 33836 42112 34060 42140
rect 33836 42100 33842 42112
rect 34054 42100 34060 42112
rect 34112 42100 34118 42152
rect 6454 42032 6460 42084
rect 6512 42072 6518 42084
rect 22554 42072 22560 42084
rect 6512 42044 22560 42072
rect 6512 42032 6518 42044
rect 22554 42032 22560 42044
rect 22612 42032 22618 42084
rect 1765 42007 1823 42013
rect 1765 41973 1777 42007
rect 1811 42004 1823 42007
rect 2130 42004 2136 42016
rect 1811 41976 2136 42004
rect 1811 41973 1823 41976
rect 1765 41967 1823 41973
rect 2130 41964 2136 41976
rect 2188 41964 2194 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 53558 41556 53564 41608
rect 53616 41596 53622 41608
rect 56965 41599 57023 41605
rect 56965 41596 56977 41599
rect 53616 41568 56977 41596
rect 53616 41556 53622 41568
rect 56965 41565 56977 41568
rect 57011 41565 57023 41599
rect 56965 41559 57023 41565
rect 57241 41599 57299 41605
rect 57241 41565 57253 41599
rect 57287 41596 57299 41599
rect 58986 41596 58992 41608
rect 57287 41568 58992 41596
rect 57287 41565 57299 41568
rect 57241 41559 57299 41565
rect 58986 41556 58992 41568
rect 59044 41556 59050 41608
rect 934 41488 940 41540
rect 992 41528 998 41540
rect 1673 41531 1731 41537
rect 1673 41528 1685 41531
rect 992 41500 1685 41528
rect 992 41488 998 41500
rect 1673 41497 1685 41500
rect 1719 41497 1731 41531
rect 1673 41491 1731 41497
rect 2041 41531 2099 41537
rect 2041 41497 2053 41531
rect 2087 41528 2099 41531
rect 6362 41528 6368 41540
rect 2087 41500 6368 41528
rect 2087 41497 2099 41500
rect 2041 41491 2099 41497
rect 6362 41488 6368 41500
rect 6420 41488 6426 41540
rect 57977 41531 58035 41537
rect 57977 41497 57989 41531
rect 58023 41528 58035 41531
rect 58710 41528 58716 41540
rect 58023 41500 58716 41528
rect 58023 41497 58035 41500
rect 57977 41491 58035 41497
rect 58710 41488 58716 41500
rect 58768 41488 58774 41540
rect 50062 41420 50068 41472
rect 50120 41460 50126 41472
rect 53834 41460 53840 41472
rect 50120 41432 53840 41460
rect 50120 41420 50126 41432
rect 53834 41420 53840 41432
rect 53892 41420 53898 41472
rect 58253 41463 58311 41469
rect 58253 41429 58265 41463
rect 58299 41460 58311 41463
rect 58618 41460 58624 41472
rect 58299 41432 58624 41460
rect 58299 41429 58311 41432
rect 58253 41423 58311 41429
rect 58618 41420 58624 41432
rect 58676 41420 58682 41472
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 934 41080 940 41132
rect 992 41120 998 41132
rect 1673 41123 1731 41129
rect 1673 41120 1685 41123
rect 992 41092 1685 41120
rect 992 41080 998 41092
rect 1673 41089 1685 41092
rect 1719 41089 1731 41123
rect 1673 41083 1731 41089
rect 1765 40919 1823 40925
rect 1765 40885 1777 40919
rect 1811 40916 1823 40919
rect 21174 40916 21180 40928
rect 1811 40888 21180 40916
rect 1811 40885 1823 40888
rect 1765 40879 1823 40885
rect 21174 40876 21180 40888
rect 21232 40876 21238 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 28442 40672 28448 40724
rect 28500 40712 28506 40724
rect 41414 40712 41420 40724
rect 28500 40684 41420 40712
rect 28500 40672 28506 40684
rect 41414 40672 41420 40684
rect 41472 40672 41478 40724
rect 54662 40468 54668 40520
rect 54720 40508 54726 40520
rect 57885 40511 57943 40517
rect 57885 40508 57897 40511
rect 54720 40480 57897 40508
rect 54720 40468 54726 40480
rect 57885 40477 57897 40480
rect 57931 40477 57943 40511
rect 57885 40471 57943 40477
rect 934 40400 940 40452
rect 992 40440 998 40452
rect 1673 40443 1731 40449
rect 1673 40440 1685 40443
rect 992 40412 1685 40440
rect 992 40400 998 40412
rect 1673 40409 1685 40412
rect 1719 40409 1731 40443
rect 1673 40403 1731 40409
rect 57057 40443 57115 40449
rect 57057 40409 57069 40443
rect 57103 40440 57115 40443
rect 58161 40443 58219 40449
rect 57103 40412 58112 40440
rect 57103 40409 57115 40412
rect 57057 40403 57115 40409
rect 1765 40375 1823 40381
rect 1765 40341 1777 40375
rect 1811 40372 1823 40375
rect 11698 40372 11704 40384
rect 1811 40344 11704 40372
rect 1811 40341 1823 40344
rect 1765 40335 1823 40341
rect 11698 40332 11704 40344
rect 11756 40332 11762 40384
rect 56042 40332 56048 40384
rect 56100 40372 56106 40384
rect 57149 40375 57207 40381
rect 57149 40372 57161 40375
rect 56100 40344 57161 40372
rect 56100 40332 56106 40344
rect 57149 40341 57161 40344
rect 57195 40341 57207 40375
rect 58084 40372 58112 40412
rect 58161 40409 58173 40443
rect 58207 40440 58219 40443
rect 58986 40440 58992 40452
rect 58207 40412 58992 40440
rect 58207 40409 58219 40412
rect 58161 40403 58219 40409
rect 58986 40400 58992 40412
rect 59044 40400 59050 40452
rect 58710 40372 58716 40384
rect 58084 40344 58716 40372
rect 57149 40335 57207 40341
rect 58710 40332 58716 40344
rect 58768 40332 58774 40384
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 20898 40128 20904 40180
rect 20956 40128 20962 40180
rect 58342 40128 58348 40180
rect 58400 40168 58406 40180
rect 58710 40168 58716 40180
rect 58400 40140 58716 40168
rect 58400 40128 58406 40140
rect 58710 40128 58716 40140
rect 58768 40128 58774 40180
rect 1026 40060 1032 40112
rect 1084 40100 1090 40112
rect 1673 40103 1731 40109
rect 1673 40100 1685 40103
rect 1084 40072 1685 40100
rect 1084 40060 1090 40072
rect 1673 40069 1685 40072
rect 1719 40069 1731 40103
rect 1673 40063 1731 40069
rect 20916 40041 20944 40128
rect 21082 40060 21088 40112
rect 21140 40060 21146 40112
rect 21174 40060 21180 40112
rect 21232 40060 21238 40112
rect 20901 40035 20959 40041
rect 20901 40001 20913 40035
rect 20947 40001 20959 40035
rect 20901 39995 20959 40001
rect 21269 40035 21327 40041
rect 21269 40001 21281 40035
rect 21315 40032 21327 40035
rect 21634 40032 21640 40044
rect 21315 40004 21640 40032
rect 21315 40001 21327 40004
rect 21269 39995 21327 40001
rect 21634 39992 21640 40004
rect 21692 39992 21698 40044
rect 1765 39831 1823 39837
rect 1765 39797 1777 39831
rect 1811 39828 1823 39831
rect 2590 39828 2596 39840
rect 1811 39800 2596 39828
rect 1811 39797 1823 39800
rect 1765 39791 1823 39797
rect 2590 39788 2596 39800
rect 2648 39788 2654 39840
rect 21453 39831 21511 39837
rect 21453 39797 21465 39831
rect 21499 39828 21511 39831
rect 22278 39828 22284 39840
rect 21499 39800 22284 39828
rect 21499 39797 21511 39800
rect 21453 39791 21511 39797
rect 22278 39788 22284 39800
rect 22336 39788 22342 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 2682 39516 2688 39568
rect 2740 39516 2746 39568
rect 2869 39559 2927 39565
rect 2869 39525 2881 39559
rect 2915 39556 2927 39559
rect 22646 39556 22652 39568
rect 2915 39528 22652 39556
rect 2915 39525 2927 39528
rect 2869 39519 2927 39525
rect 22646 39516 22652 39528
rect 22704 39516 22710 39568
rect 2222 39448 2228 39500
rect 2280 39488 2286 39500
rect 2700 39488 2728 39516
rect 2280 39460 2728 39488
rect 2280 39448 2286 39460
rect 2314 39380 2320 39432
rect 2372 39380 2378 39432
rect 2516 39429 2544 39460
rect 2501 39423 2559 39429
rect 2501 39389 2513 39423
rect 2547 39389 2559 39423
rect 2501 39383 2559 39389
rect 2590 39380 2596 39432
rect 2648 39380 2654 39432
rect 2682 39380 2688 39432
rect 2740 39429 2746 39432
rect 2740 39420 2748 39429
rect 57057 39423 57115 39429
rect 2740 39392 2785 39420
rect 2740 39383 2748 39392
rect 57057 39389 57069 39423
rect 57103 39420 57115 39423
rect 58986 39420 58992 39432
rect 57103 39392 58992 39420
rect 57103 39389 57115 39392
rect 57057 39383 57115 39389
rect 2740 39380 2746 39383
rect 58986 39380 58992 39392
rect 59044 39380 59050 39432
rect 934 39312 940 39364
rect 992 39352 998 39364
rect 1673 39355 1731 39361
rect 1673 39352 1685 39355
rect 992 39324 1685 39352
rect 992 39312 998 39324
rect 1673 39321 1685 39324
rect 1719 39321 1731 39355
rect 1673 39315 1731 39321
rect 29638 39312 29644 39364
rect 29696 39352 29702 39364
rect 53466 39352 53472 39364
rect 29696 39324 53472 39352
rect 29696 39312 29702 39324
rect 53466 39312 53472 39324
rect 53524 39312 53530 39364
rect 57974 39312 57980 39364
rect 58032 39312 58038 39364
rect 58342 39312 58348 39364
rect 58400 39312 58406 39364
rect 1765 39287 1823 39293
rect 1765 39253 1777 39287
rect 1811 39284 1823 39287
rect 3050 39284 3056 39296
rect 1811 39256 3056 39284
rect 1811 39253 1823 39256
rect 1765 39247 1823 39253
rect 3050 39244 3056 39256
rect 3108 39244 3114 39296
rect 33502 39244 33508 39296
rect 33560 39284 33566 39296
rect 57149 39287 57207 39293
rect 57149 39284 57161 39287
rect 33560 39256 57161 39284
rect 33560 39244 33566 39256
rect 57149 39253 57161 39256
rect 57195 39253 57207 39287
rect 57149 39247 57207 39253
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 1026 38904 1032 38956
rect 1084 38944 1090 38956
rect 1673 38947 1731 38953
rect 1673 38944 1685 38947
rect 1084 38916 1685 38944
rect 1084 38904 1090 38916
rect 1673 38913 1685 38916
rect 1719 38913 1731 38947
rect 1673 38907 1731 38913
rect 20530 38904 20536 38956
rect 20588 38944 20594 38956
rect 22005 38947 22063 38953
rect 22005 38944 22017 38947
rect 20588 38916 22017 38944
rect 20588 38904 20594 38916
rect 22005 38913 22017 38916
rect 22051 38913 22063 38947
rect 22005 38907 22063 38913
rect 22278 38904 22284 38956
rect 22336 38904 22342 38956
rect 22462 38836 22468 38888
rect 22520 38836 22526 38888
rect 19978 38768 19984 38820
rect 20036 38808 20042 38820
rect 20254 38808 20260 38820
rect 20036 38780 20260 38808
rect 20036 38768 20042 38780
rect 20254 38768 20260 38780
rect 20312 38768 20318 38820
rect 22097 38811 22155 38817
rect 22097 38777 22109 38811
rect 22143 38808 22155 38811
rect 23106 38808 23112 38820
rect 22143 38780 23112 38808
rect 22143 38777 22155 38780
rect 22097 38771 22155 38777
rect 23106 38768 23112 38780
rect 23164 38768 23170 38820
rect 1765 38743 1823 38749
rect 1765 38709 1777 38743
rect 1811 38740 1823 38743
rect 19426 38740 19432 38752
rect 1811 38712 19432 38740
rect 1811 38709 1823 38712
rect 1765 38703 1823 38709
rect 19426 38700 19432 38712
rect 19484 38700 19490 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 16206 38496 16212 38548
rect 16264 38536 16270 38548
rect 20073 38539 20131 38545
rect 20073 38536 20085 38539
rect 16264 38508 20085 38536
rect 16264 38496 16270 38508
rect 20073 38505 20085 38508
rect 20119 38505 20131 38539
rect 20073 38499 20131 38505
rect 20898 38496 20904 38548
rect 20956 38536 20962 38548
rect 21082 38536 21088 38548
rect 20956 38508 21088 38536
rect 20956 38496 20962 38508
rect 21082 38496 21088 38508
rect 21140 38536 21146 38548
rect 25314 38536 25320 38548
rect 21140 38508 25320 38536
rect 21140 38496 21146 38508
rect 25314 38496 25320 38508
rect 25372 38496 25378 38548
rect 1854 38428 1860 38480
rect 1912 38468 1918 38480
rect 20990 38468 20996 38480
rect 1912 38440 20996 38468
rect 1912 38428 1918 38440
rect 20990 38428 20996 38440
rect 21048 38428 21054 38480
rect 23106 38428 23112 38480
rect 23164 38468 23170 38480
rect 23382 38468 23388 38480
rect 23164 38440 23388 38468
rect 23164 38428 23170 38440
rect 1670 38360 1676 38412
rect 1728 38400 1734 38412
rect 1728 38372 2636 38400
rect 1728 38360 1734 38372
rect 1946 38292 1952 38344
rect 2004 38332 2010 38344
rect 2041 38335 2099 38341
rect 2041 38332 2053 38335
rect 2004 38304 2053 38332
rect 2004 38292 2010 38304
rect 2041 38301 2053 38304
rect 2087 38301 2099 38335
rect 2041 38295 2099 38301
rect 2406 38292 2412 38344
rect 2464 38292 2470 38344
rect 2608 38332 2636 38372
rect 3050 38360 3056 38412
rect 3108 38360 3114 38412
rect 11698 38360 11704 38412
rect 11756 38400 11762 38412
rect 11756 38372 20484 38400
rect 11756 38360 11762 38372
rect 2682 38332 2688 38344
rect 2608 38304 2688 38332
rect 2682 38292 2688 38304
rect 2740 38332 2746 38344
rect 3237 38335 3295 38341
rect 3237 38332 3249 38335
rect 2740 38304 3249 38332
rect 2740 38292 2746 38304
rect 3237 38301 3249 38304
rect 3283 38301 3295 38335
rect 3237 38295 3295 38301
rect 3421 38335 3479 38341
rect 3421 38301 3433 38335
rect 3467 38332 3479 38335
rect 20257 38335 20315 38341
rect 20257 38332 20269 38335
rect 3467 38304 20269 38332
rect 3467 38301 3479 38304
rect 3421 38295 3479 38301
rect 20257 38301 20269 38304
rect 20303 38301 20315 38335
rect 20257 38295 20315 38301
rect 20346 38292 20352 38344
rect 20404 38292 20410 38344
rect 2225 38267 2283 38273
rect 2225 38233 2237 38267
rect 2271 38233 2283 38267
rect 2225 38227 2283 38233
rect 2240 38196 2268 38227
rect 2314 38224 2320 38276
rect 2372 38224 2378 38276
rect 19242 38264 19248 38276
rect 2516 38236 19248 38264
rect 2516 38196 2544 38236
rect 19242 38224 19248 38236
rect 19300 38224 19306 38276
rect 20073 38267 20131 38273
rect 20073 38233 20085 38267
rect 20119 38264 20131 38267
rect 20162 38264 20168 38276
rect 20119 38236 20168 38264
rect 20119 38233 20131 38236
rect 20073 38227 20131 38233
rect 20162 38224 20168 38236
rect 20220 38224 20226 38276
rect 20456 38264 20484 38372
rect 20714 38360 20720 38412
rect 20772 38400 20778 38412
rect 23216 38400 23244 38440
rect 23382 38428 23388 38440
rect 23440 38428 23446 38480
rect 26970 38400 26976 38412
rect 20772 38372 23244 38400
rect 23308 38372 26976 38400
rect 20772 38360 20778 38372
rect 22922 38292 22928 38344
rect 22980 38292 22986 38344
rect 23073 38335 23131 38341
rect 23073 38301 23085 38335
rect 23119 38332 23131 38335
rect 23308 38332 23336 38372
rect 26970 38360 26976 38372
rect 27028 38360 27034 38412
rect 23119 38304 23336 38332
rect 23119 38301 23131 38304
rect 23073 38295 23131 38301
rect 23382 38292 23388 38344
rect 23440 38341 23446 38344
rect 23440 38332 23448 38341
rect 23440 38304 23485 38332
rect 23440 38295 23448 38304
rect 23440 38292 23446 38295
rect 46842 38292 46848 38344
rect 46900 38332 46906 38344
rect 57885 38335 57943 38341
rect 57885 38332 57897 38335
rect 46900 38304 57897 38332
rect 46900 38292 46906 38304
rect 57885 38301 57897 38304
rect 57931 38301 57943 38335
rect 57885 38295 57943 38301
rect 20456 38236 22094 38264
rect 2240 38168 2544 38196
rect 2590 38156 2596 38208
rect 2648 38156 2654 38208
rect 19797 38199 19855 38205
rect 19797 38165 19809 38199
rect 19843 38196 19855 38199
rect 20346 38196 20352 38208
rect 19843 38168 20352 38196
rect 19843 38165 19855 38168
rect 19797 38159 19855 38165
rect 20346 38156 20352 38168
rect 20404 38156 20410 38208
rect 20533 38199 20591 38205
rect 20533 38165 20545 38199
rect 20579 38196 20591 38199
rect 21726 38196 21732 38208
rect 20579 38168 21732 38196
rect 20579 38165 20591 38168
rect 20533 38159 20591 38165
rect 21726 38156 21732 38168
rect 21784 38156 21790 38208
rect 22066 38196 22094 38236
rect 23198 38224 23204 38276
rect 23256 38224 23262 38276
rect 23293 38267 23351 38273
rect 23293 38233 23305 38267
rect 23339 38233 23351 38267
rect 23293 38227 23351 38233
rect 23308 38196 23336 38227
rect 58158 38224 58164 38276
rect 58216 38224 58222 38276
rect 22066 38168 23336 38196
rect 23566 38156 23572 38208
rect 23624 38156 23630 38208
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 2590 37952 2596 38004
rect 2648 37992 2654 38004
rect 16206 37992 16212 38004
rect 2648 37964 16212 37992
rect 2648 37952 2654 37964
rect 16206 37952 16212 37964
rect 16264 37952 16270 38004
rect 20349 37995 20407 38001
rect 19536 37964 19840 37992
rect 5902 37884 5908 37936
rect 5960 37924 5966 37936
rect 19536 37924 19564 37964
rect 5960 37896 19564 37924
rect 5960 37884 5966 37896
rect 19702 37884 19708 37936
rect 19760 37884 19766 37936
rect 19812 37924 19840 37964
rect 20349 37961 20361 37995
rect 20395 37992 20407 37995
rect 20806 37992 20812 38004
rect 20395 37964 20812 37992
rect 20395 37961 20407 37964
rect 20349 37955 20407 37961
rect 20806 37952 20812 37964
rect 20864 37952 20870 38004
rect 20990 37952 20996 38004
rect 21048 37952 21054 38004
rect 23293 37995 23351 38001
rect 23293 37961 23305 37995
rect 23339 37992 23351 37995
rect 23339 37964 23796 37992
rect 23339 37961 23351 37964
rect 23293 37955 23351 37961
rect 19812 37896 22784 37924
rect 934 37816 940 37868
rect 992 37856 998 37868
rect 1673 37859 1731 37865
rect 1673 37856 1685 37859
rect 992 37828 1685 37856
rect 992 37816 998 37828
rect 1673 37825 1685 37828
rect 1719 37825 1731 37859
rect 1673 37819 1731 37825
rect 16666 37816 16672 37868
rect 16724 37856 16730 37868
rect 16945 37859 17003 37865
rect 16945 37856 16957 37859
rect 16724 37828 16957 37856
rect 16724 37816 16730 37828
rect 16945 37825 16957 37828
rect 16991 37825 17003 37859
rect 16945 37819 17003 37825
rect 19334 37816 19340 37868
rect 19392 37816 19398 37868
rect 19457 37859 19515 37865
rect 19457 37825 19469 37859
rect 19503 37856 19515 37859
rect 19613 37859 19671 37865
rect 19503 37825 19528 37856
rect 19457 37819 19528 37825
rect 19613 37825 19625 37859
rect 19659 37856 19671 37859
rect 19843 37859 19901 37865
rect 19659 37828 19748 37856
rect 19659 37825 19671 37828
rect 19613 37819 19671 37825
rect 17497 37791 17555 37797
rect 17497 37757 17509 37791
rect 17543 37757 17555 37791
rect 17497 37751 17555 37757
rect 1854 37680 1860 37732
rect 1912 37680 1918 37732
rect 17512 37652 17540 37751
rect 19500 37720 19528 37819
rect 19720 37788 19748 37828
rect 19843 37825 19855 37859
rect 19889 37856 19901 37859
rect 20714 37856 20720 37868
rect 19889 37828 20720 37856
rect 19889 37825 19901 37828
rect 19843 37819 19901 37825
rect 20714 37816 20720 37828
rect 20772 37816 20778 37868
rect 20806 37816 20812 37868
rect 20864 37816 20870 37868
rect 21082 37816 21088 37868
rect 21140 37856 21146 37868
rect 21358 37856 21364 37868
rect 21140 37828 21364 37856
rect 21140 37816 21146 37828
rect 21358 37816 21364 37828
rect 21416 37816 21422 37868
rect 22756 37865 22784 37896
rect 22830 37884 22836 37936
rect 22888 37924 22894 37936
rect 23768 37933 23796 37964
rect 22925 37927 22983 37933
rect 22925 37924 22937 37927
rect 22888 37896 22937 37924
rect 22888 37884 22894 37896
rect 22925 37893 22937 37896
rect 22971 37893 22983 37927
rect 22925 37887 22983 37893
rect 23753 37927 23811 37933
rect 23753 37893 23765 37927
rect 23799 37893 23811 37927
rect 23753 37887 23811 37893
rect 24762 37884 24768 37936
rect 24820 37924 24826 37936
rect 25225 37927 25283 37933
rect 25225 37924 25237 37927
rect 24820 37896 25237 37924
rect 24820 37884 24826 37896
rect 25225 37893 25237 37896
rect 25271 37893 25283 37927
rect 25225 37887 25283 37893
rect 22741 37859 22799 37865
rect 22741 37825 22753 37859
rect 22787 37825 22799 37859
rect 22741 37819 22799 37825
rect 23014 37816 23020 37868
rect 23072 37816 23078 37868
rect 23109 37859 23167 37865
rect 23109 37825 23121 37859
rect 23155 37825 23167 37859
rect 23109 37819 23167 37825
rect 20622 37788 20628 37800
rect 19720 37760 20628 37788
rect 20622 37748 20628 37760
rect 20680 37748 20686 37800
rect 20824 37788 20852 37816
rect 21450 37788 21456 37800
rect 20824 37760 21456 37788
rect 21450 37748 21456 37760
rect 21508 37748 21514 37800
rect 22465 37791 22523 37797
rect 22465 37757 22477 37791
rect 22511 37788 22523 37791
rect 23032 37788 23060 37816
rect 22511 37760 23060 37788
rect 22511 37757 22523 37760
rect 22465 37751 22523 37757
rect 19794 37720 19800 37732
rect 19500 37692 19800 37720
rect 19794 37680 19800 37692
rect 19852 37680 19858 37732
rect 19904 37692 20760 37720
rect 19904 37652 19932 37692
rect 17512 37624 19932 37652
rect 19978 37612 19984 37664
rect 20036 37612 20042 37664
rect 20622 37612 20628 37664
rect 20680 37612 20686 37664
rect 20732 37652 20760 37692
rect 20806 37680 20812 37732
rect 20864 37720 20870 37732
rect 23124 37720 23152 37819
rect 23842 37816 23848 37868
rect 23900 37856 23906 37868
rect 23983 37859 24041 37865
rect 23983 37856 23995 37859
rect 23900 37828 23995 37856
rect 23900 37816 23906 37828
rect 23983 37825 23995 37828
rect 24029 37825 24041 37859
rect 23983 37819 24041 37825
rect 24949 37859 25007 37865
rect 24949 37825 24961 37859
rect 24995 37825 25007 37859
rect 24949 37819 25007 37825
rect 24118 37748 24124 37800
rect 24176 37788 24182 37800
rect 24394 37788 24400 37800
rect 24176 37760 24400 37788
rect 24176 37748 24182 37760
rect 24394 37748 24400 37760
rect 24452 37748 24458 37800
rect 24964 37788 24992 37819
rect 25130 37816 25136 37868
rect 25188 37816 25194 37868
rect 25314 37816 25320 37868
rect 25372 37816 25378 37868
rect 58066 37816 58072 37868
rect 58124 37816 58130 37868
rect 28258 37788 28264 37800
rect 24964 37760 28264 37788
rect 28258 37748 28264 37760
rect 28316 37748 28322 37800
rect 20864 37692 23152 37720
rect 23918 37723 23976 37729
rect 20864 37680 20870 37692
rect 23918 37689 23930 37723
rect 23964 37720 23976 37723
rect 25501 37723 25559 37729
rect 25501 37720 25513 37723
rect 23964 37692 25513 37720
rect 23964 37689 23976 37692
rect 23918 37683 23976 37689
rect 25501 37689 25513 37692
rect 25547 37689 25559 37723
rect 25501 37683 25559 37689
rect 22830 37652 22836 37664
rect 20732 37624 22836 37652
rect 22830 37612 22836 37624
rect 22888 37612 22894 37664
rect 24026 37612 24032 37664
rect 24084 37652 24090 37664
rect 24213 37655 24271 37661
rect 24213 37652 24225 37655
rect 24084 37624 24225 37652
rect 24084 37612 24090 37624
rect 24213 37621 24225 37624
rect 24259 37621 24271 37655
rect 24213 37615 24271 37621
rect 58253 37655 58311 37661
rect 58253 37621 58265 37655
rect 58299 37652 58311 37655
rect 59170 37652 59176 37664
rect 58299 37624 59176 37652
rect 58299 37621 58311 37624
rect 58253 37615 58311 37621
rect 59170 37612 59176 37624
rect 59228 37612 59234 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 19242 37408 19248 37460
rect 19300 37448 19306 37460
rect 21082 37448 21088 37460
rect 19300 37420 21088 37448
rect 19300 37408 19306 37420
rect 21082 37408 21088 37420
rect 21140 37408 21146 37460
rect 19794 37340 19800 37392
rect 19852 37380 19858 37392
rect 20346 37380 20352 37392
rect 19852 37352 20352 37380
rect 19852 37340 19858 37352
rect 20346 37340 20352 37352
rect 20404 37340 20410 37392
rect 20714 37340 20720 37392
rect 20772 37380 20778 37392
rect 22186 37380 22192 37392
rect 20772 37352 22192 37380
rect 20772 37340 20778 37352
rect 22186 37340 22192 37352
rect 22244 37340 22250 37392
rect 20898 37312 20904 37324
rect 5920 37284 6684 37312
rect 5920 37253 5948 37284
rect 5905 37247 5963 37253
rect 5905 37213 5917 37247
rect 5951 37213 5963 37247
rect 5905 37207 5963 37213
rect 5994 37204 6000 37256
rect 6052 37204 6058 37256
rect 6270 37204 6276 37256
rect 6328 37204 6334 37256
rect 6549 37247 6607 37253
rect 6549 37213 6561 37247
rect 6595 37213 6607 37247
rect 6549 37207 6607 37213
rect 2406 37136 2412 37188
rect 2464 37176 2470 37188
rect 2464 37148 5764 37176
rect 2464 37136 2470 37148
rect 5534 37068 5540 37120
rect 5592 37068 5598 37120
rect 5736 37108 5764 37148
rect 6564 37108 6592 37207
rect 6656 37176 6684 37284
rect 20180 37284 20904 37312
rect 6730 37204 6736 37256
rect 6788 37204 6794 37256
rect 19334 37204 19340 37256
rect 19392 37244 19398 37256
rect 19613 37247 19671 37253
rect 19613 37244 19625 37247
rect 19392 37216 19625 37244
rect 19392 37204 19398 37216
rect 19613 37213 19625 37216
rect 19659 37213 19671 37247
rect 19613 37207 19671 37213
rect 18874 37176 18880 37188
rect 6656 37148 18880 37176
rect 18874 37136 18880 37148
rect 18932 37136 18938 37188
rect 5736 37080 6592 37108
rect 19628 37108 19656 37207
rect 20180 37188 20208 37284
rect 20898 37272 20904 37284
rect 20956 37272 20962 37324
rect 21082 37272 21088 37324
rect 21140 37272 21146 37324
rect 31110 37272 31116 37324
rect 31168 37312 31174 37324
rect 33502 37312 33508 37324
rect 31168 37284 33508 37312
rect 31168 37272 31174 37284
rect 33502 37272 33508 37284
rect 33560 37272 33566 37324
rect 53668 37284 53880 37312
rect 20530 37204 20536 37256
rect 20588 37244 20594 37256
rect 20809 37247 20867 37253
rect 20809 37244 20821 37247
rect 20588 37216 20821 37244
rect 20588 37204 20594 37216
rect 20809 37213 20821 37216
rect 20855 37213 20867 37247
rect 28350 37244 28356 37256
rect 20809 37207 20867 37213
rect 20916 37216 28356 37244
rect 20162 37136 20168 37188
rect 20220 37136 20226 37188
rect 20916 37176 20944 37216
rect 28350 37204 28356 37216
rect 28408 37204 28414 37256
rect 53466 37204 53472 37256
rect 53524 37244 53530 37256
rect 53668 37244 53696 37284
rect 53524 37216 53696 37244
rect 53524 37204 53530 37216
rect 53742 37204 53748 37256
rect 53800 37204 53806 37256
rect 53852 37244 53880 37284
rect 54118 37247 54176 37253
rect 54118 37244 54130 37247
rect 53852 37216 54130 37244
rect 54118 37213 54130 37216
rect 54164 37213 54176 37247
rect 54118 37207 54176 37213
rect 54478 37204 54484 37256
rect 54536 37244 54542 37256
rect 57885 37247 57943 37253
rect 57885 37244 57897 37247
rect 54536 37216 57897 37244
rect 54536 37204 54542 37216
rect 57885 37213 57897 37216
rect 57931 37213 57943 37247
rect 57885 37207 57943 37213
rect 20364 37148 20944 37176
rect 26206 37148 45554 37176
rect 20364 37108 20392 37148
rect 19628 37080 20392 37108
rect 20438 37068 20444 37120
rect 20496 37108 20502 37120
rect 26206 37108 26234 37148
rect 20496 37080 26234 37108
rect 45526 37108 45554 37148
rect 53834 37136 53840 37188
rect 53892 37176 53898 37188
rect 53929 37179 53987 37185
rect 53929 37176 53941 37179
rect 53892 37148 53941 37176
rect 53892 37136 53898 37148
rect 53929 37145 53941 37148
rect 53975 37145 53987 37179
rect 53929 37139 53987 37145
rect 54021 37179 54079 37185
rect 54021 37145 54033 37179
rect 54067 37176 54079 37179
rect 56686 37176 56692 37188
rect 54067 37148 56692 37176
rect 54067 37145 54079 37148
rect 54021 37139 54079 37145
rect 56686 37136 56692 37148
rect 56744 37136 56750 37188
rect 58158 37136 58164 37188
rect 58216 37136 58222 37188
rect 54305 37111 54363 37117
rect 54305 37108 54317 37111
rect 45526 37080 54317 37108
rect 20496 37068 20502 37080
rect 54305 37077 54317 37080
rect 54351 37077 54363 37111
rect 54305 37071 54363 37077
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 5994 36864 6000 36916
rect 6052 36904 6058 36916
rect 42978 36904 42984 36916
rect 6052 36876 42984 36904
rect 6052 36864 6058 36876
rect 42978 36864 42984 36876
rect 43036 36864 43042 36916
rect 18785 36839 18843 36845
rect 18785 36805 18797 36839
rect 18831 36836 18843 36839
rect 21818 36836 21824 36848
rect 18831 36808 21824 36836
rect 18831 36805 18843 36808
rect 18785 36799 18843 36805
rect 21818 36796 21824 36808
rect 21876 36796 21882 36848
rect 23477 36839 23535 36845
rect 23477 36805 23489 36839
rect 23523 36836 23535 36839
rect 23753 36839 23811 36845
rect 23753 36836 23765 36839
rect 23523 36808 23765 36836
rect 23523 36805 23535 36808
rect 23477 36799 23535 36805
rect 23753 36805 23765 36808
rect 23799 36836 23811 36839
rect 53929 36839 53987 36845
rect 23799 36808 26234 36836
rect 23799 36805 23811 36808
rect 23753 36799 23811 36805
rect 934 36728 940 36780
rect 992 36768 998 36780
rect 1581 36771 1639 36777
rect 1581 36768 1593 36771
rect 992 36740 1593 36768
rect 992 36728 998 36740
rect 1581 36737 1593 36740
rect 1627 36737 1639 36771
rect 1581 36731 1639 36737
rect 16574 36728 16580 36780
rect 16632 36768 16638 36780
rect 18509 36771 18567 36777
rect 18509 36768 18521 36771
rect 16632 36740 18521 36768
rect 16632 36728 16638 36740
rect 18509 36737 18521 36740
rect 18555 36737 18567 36771
rect 18509 36731 18567 36737
rect 18693 36771 18751 36777
rect 18693 36737 18705 36771
rect 18739 36737 18751 36771
rect 18693 36731 18751 36737
rect 18708 36700 18736 36731
rect 18874 36728 18880 36780
rect 18932 36768 18938 36780
rect 18932 36740 19380 36768
rect 18932 36728 18938 36740
rect 19242 36700 19248 36712
rect 18708 36672 19248 36700
rect 19242 36660 19248 36672
rect 19300 36660 19306 36712
rect 19352 36700 19380 36740
rect 19426 36728 19432 36780
rect 19484 36768 19490 36780
rect 19521 36771 19579 36777
rect 19521 36768 19533 36771
rect 19484 36740 19533 36768
rect 19484 36728 19490 36740
rect 19521 36737 19533 36740
rect 19567 36737 19579 36771
rect 19521 36731 19579 36737
rect 20349 36771 20407 36777
rect 20349 36737 20361 36771
rect 20395 36768 20407 36771
rect 20714 36768 20720 36780
rect 20395 36740 20720 36768
rect 20395 36737 20407 36740
rect 20349 36731 20407 36737
rect 20364 36700 20392 36731
rect 20714 36728 20720 36740
rect 20772 36728 20778 36780
rect 20993 36771 21051 36777
rect 20993 36768 21005 36771
rect 20916 36740 21005 36768
rect 19352 36672 20392 36700
rect 19061 36635 19119 36641
rect 19061 36601 19073 36635
rect 19107 36632 19119 36635
rect 20916 36632 20944 36740
rect 20993 36737 21005 36740
rect 21039 36737 21051 36771
rect 20993 36731 21051 36737
rect 23934 36728 23940 36780
rect 23992 36768 23998 36780
rect 24029 36771 24087 36777
rect 24029 36768 24041 36771
rect 23992 36740 24041 36768
rect 23992 36728 23998 36740
rect 24029 36737 24041 36740
rect 24075 36768 24087 36771
rect 24118 36768 24124 36780
rect 24075 36740 24124 36768
rect 24075 36737 24087 36740
rect 24029 36731 24087 36737
rect 24118 36728 24124 36740
rect 24176 36728 24182 36780
rect 21085 36703 21143 36709
rect 21085 36669 21097 36703
rect 21131 36700 21143 36703
rect 21174 36700 21180 36712
rect 21131 36672 21180 36700
rect 21131 36669 21143 36672
rect 21085 36663 21143 36669
rect 21174 36660 21180 36672
rect 21232 36660 21238 36712
rect 23842 36660 23848 36712
rect 23900 36660 23906 36712
rect 26206 36700 26234 36808
rect 53929 36805 53941 36839
rect 53975 36836 53987 36839
rect 57330 36836 57336 36848
rect 53975 36808 57336 36836
rect 53975 36805 53987 36808
rect 53929 36799 53987 36805
rect 57330 36796 57336 36808
rect 57388 36796 57394 36848
rect 53650 36728 53656 36780
rect 53708 36728 53714 36780
rect 53834 36728 53840 36780
rect 53892 36728 53898 36780
rect 54026 36771 54084 36777
rect 54026 36768 54038 36771
rect 53944 36740 54038 36768
rect 39942 36700 39948 36712
rect 26206 36672 39948 36700
rect 39942 36660 39948 36672
rect 40000 36660 40006 36712
rect 53944 36700 53972 36740
rect 54026 36737 54038 36740
rect 54072 36737 54084 36771
rect 54026 36731 54084 36737
rect 53484 36672 53972 36700
rect 53484 36644 53512 36672
rect 19107 36604 20944 36632
rect 19107 36601 19119 36604
rect 19061 36595 19119 36601
rect 21818 36592 21824 36644
rect 21876 36632 21882 36644
rect 39114 36632 39120 36644
rect 21876 36604 39120 36632
rect 21876 36592 21882 36604
rect 39114 36592 39120 36604
rect 39172 36592 39178 36644
rect 40862 36592 40868 36644
rect 40920 36632 40926 36644
rect 53466 36632 53472 36644
rect 40920 36604 53472 36632
rect 40920 36592 40926 36604
rect 53466 36592 53472 36604
rect 53524 36592 53530 36644
rect 1765 36567 1823 36573
rect 1765 36533 1777 36567
rect 1811 36564 1823 36567
rect 3418 36564 3424 36576
rect 1811 36536 3424 36564
rect 1811 36533 1823 36536
rect 1765 36527 1823 36533
rect 3418 36524 3424 36536
rect 3476 36524 3482 36576
rect 20990 36524 20996 36576
rect 21048 36524 21054 36576
rect 21358 36524 21364 36576
rect 21416 36524 21422 36576
rect 23474 36524 23480 36576
rect 23532 36564 23538 36576
rect 23753 36567 23811 36573
rect 23753 36564 23765 36567
rect 23532 36536 23765 36564
rect 23532 36524 23538 36536
rect 23753 36533 23765 36536
rect 23799 36533 23811 36567
rect 23753 36527 23811 36533
rect 24213 36567 24271 36573
rect 24213 36533 24225 36567
rect 24259 36564 24271 36567
rect 24578 36564 24584 36576
rect 24259 36536 24584 36564
rect 24259 36533 24271 36536
rect 24213 36527 24271 36533
rect 24578 36524 24584 36536
rect 24636 36524 24642 36576
rect 54202 36524 54208 36576
rect 54260 36524 54266 36576
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1765 36363 1823 36369
rect 1765 36329 1777 36363
rect 1811 36360 1823 36363
rect 6730 36360 6736 36372
rect 1811 36332 6736 36360
rect 1811 36329 1823 36332
rect 1765 36323 1823 36329
rect 6730 36320 6736 36332
rect 6788 36320 6794 36372
rect 23474 36360 23480 36372
rect 6886 36332 23480 36360
rect 3053 36295 3111 36301
rect 3053 36261 3065 36295
rect 3099 36292 3111 36295
rect 6886 36292 6914 36332
rect 23474 36320 23480 36332
rect 23532 36320 23538 36372
rect 23842 36320 23848 36372
rect 23900 36320 23906 36372
rect 54202 36360 54208 36372
rect 26206 36332 54208 36360
rect 21358 36292 21364 36304
rect 3099 36264 6914 36292
rect 20180 36264 21364 36292
rect 3099 36261 3111 36264
rect 3053 36255 3111 36261
rect 2406 36184 2412 36236
rect 2464 36224 2470 36236
rect 2464 36196 2912 36224
rect 2464 36184 2470 36196
rect 2498 36116 2504 36168
rect 2556 36116 2562 36168
rect 2884 36165 2912 36196
rect 20180 36165 20208 36264
rect 21358 36252 21364 36264
rect 21416 36252 21422 36304
rect 21450 36252 21456 36304
rect 21508 36292 21514 36304
rect 26206 36292 26234 36332
rect 54202 36320 54208 36332
rect 54260 36320 54266 36372
rect 21508 36264 26234 36292
rect 21508 36252 21514 36264
rect 20257 36227 20315 36233
rect 20257 36193 20269 36227
rect 20303 36224 20315 36227
rect 20622 36224 20628 36236
rect 20303 36196 20628 36224
rect 20303 36193 20315 36196
rect 20257 36187 20315 36193
rect 20622 36184 20628 36196
rect 20680 36184 20686 36236
rect 20714 36184 20720 36236
rect 20772 36184 20778 36236
rect 22664 36196 23428 36224
rect 2874 36159 2932 36165
rect 2874 36125 2886 36159
rect 2920 36125 2932 36159
rect 2874 36119 2932 36125
rect 20165 36159 20223 36165
rect 20165 36125 20177 36159
rect 20211 36125 20223 36159
rect 20165 36119 20223 36125
rect 20441 36159 20499 36165
rect 20441 36125 20453 36159
rect 20487 36125 20499 36159
rect 20441 36119 20499 36125
rect 934 36048 940 36100
rect 992 36088 998 36100
rect 1673 36091 1731 36097
rect 1673 36088 1685 36091
rect 992 36060 1685 36088
rect 992 36048 998 36060
rect 1673 36057 1685 36060
rect 1719 36057 1731 36091
rect 1673 36051 1731 36057
rect 2222 36048 2228 36100
rect 2280 36088 2286 36100
rect 2685 36091 2743 36097
rect 2685 36088 2697 36091
rect 2280 36060 2697 36088
rect 2280 36048 2286 36060
rect 2685 36057 2697 36060
rect 2731 36057 2743 36091
rect 2685 36051 2743 36057
rect 2700 36020 2728 36051
rect 2774 36048 2780 36100
rect 2832 36048 2838 36100
rect 16666 36088 16672 36100
rect 6886 36060 16672 36088
rect 6886 36020 6914 36060
rect 16666 36048 16672 36060
rect 16724 36048 16730 36100
rect 19978 36048 19984 36100
rect 20036 36088 20042 36100
rect 20456 36088 20484 36119
rect 22278 36116 22284 36168
rect 22336 36116 22342 36168
rect 22554 36116 22560 36168
rect 22612 36116 22618 36168
rect 22664 36165 22692 36196
rect 23400 36168 23428 36196
rect 23566 36184 23572 36236
rect 23624 36224 23630 36236
rect 23624 36196 24808 36224
rect 23624 36184 23630 36196
rect 22649 36159 22707 36165
rect 22649 36125 22661 36159
rect 22695 36125 22707 36159
rect 22649 36119 22707 36125
rect 23290 36116 23296 36168
rect 23348 36116 23354 36168
rect 23382 36116 23388 36168
rect 23440 36156 23446 36168
rect 23661 36159 23719 36165
rect 23661 36156 23673 36159
rect 23440 36128 23673 36156
rect 23440 36116 23446 36128
rect 23661 36125 23673 36128
rect 23707 36156 23719 36159
rect 24302 36156 24308 36168
rect 23707 36128 24308 36156
rect 23707 36125 23719 36128
rect 23661 36119 23719 36125
rect 24302 36116 24308 36128
rect 24360 36116 24366 36168
rect 24578 36116 24584 36168
rect 24636 36116 24642 36168
rect 24780 36165 24808 36196
rect 24765 36159 24823 36165
rect 24765 36125 24777 36159
rect 24811 36125 24823 36159
rect 24765 36119 24823 36125
rect 20036 36060 20484 36088
rect 22465 36091 22523 36097
rect 20036 36048 20042 36060
rect 22465 36057 22477 36091
rect 22511 36057 22523 36091
rect 23477 36091 23535 36097
rect 23477 36088 23489 36091
rect 22465 36051 22523 36057
rect 22664 36060 23489 36088
rect 2700 35992 6914 36020
rect 22186 35980 22192 36032
rect 22244 36020 22250 36032
rect 22480 36020 22508 36051
rect 22664 36020 22692 36060
rect 23477 36057 23489 36060
rect 23523 36057 23535 36091
rect 23477 36051 23535 36057
rect 22244 35992 22692 36020
rect 22244 35980 22250 35992
rect 22738 35980 22744 36032
rect 22796 36020 22802 36032
rect 22833 36023 22891 36029
rect 22833 36020 22845 36023
rect 22796 35992 22845 36020
rect 22796 35980 22802 35992
rect 22833 35989 22845 35992
rect 22879 35989 22891 36023
rect 23492 36020 23520 36051
rect 23566 36048 23572 36100
rect 23624 36048 23630 36100
rect 25133 36091 25191 36097
rect 25133 36057 25145 36091
rect 25179 36088 25191 36091
rect 25222 36088 25228 36100
rect 25179 36060 25228 36088
rect 25179 36057 25191 36060
rect 25133 36051 25191 36057
rect 25222 36048 25228 36060
rect 25280 36048 25286 36100
rect 57974 36048 57980 36100
rect 58032 36048 58038 36100
rect 58345 36091 58403 36097
rect 58345 36057 58357 36091
rect 58391 36088 58403 36091
rect 59262 36088 59268 36100
rect 58391 36060 59268 36088
rect 58391 36057 58403 36060
rect 58345 36051 58403 36057
rect 59262 36048 59268 36060
rect 59320 36048 59326 36100
rect 24946 36020 24952 36032
rect 23492 35992 24952 36020
rect 22833 35983 22891 35989
rect 24946 35980 24952 35992
rect 25004 35980 25010 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1578 35776 1584 35828
rect 1636 35816 1642 35828
rect 1765 35819 1823 35825
rect 1765 35816 1777 35819
rect 1636 35788 1777 35816
rect 1636 35776 1642 35788
rect 1765 35785 1777 35788
rect 1811 35785 1823 35819
rect 1765 35779 1823 35785
rect 19797 35819 19855 35825
rect 19797 35785 19809 35819
rect 19843 35816 19855 35819
rect 20990 35816 20996 35828
rect 19843 35788 20996 35816
rect 19843 35785 19855 35788
rect 19797 35779 19855 35785
rect 20990 35776 20996 35788
rect 21048 35776 21054 35828
rect 25130 35776 25136 35828
rect 25188 35816 25194 35828
rect 41690 35816 41696 35828
rect 25188 35788 40448 35816
rect 25188 35776 25194 35788
rect 18782 35708 18788 35760
rect 18840 35748 18846 35760
rect 19521 35751 19579 35757
rect 19521 35748 19533 35751
rect 18840 35720 19533 35748
rect 18840 35708 18846 35720
rect 19521 35717 19533 35720
rect 19567 35717 19579 35751
rect 19521 35711 19579 35717
rect 21082 35708 21088 35760
rect 21140 35748 21146 35760
rect 40420 35757 40448 35788
rect 40512 35788 41696 35816
rect 40405 35751 40463 35757
rect 21140 35720 22094 35748
rect 21140 35708 21146 35720
rect 934 35640 940 35692
rect 992 35680 998 35692
rect 1673 35683 1731 35689
rect 1673 35680 1685 35683
rect 992 35652 1685 35680
rect 992 35640 998 35652
rect 1673 35649 1685 35652
rect 1719 35649 1731 35683
rect 1673 35643 1731 35649
rect 18874 35640 18880 35692
rect 18932 35680 18938 35692
rect 19245 35683 19303 35689
rect 19245 35680 19257 35683
rect 18932 35652 19257 35680
rect 18932 35640 18938 35652
rect 19245 35649 19257 35652
rect 19291 35649 19303 35683
rect 19245 35643 19303 35649
rect 19429 35683 19487 35689
rect 19429 35649 19441 35683
rect 19475 35649 19487 35683
rect 19429 35643 19487 35649
rect 19613 35683 19671 35689
rect 19613 35649 19625 35683
rect 19659 35680 19671 35683
rect 20162 35680 20168 35692
rect 19659 35652 20168 35680
rect 19659 35649 19671 35652
rect 19613 35643 19671 35649
rect 19444 35612 19472 35643
rect 20162 35640 20168 35652
rect 20220 35640 20226 35692
rect 22066 35680 22094 35720
rect 40405 35717 40417 35751
rect 40451 35717 40463 35751
rect 40405 35711 40463 35717
rect 40512 35689 40540 35788
rect 41690 35776 41696 35788
rect 41748 35776 41754 35828
rect 22649 35683 22707 35689
rect 22649 35680 22661 35683
rect 22066 35652 22661 35680
rect 22649 35649 22661 35652
rect 22695 35649 22707 35683
rect 22649 35643 22707 35649
rect 40221 35683 40279 35689
rect 40221 35649 40233 35683
rect 40267 35649 40279 35683
rect 40221 35643 40279 35649
rect 40497 35683 40555 35689
rect 40497 35649 40509 35683
rect 40543 35649 40555 35683
rect 40497 35643 40555 35649
rect 21082 35612 21088 35624
rect 19444 35584 21088 35612
rect 21082 35572 21088 35584
rect 21140 35572 21146 35624
rect 23382 35572 23388 35624
rect 23440 35572 23446 35624
rect 40236 35612 40264 35643
rect 40586 35640 40592 35692
rect 40644 35640 40650 35692
rect 47670 35612 47676 35624
rect 40236 35584 47676 35612
rect 47670 35572 47676 35584
rect 47728 35572 47734 35624
rect 39942 35504 39948 35556
rect 40000 35544 40006 35556
rect 40773 35547 40831 35553
rect 40773 35544 40785 35547
rect 40000 35516 40785 35544
rect 40000 35504 40006 35516
rect 40773 35513 40785 35516
rect 40819 35513 40831 35547
rect 40773 35507 40831 35513
rect 18874 35436 18880 35488
rect 18932 35436 18938 35488
rect 33778 35436 33784 35488
rect 33836 35476 33842 35488
rect 40586 35476 40592 35488
rect 33836 35448 40592 35476
rect 33836 35436 33842 35448
rect 40586 35436 40592 35448
rect 40644 35436 40650 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 22738 35232 22744 35284
rect 22796 35232 22802 35284
rect 23566 35232 23572 35284
rect 23624 35272 23630 35284
rect 37366 35272 37372 35284
rect 23624 35244 37372 35272
rect 23624 35232 23630 35244
rect 37366 35232 37372 35244
rect 37424 35232 37430 35284
rect 1857 35207 1915 35213
rect 1857 35173 1869 35207
rect 1903 35204 1915 35207
rect 2774 35204 2780 35216
rect 1903 35176 2780 35204
rect 1903 35173 1915 35176
rect 1857 35167 1915 35173
rect 2774 35164 2780 35176
rect 2832 35164 2838 35216
rect 22278 35164 22284 35216
rect 22336 35204 22342 35216
rect 55674 35204 55680 35216
rect 22336 35176 55680 35204
rect 22336 35164 22342 35176
rect 55674 35164 55680 35176
rect 55732 35164 55738 35216
rect 22649 35139 22707 35145
rect 22649 35105 22661 35139
rect 22695 35136 22707 35139
rect 22695 35108 35894 35136
rect 22695 35105 22707 35108
rect 22649 35099 22707 35105
rect 21174 35028 21180 35080
rect 21232 35068 21238 35080
rect 22741 35071 22799 35077
rect 22741 35068 22753 35071
rect 21232 35040 22753 35068
rect 21232 35028 21238 35040
rect 22741 35037 22753 35040
rect 22787 35068 22799 35071
rect 24394 35068 24400 35080
rect 22787 35040 24400 35068
rect 22787 35037 22799 35040
rect 22741 35031 22799 35037
rect 24394 35028 24400 35040
rect 24452 35068 24458 35080
rect 26970 35068 26976 35080
rect 24452 35040 26976 35068
rect 24452 35028 24458 35040
rect 26970 35028 26976 35040
rect 27028 35028 27034 35080
rect 934 34960 940 35012
rect 992 35000 998 35012
rect 1673 35003 1731 35009
rect 1673 35000 1685 35003
rect 992 34972 1685 35000
rect 992 34960 998 34972
rect 1673 34969 1685 34972
rect 1719 34969 1731 35003
rect 1673 34963 1731 34969
rect 22465 35003 22523 35009
rect 22465 34969 22477 35003
rect 22511 35000 22523 35003
rect 22646 35000 22652 35012
rect 22511 34972 22652 35000
rect 22511 34969 22523 34972
rect 22465 34963 22523 34969
rect 22646 34960 22652 34972
rect 22704 34960 22710 35012
rect 22922 34892 22928 34944
rect 22980 34892 22986 34944
rect 35866 34932 35894 35108
rect 40034 35028 40040 35080
rect 40092 35028 40098 35080
rect 40310 35028 40316 35080
rect 40368 35028 40374 35080
rect 40405 35071 40463 35077
rect 40405 35037 40417 35071
rect 40451 35068 40463 35071
rect 40494 35068 40500 35080
rect 40451 35040 40500 35068
rect 40451 35037 40463 35040
rect 40405 35031 40463 35037
rect 40494 35028 40500 35040
rect 40552 35028 40558 35080
rect 54938 35028 54944 35080
rect 54996 35068 55002 35080
rect 57885 35071 57943 35077
rect 57885 35068 57897 35071
rect 54996 35040 57897 35068
rect 54996 35028 55002 35040
rect 57885 35037 57897 35040
rect 57931 35037 57943 35071
rect 57885 35031 57943 35037
rect 37366 34960 37372 35012
rect 37424 35000 37430 35012
rect 40221 35003 40279 35009
rect 40221 35000 40233 35003
rect 37424 34972 40233 35000
rect 37424 34960 37430 34972
rect 40221 34969 40233 34972
rect 40267 34969 40279 35003
rect 40221 34963 40279 34969
rect 58158 34960 58164 35012
rect 58216 34960 58222 35012
rect 40589 34935 40647 34941
rect 40589 34932 40601 34935
rect 35866 34904 40601 34932
rect 40589 34901 40601 34904
rect 40635 34901 40647 34935
rect 40589 34895 40647 34901
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 20254 34688 20260 34740
rect 20312 34728 20318 34740
rect 22370 34728 22376 34740
rect 20312 34700 22376 34728
rect 20312 34688 20318 34700
rect 22370 34688 22376 34700
rect 22428 34688 22434 34740
rect 58253 34731 58311 34737
rect 58253 34697 58265 34731
rect 58299 34728 58311 34731
rect 59354 34728 59360 34740
rect 58299 34700 59360 34728
rect 58299 34697 58311 34700
rect 58253 34691 58311 34697
rect 59354 34688 59360 34700
rect 59412 34688 59418 34740
rect 19426 34620 19432 34672
rect 19484 34660 19490 34672
rect 24854 34660 24860 34672
rect 19484 34632 24860 34660
rect 19484 34620 19490 34632
rect 24854 34620 24860 34632
rect 24912 34620 24918 34672
rect 58069 34595 58127 34601
rect 58069 34561 58081 34595
rect 58115 34592 58127 34595
rect 58986 34592 58992 34604
rect 58115 34564 58992 34592
rect 58115 34561 58127 34564
rect 58069 34555 58127 34561
rect 58986 34552 58992 34564
rect 59044 34552 59050 34604
rect 20070 34484 20076 34536
rect 20128 34524 20134 34536
rect 23382 34524 23388 34536
rect 20128 34496 23388 34524
rect 20128 34484 20134 34496
rect 23382 34484 23388 34496
rect 23440 34484 23446 34536
rect 47578 34484 47584 34536
rect 47636 34524 47642 34536
rect 54662 34524 54668 34536
rect 47636 34496 54668 34524
rect 47636 34484 47642 34496
rect 54662 34484 54668 34496
rect 54720 34484 54726 34536
rect 40034 34416 40040 34468
rect 40092 34456 40098 34468
rect 44358 34456 44364 34468
rect 40092 34428 44364 34456
rect 40092 34416 40098 34428
rect 44358 34416 44364 34428
rect 44416 34416 44422 34468
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 21082 34144 21088 34196
rect 21140 34184 21146 34196
rect 23566 34184 23572 34196
rect 21140 34156 23572 34184
rect 21140 34144 21146 34156
rect 23566 34144 23572 34156
rect 23624 34184 23630 34196
rect 23842 34184 23848 34196
rect 23624 34156 23848 34184
rect 23624 34144 23630 34156
rect 23842 34144 23848 34156
rect 23900 34144 23906 34196
rect 40034 34144 40040 34196
rect 40092 34184 40098 34196
rect 40494 34184 40500 34196
rect 40092 34156 40500 34184
rect 40092 34144 40098 34156
rect 40494 34144 40500 34156
rect 40552 34144 40558 34196
rect 17310 34076 17316 34128
rect 17368 34116 17374 34128
rect 17368 34088 23336 34116
rect 17368 34076 17374 34088
rect 21910 34048 21916 34060
rect 21284 34020 21916 34048
rect 934 33940 940 33992
rect 992 33980 998 33992
rect 21284 33989 21312 34020
rect 21910 34008 21916 34020
rect 21968 34008 21974 34060
rect 21450 33989 21456 33992
rect 1673 33983 1731 33989
rect 1673 33980 1685 33983
rect 992 33952 1685 33980
rect 992 33940 998 33952
rect 1673 33949 1685 33952
rect 1719 33949 1731 33983
rect 1673 33943 1731 33949
rect 21269 33983 21327 33989
rect 21269 33949 21281 33983
rect 21315 33949 21327 33983
rect 21269 33943 21327 33949
rect 21417 33983 21456 33989
rect 21417 33949 21429 33983
rect 21417 33943 21456 33949
rect 21450 33940 21456 33943
rect 21508 33940 21514 33992
rect 21542 33940 21548 33992
rect 21600 33940 21606 33992
rect 21818 33989 21824 33992
rect 21775 33983 21824 33989
rect 21775 33949 21787 33983
rect 21821 33949 21824 33983
rect 21775 33943 21824 33949
rect 21818 33940 21824 33943
rect 21876 33940 21882 33992
rect 22465 33983 22523 33989
rect 22465 33949 22477 33983
rect 22511 33949 22523 33983
rect 22465 33943 22523 33949
rect 1857 33915 1915 33921
rect 1857 33881 1869 33915
rect 1903 33912 1915 33915
rect 21637 33915 21695 33921
rect 1903 33884 6914 33912
rect 1903 33881 1915 33884
rect 1857 33875 1915 33881
rect 6886 33844 6914 33884
rect 21637 33881 21649 33915
rect 21683 33881 21695 33915
rect 21637 33875 21695 33881
rect 21652 33844 21680 33875
rect 6886 33816 21680 33844
rect 21913 33847 21971 33853
rect 21913 33813 21925 33847
rect 21959 33844 21971 33847
rect 22480 33844 22508 33943
rect 22922 33940 22928 33992
rect 22980 33940 22986 33992
rect 23106 33872 23112 33924
rect 23164 33912 23170 33924
rect 23201 33915 23259 33921
rect 23201 33912 23213 33915
rect 23164 33884 23213 33912
rect 23164 33872 23170 33884
rect 23201 33881 23213 33884
rect 23247 33881 23259 33915
rect 23308 33912 23336 34088
rect 23474 34076 23480 34128
rect 23532 34116 23538 34128
rect 23532 34088 25084 34116
rect 23532 34076 23538 34088
rect 24946 34048 24952 34060
rect 24872 34020 24952 34048
rect 24486 33940 24492 33992
rect 24544 33980 24550 33992
rect 24762 33989 24768 33992
rect 24581 33983 24639 33989
rect 24581 33980 24593 33983
rect 24544 33952 24593 33980
rect 24544 33940 24550 33952
rect 24581 33949 24593 33952
rect 24627 33949 24639 33983
rect 24581 33943 24639 33949
rect 24729 33983 24768 33989
rect 24729 33949 24741 33983
rect 24729 33943 24768 33949
rect 24762 33940 24768 33943
rect 24820 33940 24826 33992
rect 24872 33989 24900 34020
rect 24946 34008 24952 34020
rect 25004 34008 25010 34060
rect 25056 33989 25084 34088
rect 24857 33983 24915 33989
rect 24857 33949 24869 33983
rect 24903 33949 24915 33983
rect 24857 33943 24915 33949
rect 25046 33983 25104 33989
rect 25046 33949 25058 33983
rect 25092 33949 25104 33983
rect 25046 33943 25104 33949
rect 24949 33915 25007 33921
rect 24949 33912 24961 33915
rect 23308 33884 24961 33912
rect 23201 33875 23259 33881
rect 24949 33881 24961 33884
rect 24995 33881 25007 33915
rect 24949 33875 25007 33881
rect 21959 33816 22508 33844
rect 21959 33813 21971 33816
rect 21913 33807 21971 33813
rect 25038 33804 25044 33856
rect 25096 33844 25102 33856
rect 25225 33847 25283 33853
rect 25225 33844 25237 33847
rect 25096 33816 25237 33844
rect 25096 33804 25102 33816
rect 25225 33813 25237 33816
rect 25271 33813 25283 33847
rect 25225 33807 25283 33813
rect 35894 33804 35900 33856
rect 35952 33844 35958 33856
rect 36538 33844 36544 33856
rect 35952 33816 36544 33844
rect 35952 33804 35958 33816
rect 36538 33804 36544 33816
rect 36596 33804 36602 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 22296 33612 23244 33640
rect 1857 33575 1915 33581
rect 1857 33541 1869 33575
rect 1903 33572 1915 33575
rect 2314 33572 2320 33584
rect 1903 33544 2320 33572
rect 1903 33541 1915 33544
rect 1857 33535 1915 33541
rect 2314 33532 2320 33544
rect 2372 33532 2378 33584
rect 12158 33532 12164 33584
rect 12216 33572 12222 33584
rect 21177 33575 21235 33581
rect 21177 33572 21189 33575
rect 12216 33544 21189 33572
rect 12216 33532 12222 33544
rect 21177 33541 21189 33544
rect 21223 33541 21235 33575
rect 21177 33535 21235 33541
rect 22296 33516 22324 33612
rect 22370 33532 22376 33584
rect 22428 33532 22434 33584
rect 23216 33572 23244 33612
rect 24854 33600 24860 33652
rect 24912 33640 24918 33652
rect 31018 33640 31024 33652
rect 24912 33612 31024 33640
rect 24912 33600 24918 33612
rect 31018 33600 31024 33612
rect 31076 33600 31082 33652
rect 38470 33640 38476 33652
rect 36004 33612 38476 33640
rect 34698 33572 34704 33584
rect 23216 33544 34704 33572
rect 34698 33532 34704 33544
rect 34756 33532 34762 33584
rect 36004 33581 36032 33612
rect 38470 33600 38476 33612
rect 38528 33600 38534 33652
rect 35989 33575 36047 33581
rect 35989 33541 36001 33575
rect 36035 33541 36047 33575
rect 35989 33535 36047 33541
rect 934 33464 940 33516
rect 992 33504 998 33516
rect 1673 33507 1731 33513
rect 1673 33504 1685 33507
rect 992 33476 1685 33504
rect 992 33464 998 33476
rect 1673 33473 1685 33476
rect 1719 33473 1731 33507
rect 1673 33467 1731 33473
rect 20898 33464 20904 33516
rect 20956 33464 20962 33516
rect 21082 33464 21088 33516
rect 21140 33464 21146 33516
rect 21266 33464 21272 33516
rect 21324 33464 21330 33516
rect 22005 33507 22063 33513
rect 22005 33504 22017 33507
rect 21468 33476 22017 33504
rect 20346 33396 20352 33448
rect 20404 33436 20410 33448
rect 20622 33436 20628 33448
rect 20404 33408 20628 33436
rect 20404 33396 20410 33408
rect 20622 33396 20628 33408
rect 20680 33396 20686 33448
rect 21468 33377 21496 33476
rect 22005 33473 22017 33476
rect 22051 33473 22063 33507
rect 22005 33467 22063 33473
rect 22153 33507 22211 33513
rect 22153 33473 22165 33507
rect 22199 33504 22211 33507
rect 22199 33473 22232 33504
rect 22153 33467 22232 33473
rect 22204 33436 22232 33467
rect 22278 33464 22284 33516
rect 22336 33464 22342 33516
rect 22511 33507 22569 33513
rect 22511 33473 22523 33507
rect 22557 33504 22569 33507
rect 23474 33504 23480 33516
rect 22557 33476 23480 33504
rect 22557 33473 22569 33476
rect 22511 33467 22569 33473
rect 23474 33464 23480 33476
rect 23532 33464 23538 33516
rect 35894 33513 35900 33516
rect 35713 33507 35771 33513
rect 35713 33504 35725 33507
rect 26206 33476 35725 33504
rect 24946 33436 24952 33448
rect 22204 33408 24952 33436
rect 24946 33396 24952 33408
rect 25004 33396 25010 33448
rect 21453 33371 21511 33377
rect 21453 33337 21465 33371
rect 21499 33337 21511 33371
rect 21453 33331 21511 33337
rect 23566 33328 23572 33380
rect 23624 33368 23630 33380
rect 26206 33368 26234 33476
rect 35713 33473 35725 33476
rect 35759 33473 35771 33507
rect 35713 33467 35771 33473
rect 35861 33507 35900 33513
rect 35861 33473 35873 33507
rect 35861 33467 35900 33473
rect 35894 33464 35900 33467
rect 35952 33464 35958 33516
rect 36004 33368 36032 33535
rect 36078 33532 36084 33584
rect 36136 33532 36142 33584
rect 36219 33507 36277 33513
rect 36219 33473 36231 33507
rect 36265 33504 36277 33507
rect 40034 33504 40040 33516
rect 36265 33476 40040 33504
rect 36265 33473 36277 33476
rect 36219 33467 36277 33473
rect 36648 33368 36676 33476
rect 40034 33464 40040 33476
rect 40092 33464 40098 33516
rect 23624 33340 26234 33368
rect 28920 33340 36032 33368
rect 36280 33340 36676 33368
rect 23624 33328 23630 33340
rect 22646 33260 22652 33312
rect 22704 33260 22710 33312
rect 23382 33260 23388 33312
rect 23440 33300 23446 33312
rect 28920 33300 28948 33340
rect 23440 33272 28948 33300
rect 23440 33260 23446 33272
rect 31018 33260 31024 33312
rect 31076 33300 31082 33312
rect 36280 33300 36308 33340
rect 31076 33272 36308 33300
rect 36357 33303 36415 33309
rect 31076 33260 31082 33272
rect 36357 33269 36369 33303
rect 36403 33300 36415 33303
rect 37826 33300 37832 33312
rect 36403 33272 37832 33300
rect 36403 33269 36415 33272
rect 36357 33263 36415 33269
rect 37826 33260 37832 33272
rect 37884 33260 37890 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 21821 33031 21879 33037
rect 21821 32997 21833 33031
rect 21867 33028 21879 33031
rect 22646 33028 22652 33040
rect 21867 33000 22652 33028
rect 21867 32997 21879 33000
rect 21821 32991 21879 32997
rect 22646 32988 22652 33000
rect 22704 32988 22710 33040
rect 58161 32963 58219 32969
rect 58161 32929 58173 32963
rect 58207 32960 58219 32963
rect 58986 32960 58992 32972
rect 58207 32932 58992 32960
rect 58207 32929 58219 32932
rect 58161 32923 58219 32929
rect 58986 32920 58992 32932
rect 59044 32920 59050 32972
rect 21726 32852 21732 32904
rect 21784 32852 21790 32904
rect 22005 32895 22063 32901
rect 22005 32861 22017 32895
rect 22051 32892 22063 32895
rect 23566 32892 23572 32904
rect 22051 32864 23572 32892
rect 22051 32861 22063 32864
rect 22005 32855 22063 32861
rect 23566 32852 23572 32864
rect 23624 32852 23630 32904
rect 57422 32852 57428 32904
rect 57480 32892 57486 32904
rect 57885 32895 57943 32901
rect 57885 32892 57897 32895
rect 57480 32864 57897 32892
rect 57480 32852 57486 32864
rect 57885 32861 57897 32864
rect 57931 32861 57943 32895
rect 57885 32855 57943 32861
rect 934 32784 940 32836
rect 992 32824 998 32836
rect 1673 32827 1731 32833
rect 1673 32824 1685 32827
rect 992 32796 1685 32824
rect 992 32784 998 32796
rect 1673 32793 1685 32796
rect 1719 32793 1731 32827
rect 1673 32787 1731 32793
rect 22465 32827 22523 32833
rect 22465 32793 22477 32827
rect 22511 32824 22523 32827
rect 22554 32824 22560 32836
rect 22511 32796 22560 32824
rect 22511 32793 22523 32796
rect 22465 32787 22523 32793
rect 22554 32784 22560 32796
rect 22612 32784 22618 32836
rect 57057 32827 57115 32833
rect 57057 32793 57069 32827
rect 57103 32824 57115 32827
rect 58986 32824 58992 32836
rect 57103 32796 58992 32824
rect 57103 32793 57115 32796
rect 57057 32787 57115 32793
rect 58986 32784 58992 32796
rect 59044 32784 59050 32836
rect 1765 32759 1823 32765
rect 1765 32725 1777 32759
rect 1811 32756 1823 32759
rect 16574 32756 16580 32768
rect 1811 32728 16580 32756
rect 1811 32725 1823 32728
rect 1765 32719 1823 32725
rect 16574 32716 16580 32728
rect 16632 32716 16638 32768
rect 54754 32716 54760 32768
rect 54812 32756 54818 32768
rect 57149 32759 57207 32765
rect 57149 32756 57161 32759
rect 54812 32728 57161 32756
rect 54812 32716 54818 32728
rect 57149 32725 57161 32728
rect 57195 32725 57207 32759
rect 57149 32719 57207 32725
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 24762 32512 24768 32564
rect 24820 32552 24826 32564
rect 54018 32552 54024 32564
rect 24820 32524 54024 32552
rect 24820 32512 24826 32524
rect 54018 32512 54024 32524
rect 54076 32512 54082 32564
rect 23290 32444 23296 32496
rect 23348 32484 23354 32496
rect 53282 32484 53288 32496
rect 23348 32456 53288 32484
rect 23348 32444 23354 32456
rect 53282 32444 53288 32456
rect 53340 32444 53346 32496
rect 934 32376 940 32428
rect 992 32416 998 32428
rect 1673 32419 1731 32425
rect 1673 32416 1685 32419
rect 992 32388 1685 32416
rect 992 32376 998 32388
rect 1673 32385 1685 32388
rect 1719 32385 1731 32419
rect 1673 32379 1731 32385
rect 1854 32376 1860 32428
rect 1912 32416 1918 32428
rect 22002 32416 22008 32428
rect 1912 32388 22008 32416
rect 1912 32376 1918 32388
rect 22002 32376 22008 32388
rect 22060 32376 22066 32428
rect 24854 32376 24860 32428
rect 24912 32376 24918 32428
rect 24949 32419 25007 32425
rect 24949 32385 24961 32419
rect 24995 32416 25007 32419
rect 25038 32416 25044 32428
rect 24995 32388 25044 32416
rect 24995 32385 25007 32388
rect 24949 32379 25007 32385
rect 25038 32376 25044 32388
rect 25096 32376 25102 32428
rect 25133 32419 25191 32425
rect 25133 32385 25145 32419
rect 25179 32416 25191 32419
rect 37550 32416 37556 32428
rect 25179 32388 37556 32416
rect 25179 32385 25191 32388
rect 25133 32379 25191 32385
rect 37550 32376 37556 32388
rect 37608 32376 37614 32428
rect 25222 32308 25228 32360
rect 25280 32348 25286 32360
rect 25317 32351 25375 32357
rect 25317 32348 25329 32351
rect 25280 32320 25329 32348
rect 25280 32308 25286 32320
rect 25317 32317 25329 32320
rect 25363 32317 25375 32351
rect 25317 32311 25375 32317
rect 1765 32215 1823 32221
rect 1765 32181 1777 32215
rect 1811 32212 1823 32215
rect 23014 32212 23020 32224
rect 1811 32184 23020 32212
rect 1811 32181 1823 32184
rect 1765 32175 1823 32181
rect 23014 32172 23020 32184
rect 23072 32172 23078 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 59538 31940 59544 31952
rect 26206 31912 59544 31940
rect 22741 31875 22799 31881
rect 22741 31841 22753 31875
rect 22787 31872 22799 31875
rect 26206 31872 26234 31912
rect 59538 31900 59544 31912
rect 59596 31900 59602 31952
rect 22787 31844 26234 31872
rect 22787 31841 22799 31844
rect 22741 31835 22799 31841
rect 16758 31764 16764 31816
rect 16816 31804 16822 31816
rect 21818 31804 21824 31816
rect 16816 31776 21824 31804
rect 16816 31764 16822 31776
rect 21818 31764 21824 31776
rect 21876 31804 21882 31816
rect 21876 31776 22968 31804
rect 21876 31764 21882 31776
rect 22940 31736 22968 31776
rect 23014 31764 23020 31816
rect 23072 31764 23078 31816
rect 23308 31813 23336 31844
rect 23201 31807 23259 31813
rect 23201 31804 23213 31807
rect 23124 31776 23213 31804
rect 23124 31736 23152 31776
rect 23201 31773 23213 31776
rect 23247 31773 23259 31807
rect 23201 31767 23259 31773
rect 23293 31807 23351 31813
rect 23293 31773 23305 31807
rect 23339 31773 23351 31807
rect 23293 31767 23351 31773
rect 23382 31764 23388 31816
rect 23440 31764 23446 31816
rect 48958 31764 48964 31816
rect 49016 31804 49022 31816
rect 57885 31807 57943 31813
rect 57885 31804 57897 31807
rect 49016 31776 57897 31804
rect 49016 31764 49022 31776
rect 57885 31773 57897 31776
rect 57931 31773 57943 31807
rect 57885 31767 57943 31773
rect 58161 31807 58219 31813
rect 58161 31773 58173 31807
rect 58207 31804 58219 31807
rect 58986 31804 58992 31816
rect 58207 31776 58992 31804
rect 58207 31773 58219 31776
rect 58161 31767 58219 31773
rect 58986 31764 58992 31776
rect 59044 31764 59050 31816
rect 22940 31708 23152 31736
rect 23566 31628 23572 31680
rect 23624 31628 23630 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 24302 31424 24308 31476
rect 24360 31424 24366 31476
rect 24854 31424 24860 31476
rect 24912 31424 24918 31476
rect 24320 31396 24348 31424
rect 24320 31368 24716 31396
rect 934 31288 940 31340
rect 992 31328 998 31340
rect 1673 31331 1731 31337
rect 1673 31328 1685 31331
rect 992 31300 1685 31328
rect 992 31288 998 31300
rect 1673 31297 1685 31300
rect 1719 31297 1731 31331
rect 1673 31291 1731 31297
rect 24210 31288 24216 31340
rect 24268 31288 24274 31340
rect 24394 31337 24400 31340
rect 24361 31331 24400 31337
rect 24361 31297 24373 31331
rect 24361 31291 24400 31297
rect 24394 31288 24400 31291
rect 24452 31288 24458 31340
rect 24688 31337 24716 31368
rect 24489 31331 24547 31337
rect 24489 31297 24501 31331
rect 24535 31297 24547 31331
rect 24489 31291 24547 31297
rect 24581 31331 24639 31337
rect 24581 31297 24593 31331
rect 24627 31297 24639 31331
rect 24581 31291 24639 31297
rect 24678 31331 24736 31337
rect 24678 31297 24690 31331
rect 24724 31297 24736 31331
rect 24678 31291 24736 31297
rect 21542 31220 21548 31272
rect 21600 31260 21606 31272
rect 23014 31260 23020 31272
rect 21600 31232 23020 31260
rect 21600 31220 21606 31232
rect 23014 31220 23020 31232
rect 23072 31260 23078 31272
rect 24504 31260 24532 31291
rect 23072 31232 24532 31260
rect 23072 31220 23078 31232
rect 24228 31204 24256 31232
rect 23474 31152 23480 31204
rect 23532 31192 23538 31204
rect 24118 31192 24124 31204
rect 23532 31164 24124 31192
rect 23532 31152 23538 31164
rect 24118 31152 24124 31164
rect 24176 31152 24182 31204
rect 24210 31152 24216 31204
rect 24268 31152 24274 31204
rect 1765 31127 1823 31133
rect 1765 31093 1777 31127
rect 1811 31124 1823 31127
rect 24596 31124 24624 31291
rect 58066 31288 58072 31340
rect 58124 31288 58130 31340
rect 24946 31152 24952 31204
rect 25004 31192 25010 31204
rect 47486 31192 47492 31204
rect 25004 31164 47492 31192
rect 25004 31152 25010 31164
rect 47486 31152 47492 31164
rect 47544 31152 47550 31204
rect 1811 31096 24624 31124
rect 1811 31093 1823 31096
rect 1765 31087 1823 31093
rect 36354 31084 36360 31136
rect 36412 31124 36418 31136
rect 58253 31127 58311 31133
rect 58253 31124 58265 31127
rect 36412 31096 58265 31124
rect 36412 31084 36418 31096
rect 58253 31093 58265 31096
rect 58299 31093 58311 31127
rect 58253 31087 58311 31093
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 24394 30880 24400 30932
rect 24452 30920 24458 30932
rect 40678 30920 40684 30932
rect 24452 30892 40684 30920
rect 24452 30880 24458 30892
rect 40678 30880 40684 30892
rect 40736 30880 40742 30932
rect 19426 30812 19432 30864
rect 19484 30852 19490 30864
rect 19521 30855 19579 30861
rect 19521 30852 19533 30855
rect 19484 30824 19533 30852
rect 19484 30812 19490 30824
rect 19521 30821 19533 30824
rect 19567 30821 19579 30855
rect 19521 30815 19579 30821
rect 34790 30784 34796 30796
rect 19444 30756 34796 30784
rect 19444 30725 19472 30756
rect 34790 30744 34796 30756
rect 34848 30744 34854 30796
rect 19429 30719 19487 30725
rect 19429 30685 19441 30719
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30685 19763 30719
rect 19705 30679 19763 30685
rect 934 30608 940 30660
rect 992 30648 998 30660
rect 1673 30651 1731 30657
rect 1673 30648 1685 30651
rect 992 30620 1685 30648
rect 992 30608 998 30620
rect 1673 30617 1685 30620
rect 1719 30617 1731 30651
rect 1673 30611 1731 30617
rect 17770 30608 17776 30660
rect 17828 30648 17834 30660
rect 19720 30648 19748 30679
rect 22830 30676 22836 30728
rect 22888 30676 22894 30728
rect 23109 30719 23167 30725
rect 23109 30716 23121 30719
rect 22940 30688 23121 30716
rect 17828 30620 19748 30648
rect 17828 30608 17834 30620
rect 22002 30608 22008 30660
rect 22060 30648 22066 30660
rect 22940 30648 22968 30688
rect 23109 30685 23121 30688
rect 23155 30685 23167 30719
rect 23109 30679 23167 30685
rect 23198 30676 23204 30728
rect 23256 30676 23262 30728
rect 22060 30620 22968 30648
rect 22060 30608 22066 30620
rect 23014 30608 23020 30660
rect 23072 30608 23078 30660
rect 1765 30583 1823 30589
rect 1765 30549 1777 30583
rect 1811 30580 1823 30583
rect 19150 30580 19156 30592
rect 1811 30552 19156 30580
rect 1811 30549 1823 30552
rect 1765 30543 1823 30549
rect 19150 30540 19156 30552
rect 19208 30540 19214 30592
rect 19889 30583 19947 30589
rect 19889 30549 19901 30583
rect 19935 30580 19947 30583
rect 19978 30580 19984 30592
rect 19935 30552 19984 30580
rect 19935 30549 19947 30552
rect 19889 30543 19947 30549
rect 19978 30540 19984 30552
rect 20036 30540 20042 30592
rect 21910 30540 21916 30592
rect 21968 30580 21974 30592
rect 23198 30580 23204 30592
rect 21968 30552 23204 30580
rect 21968 30540 21974 30552
rect 23198 30540 23204 30552
rect 23256 30540 23262 30592
rect 23382 30540 23388 30592
rect 23440 30540 23446 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 19426 30336 19432 30388
rect 19484 30336 19490 30388
rect 22830 30336 22836 30388
rect 22888 30376 22894 30388
rect 25958 30376 25964 30388
rect 22888 30348 25964 30376
rect 22888 30336 22894 30348
rect 25958 30336 25964 30348
rect 26016 30336 26022 30388
rect 19150 30268 19156 30320
rect 19208 30268 19214 30320
rect 22281 30311 22339 30317
rect 22281 30308 22293 30311
rect 19628 30280 22293 30308
rect 1581 30243 1639 30249
rect 1581 30209 1593 30243
rect 1627 30240 1639 30243
rect 9766 30240 9772 30252
rect 1627 30212 9772 30240
rect 1627 30209 1639 30212
rect 1581 30203 1639 30209
rect 9766 30200 9772 30212
rect 9824 30200 9830 30252
rect 18782 30200 18788 30252
rect 18840 30200 18846 30252
rect 18966 30249 18972 30252
rect 18933 30243 18972 30249
rect 18933 30209 18945 30243
rect 18933 30203 18972 30209
rect 18966 30200 18972 30203
rect 19024 30200 19030 30252
rect 19058 30200 19064 30252
rect 19116 30200 19122 30252
rect 19242 30200 19248 30252
rect 19300 30249 19306 30252
rect 19300 30240 19308 30249
rect 19300 30212 19345 30240
rect 19300 30203 19308 30212
rect 19300 30200 19306 30203
rect 934 30132 940 30184
rect 992 30172 998 30184
rect 1765 30175 1823 30181
rect 1765 30172 1777 30175
rect 992 30144 1777 30172
rect 992 30132 998 30144
rect 1765 30141 1777 30144
rect 1811 30141 1823 30175
rect 1765 30135 1823 30141
rect 8938 29996 8944 30048
rect 8996 30036 9002 30048
rect 19628 30036 19656 30280
rect 22281 30277 22293 30280
rect 22327 30277 22339 30311
rect 22281 30271 22339 30277
rect 23676 30280 31754 30308
rect 22005 30243 22063 30249
rect 22005 30209 22017 30243
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 22020 30172 22048 30203
rect 22186 30200 22192 30252
rect 22244 30200 22250 30252
rect 22373 30243 22431 30249
rect 22373 30209 22385 30243
rect 22419 30240 22431 30243
rect 23198 30240 23204 30252
rect 22419 30212 23204 30240
rect 22419 30209 22431 30212
rect 22373 30203 22431 30209
rect 23198 30200 23204 30212
rect 23256 30200 23262 30252
rect 23382 30200 23388 30252
rect 23440 30200 23446 30252
rect 23477 30243 23535 30249
rect 23477 30209 23489 30243
rect 23523 30240 23535 30243
rect 23566 30240 23572 30252
rect 23523 30212 23572 30240
rect 23523 30209 23535 30212
rect 23477 30203 23535 30209
rect 23566 30200 23572 30212
rect 23624 30200 23630 30252
rect 23676 30249 23704 30280
rect 23661 30243 23719 30249
rect 23661 30209 23673 30243
rect 23707 30209 23719 30243
rect 23661 30203 23719 30209
rect 23842 30200 23848 30252
rect 23900 30200 23906 30252
rect 31726 30240 31754 30280
rect 40586 30240 40592 30252
rect 31726 30212 40592 30240
rect 40586 30200 40592 30212
rect 40644 30200 40650 30252
rect 40678 30200 40684 30252
rect 40736 30240 40742 30252
rect 46474 30240 46480 30252
rect 40736 30212 46480 30240
rect 40736 30200 40742 30212
rect 46474 30200 46480 30212
rect 46532 30200 46538 30252
rect 30374 30172 30380 30184
rect 22020 30144 22094 30172
rect 22066 30104 22094 30144
rect 23400 30144 30380 30172
rect 22066 30076 23244 30104
rect 8996 30008 19656 30036
rect 22557 30039 22615 30045
rect 8996 29996 9002 30008
rect 22557 30005 22569 30039
rect 22603 30036 22615 30039
rect 22830 30036 22836 30048
rect 22603 30008 22836 30036
rect 22603 30005 22615 30008
rect 22557 29999 22615 30005
rect 22830 29996 22836 30008
rect 22888 29996 22894 30048
rect 23106 29996 23112 30048
rect 23164 29996 23170 30048
rect 23216 30036 23244 30076
rect 23400 30036 23428 30144
rect 30374 30132 30380 30144
rect 30432 30132 30438 30184
rect 23216 30008 23428 30036
rect 23569 30039 23627 30045
rect 23569 30005 23581 30039
rect 23615 30036 23627 30039
rect 23658 30036 23664 30048
rect 23615 30008 23664 30036
rect 23615 30005 23627 30008
rect 23569 29999 23627 30005
rect 23658 29996 23664 30008
rect 23716 30036 23722 30048
rect 23842 30036 23848 30048
rect 23716 30008 23848 30036
rect 23716 29996 23722 30008
rect 23842 29996 23848 30008
rect 23900 29996 23906 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 27338 29832 27344 29844
rect 6886 29804 27344 29832
rect 6362 29724 6368 29776
rect 6420 29764 6426 29776
rect 6886 29764 6914 29804
rect 27338 29792 27344 29804
rect 27396 29792 27402 29844
rect 6420 29736 6914 29764
rect 6420 29724 6426 29736
rect 18782 29724 18788 29776
rect 18840 29764 18846 29776
rect 24486 29764 24492 29776
rect 18840 29736 24492 29764
rect 18840 29724 18846 29736
rect 24486 29724 24492 29736
rect 24544 29724 24550 29776
rect 19058 29656 19064 29708
rect 19116 29696 19122 29708
rect 22186 29696 22192 29708
rect 19116 29668 22192 29696
rect 19116 29656 19122 29668
rect 22186 29656 22192 29668
rect 22244 29656 22250 29708
rect 23106 29696 23112 29708
rect 22572 29668 23112 29696
rect 1581 29631 1639 29637
rect 1581 29597 1593 29631
rect 1627 29628 1639 29631
rect 1946 29628 1952 29640
rect 1627 29600 1952 29628
rect 1627 29597 1639 29600
rect 1581 29591 1639 29597
rect 1946 29588 1952 29600
rect 2004 29588 2010 29640
rect 22572 29637 22600 29668
rect 23106 29656 23112 29668
rect 23164 29656 23170 29708
rect 23198 29656 23204 29708
rect 23256 29696 23262 29708
rect 25406 29696 25412 29708
rect 23256 29668 25412 29696
rect 23256 29656 23262 29668
rect 25406 29656 25412 29668
rect 25464 29656 25470 29708
rect 48866 29696 48872 29708
rect 26896 29668 48872 29696
rect 22557 29631 22615 29637
rect 22557 29597 22569 29631
rect 22603 29597 22615 29631
rect 22557 29591 22615 29597
rect 22646 29588 22652 29640
rect 22704 29588 22710 29640
rect 22830 29588 22836 29640
rect 22888 29588 22894 29640
rect 934 29520 940 29572
rect 992 29560 998 29572
rect 1857 29563 1915 29569
rect 1857 29560 1869 29563
rect 992 29532 1869 29560
rect 992 29520 998 29532
rect 1857 29529 1869 29532
rect 1903 29529 1915 29563
rect 1857 29523 1915 29529
rect 21450 29520 21456 29572
rect 21508 29560 21514 29572
rect 26896 29560 26924 29668
rect 48866 29656 48872 29668
rect 48924 29656 48930 29708
rect 58158 29656 58164 29708
rect 58216 29656 58222 29708
rect 27062 29588 27068 29640
rect 27120 29628 27126 29640
rect 40310 29628 40316 29640
rect 27120 29600 40316 29628
rect 27120 29588 27126 29600
rect 40310 29588 40316 29600
rect 40368 29588 40374 29640
rect 43346 29588 43352 29640
rect 43404 29628 43410 29640
rect 56042 29628 56048 29640
rect 43404 29600 56048 29628
rect 43404 29588 43410 29600
rect 56042 29588 56048 29600
rect 56100 29588 56106 29640
rect 57238 29588 57244 29640
rect 57296 29628 57302 29640
rect 57885 29631 57943 29637
rect 57885 29628 57897 29631
rect 57296 29600 57897 29628
rect 57296 29588 57302 29600
rect 57885 29597 57897 29600
rect 57931 29597 57943 29631
rect 57885 29591 57943 29597
rect 21508 29532 26924 29560
rect 57057 29563 57115 29569
rect 21508 29520 21514 29532
rect 57057 29529 57069 29563
rect 57103 29560 57115 29563
rect 58986 29560 58992 29572
rect 57103 29532 58992 29560
rect 57103 29529 57115 29532
rect 57057 29523 57115 29529
rect 58986 29520 58992 29532
rect 59044 29520 59050 29572
rect 22922 29452 22928 29504
rect 22980 29492 22986 29504
rect 23017 29495 23075 29501
rect 23017 29492 23029 29495
rect 22980 29464 23029 29492
rect 22980 29452 22986 29464
rect 23017 29461 23029 29464
rect 23063 29461 23075 29495
rect 23017 29455 23075 29461
rect 33778 29452 33784 29504
rect 33836 29492 33842 29504
rect 57149 29495 57207 29501
rect 57149 29492 57161 29495
rect 33836 29464 57161 29492
rect 33836 29452 33842 29464
rect 57149 29461 57161 29464
rect 57195 29461 57207 29495
rect 57149 29455 57207 29461
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 9766 29248 9772 29300
rect 9824 29248 9830 29300
rect 19242 29248 19248 29300
rect 19300 29288 19306 29300
rect 24302 29288 24308 29300
rect 19300 29260 24308 29288
rect 19300 29248 19306 29260
rect 24302 29248 24308 29260
rect 24360 29248 24366 29300
rect 9398 29112 9404 29164
rect 9456 29112 9462 29164
rect 9555 29155 9613 29161
rect 9555 29121 9567 29155
rect 9601 29152 9613 29155
rect 19058 29152 19064 29164
rect 9601 29124 19064 29152
rect 9601 29121 9613 29124
rect 9555 29115 9613 29121
rect 19058 29112 19064 29124
rect 19116 29112 19122 29164
rect 24486 28976 24492 29028
rect 24544 29016 24550 29028
rect 30834 29016 30840 29028
rect 24544 28988 30840 29016
rect 24544 28976 24550 28988
rect 30834 28976 30840 28988
rect 30892 28976 30898 29028
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 1670 28636 1676 28688
rect 1728 28676 1734 28688
rect 2590 28676 2596 28688
rect 1728 28648 2596 28676
rect 1728 28636 1734 28648
rect 2590 28636 2596 28648
rect 2648 28636 2654 28688
rect 934 28568 940 28620
rect 992 28608 998 28620
rect 1765 28611 1823 28617
rect 1765 28608 1777 28611
rect 992 28580 1777 28608
rect 992 28568 998 28580
rect 1765 28577 1777 28580
rect 1811 28577 1823 28611
rect 9398 28608 9404 28620
rect 1765 28571 1823 28577
rect 2516 28580 9404 28608
rect 2516 28549 2544 28580
rect 9398 28568 9404 28580
rect 9456 28568 9462 28620
rect 21634 28608 21640 28620
rect 16546 28580 21640 28608
rect 1581 28543 1639 28549
rect 1581 28509 1593 28543
rect 1627 28509 1639 28543
rect 1581 28503 1639 28509
rect 2501 28543 2559 28549
rect 2501 28509 2513 28543
rect 2547 28509 2559 28543
rect 2501 28503 2559 28509
rect 1596 28472 1624 28503
rect 2590 28500 2596 28552
rect 2648 28540 2654 28552
rect 16546 28540 16574 28580
rect 21634 28568 21640 28580
rect 21692 28568 21698 28620
rect 2648 28512 16574 28540
rect 2648 28500 2654 28512
rect 54662 28500 54668 28552
rect 54720 28540 54726 28552
rect 57885 28543 57943 28549
rect 57885 28540 57897 28543
rect 54720 28512 57897 28540
rect 54720 28500 54726 28512
rect 57885 28509 57897 28512
rect 57931 28509 57943 28543
rect 57885 28503 57943 28509
rect 2869 28475 2927 28481
rect 2869 28472 2881 28475
rect 1596 28444 2881 28472
rect 2869 28441 2881 28444
rect 2915 28441 2927 28475
rect 2869 28435 2927 28441
rect 28258 28432 28264 28484
rect 28316 28472 28322 28484
rect 49786 28472 49792 28484
rect 28316 28444 49792 28472
rect 28316 28432 28322 28444
rect 49786 28432 49792 28444
rect 49844 28432 49850 28484
rect 58158 28432 58164 28484
rect 58216 28432 58222 28484
rect 25958 28364 25964 28416
rect 26016 28404 26022 28416
rect 47394 28404 47400 28416
rect 26016 28376 47400 28404
rect 26016 28364 26022 28376
rect 47394 28364 47400 28376
rect 47452 28364 47458 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 1581 28067 1639 28073
rect 1581 28033 1593 28067
rect 1627 28064 1639 28067
rect 2314 28064 2320 28076
rect 1627 28036 2320 28064
rect 1627 28033 1639 28036
rect 1581 28027 1639 28033
rect 2314 28024 2320 28036
rect 2372 28024 2378 28076
rect 934 27956 940 28008
rect 992 27996 998 28008
rect 1765 27999 1823 28005
rect 1765 27996 1777 27999
rect 992 27968 1777 27996
rect 992 27956 998 27968
rect 1765 27965 1777 27968
rect 1811 27965 1823 27999
rect 1765 27959 1823 27965
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 34238 27548 34244 27600
rect 34296 27588 34302 27600
rect 35434 27588 35440 27600
rect 34296 27560 35440 27588
rect 34296 27548 34302 27560
rect 35434 27548 35440 27560
rect 35492 27548 35498 27600
rect 1578 27412 1584 27464
rect 1636 27412 1642 27464
rect 57977 27455 58035 27461
rect 57977 27421 57989 27455
rect 58023 27452 58035 27455
rect 58986 27452 58992 27464
rect 58023 27424 58992 27452
rect 58023 27421 58035 27424
rect 57977 27415 58035 27421
rect 58986 27412 58992 27424
rect 59044 27412 59050 27464
rect 934 27344 940 27396
rect 992 27384 998 27396
rect 1857 27387 1915 27393
rect 1857 27384 1869 27387
rect 992 27356 1869 27384
rect 992 27344 998 27356
rect 1857 27353 1869 27356
rect 1903 27353 1915 27387
rect 1857 27347 1915 27353
rect 34606 27276 34612 27328
rect 34664 27316 34670 27328
rect 58069 27319 58127 27325
rect 58069 27316 58081 27319
rect 34664 27288 58081 27316
rect 34664 27276 34670 27288
rect 58069 27285 58081 27288
rect 58115 27285 58127 27319
rect 58069 27279 58127 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 1578 27072 1584 27124
rect 1636 27112 1642 27124
rect 2869 27115 2927 27121
rect 2869 27112 2881 27115
rect 1636 27084 2881 27112
rect 1636 27072 1642 27084
rect 2869 27081 2881 27084
rect 2915 27081 2927 27115
rect 2869 27075 2927 27081
rect 6886 27084 24348 27112
rect 2406 27004 2412 27056
rect 2464 27044 2470 27056
rect 2464 27016 2636 27044
rect 2464 27004 2470 27016
rect 2608 26988 2636 27016
rect 1581 26979 1639 26985
rect 1581 26945 1593 26979
rect 1627 26976 1639 26979
rect 1670 26976 1676 26988
rect 1627 26948 1676 26976
rect 1627 26945 1639 26948
rect 1581 26939 1639 26945
rect 1670 26936 1676 26948
rect 1728 26936 1734 26988
rect 2498 26936 2504 26988
rect 2556 26936 2562 26988
rect 2590 26936 2596 26988
rect 2648 26936 2654 26988
rect 934 26868 940 26920
rect 992 26908 998 26920
rect 1765 26911 1823 26917
rect 1765 26908 1777 26911
rect 992 26880 1777 26908
rect 992 26868 998 26880
rect 1765 26877 1777 26880
rect 1811 26877 1823 26911
rect 1765 26871 1823 26877
rect 2130 26868 2136 26920
rect 2188 26908 2194 26920
rect 6886 26908 6914 27084
rect 21634 27004 21640 27056
rect 21692 27044 21698 27056
rect 23842 27044 23848 27056
rect 21692 27016 22876 27044
rect 21692 27004 21698 27016
rect 7834 26936 7840 26988
rect 7892 26976 7898 26988
rect 22741 26979 22799 26985
rect 22741 26976 22753 26979
rect 7892 26948 22753 26976
rect 7892 26936 7898 26948
rect 22741 26945 22753 26948
rect 22787 26945 22799 26979
rect 22741 26939 22799 26945
rect 22848 26908 22876 27016
rect 23492 27016 23848 27044
rect 23492 26988 23520 27016
rect 23842 27004 23848 27016
rect 23900 27004 23906 27056
rect 24320 27053 24348 27084
rect 24305 27047 24363 27053
rect 24305 27013 24317 27047
rect 24351 27013 24363 27047
rect 27062 27044 27068 27056
rect 24305 27007 24363 27013
rect 24504 27016 27068 27044
rect 23017 26979 23075 26985
rect 23017 26945 23029 26979
rect 23063 26976 23075 26979
rect 23474 26976 23480 26988
rect 23063 26948 23480 26976
rect 23063 26945 23075 26948
rect 23017 26939 23075 26945
rect 23474 26936 23480 26948
rect 23532 26936 23538 26988
rect 23658 26936 23664 26988
rect 23716 26976 23722 26988
rect 23937 26979 23995 26985
rect 23937 26976 23949 26979
rect 23716 26948 23949 26976
rect 23716 26936 23722 26948
rect 23937 26945 23949 26948
rect 23983 26945 23995 26979
rect 23937 26939 23995 26945
rect 24085 26979 24143 26985
rect 24085 26945 24097 26979
rect 24131 26976 24143 26979
rect 24131 26945 24164 26976
rect 24085 26939 24164 26945
rect 2188 26880 6914 26908
rect 22756 26880 22876 26908
rect 2188 26868 2194 26880
rect 22756 26772 22784 26880
rect 23198 26868 23204 26920
rect 23256 26868 23262 26920
rect 24136 26908 24164 26939
rect 24210 26936 24216 26988
rect 24268 26936 24274 26988
rect 24394 26936 24400 26988
rect 24452 26985 24458 26988
rect 24452 26976 24460 26985
rect 24504 26976 24532 27016
rect 27062 27004 27068 27016
rect 27120 27004 27126 27056
rect 24452 26948 24532 26976
rect 24452 26939 24460 26948
rect 24452 26936 24458 26939
rect 26878 26936 26884 26988
rect 26936 26976 26942 26988
rect 27890 26976 27896 26988
rect 26936 26948 27896 26976
rect 26936 26936 26942 26948
rect 27890 26936 27896 26948
rect 27948 26936 27954 26988
rect 24136 26880 27936 26908
rect 22833 26843 22891 26849
rect 22833 26809 22845 26843
rect 22879 26840 22891 26843
rect 24581 26843 24639 26849
rect 24581 26840 24593 26843
rect 22879 26812 24593 26840
rect 22879 26809 22891 26812
rect 22833 26803 22891 26809
rect 24581 26809 24593 26812
rect 24627 26809 24639 26843
rect 24581 26803 24639 26809
rect 24394 26772 24400 26784
rect 22756 26744 24400 26772
rect 24394 26732 24400 26744
rect 24452 26732 24458 26784
rect 27908 26772 27936 26880
rect 30374 26868 30380 26920
rect 30432 26908 30438 26920
rect 55214 26908 55220 26920
rect 30432 26880 55220 26908
rect 30432 26868 30438 26880
rect 55214 26868 55220 26880
rect 55272 26868 55278 26920
rect 48774 26772 48780 26784
rect 27908 26744 48780 26772
rect 48774 26732 48780 26744
rect 48832 26732 48838 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 23658 26528 23664 26580
rect 23716 26528 23722 26580
rect 28994 26432 29000 26444
rect 23124 26404 29000 26432
rect 23124 26373 23152 26404
rect 28994 26392 29000 26404
rect 29052 26392 29058 26444
rect 58158 26392 58164 26444
rect 58216 26392 58222 26444
rect 23109 26367 23167 26373
rect 23109 26333 23121 26367
rect 23155 26333 23167 26367
rect 23109 26327 23167 26333
rect 23382 26324 23388 26376
rect 23440 26324 23446 26376
rect 23477 26367 23535 26373
rect 23477 26333 23489 26367
rect 23523 26364 23535 26367
rect 23566 26364 23572 26376
rect 23523 26336 23572 26364
rect 23523 26333 23535 26336
rect 23477 26327 23535 26333
rect 23566 26324 23572 26336
rect 23624 26364 23630 26376
rect 24118 26364 24124 26376
rect 23624 26336 24124 26364
rect 23624 26324 23630 26336
rect 24118 26324 24124 26336
rect 24176 26324 24182 26376
rect 56318 26324 56324 26376
rect 56376 26364 56382 26376
rect 57885 26367 57943 26373
rect 57885 26364 57897 26367
rect 56376 26336 57897 26364
rect 56376 26324 56382 26336
rect 57885 26333 57897 26336
rect 57931 26333 57943 26367
rect 57885 26327 57943 26333
rect 18506 26256 18512 26308
rect 18564 26296 18570 26308
rect 23293 26299 23351 26305
rect 23293 26296 23305 26299
rect 18564 26268 23305 26296
rect 18564 26256 18570 26268
rect 23293 26265 23305 26268
rect 23339 26296 23351 26299
rect 23934 26296 23940 26308
rect 23339 26268 23940 26296
rect 23339 26265 23351 26268
rect 23293 26259 23351 26265
rect 23934 26256 23940 26268
rect 23992 26256 23998 26308
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 1581 25891 1639 25897
rect 1581 25857 1593 25891
rect 1627 25888 1639 25891
rect 1627 25860 6914 25888
rect 1627 25857 1639 25860
rect 1581 25851 1639 25857
rect 934 25780 940 25832
rect 992 25820 998 25832
rect 1765 25823 1823 25829
rect 1765 25820 1777 25823
rect 992 25792 1777 25820
rect 992 25780 998 25792
rect 1765 25789 1777 25792
rect 1811 25789 1823 25823
rect 1765 25783 1823 25789
rect 6886 25684 6914 25860
rect 9398 25848 9404 25900
rect 9456 25888 9462 25900
rect 10686 25888 10692 25900
rect 9456 25860 10692 25888
rect 9456 25848 9462 25860
rect 10686 25848 10692 25860
rect 10744 25848 10750 25900
rect 10843 25891 10901 25897
rect 10843 25857 10855 25891
rect 10889 25888 10901 25891
rect 26878 25888 26884 25900
rect 10889 25860 26884 25888
rect 10889 25857 10901 25860
rect 10843 25851 10901 25857
rect 26878 25848 26884 25860
rect 26936 25848 26942 25900
rect 58066 25848 58072 25900
rect 58124 25848 58130 25900
rect 34054 25780 34060 25832
rect 34112 25820 34118 25832
rect 39298 25820 39304 25832
rect 34112 25792 39304 25820
rect 34112 25780 34118 25792
rect 39298 25780 39304 25792
rect 39356 25780 39362 25832
rect 28994 25712 29000 25764
rect 29052 25752 29058 25764
rect 44726 25752 44732 25764
rect 29052 25724 44732 25752
rect 29052 25712 29058 25724
rect 44726 25712 44732 25724
rect 44784 25712 44790 25764
rect 10873 25687 10931 25693
rect 10873 25684 10885 25687
rect 6886 25656 10885 25684
rect 10873 25653 10885 25656
rect 10919 25653 10931 25687
rect 10873 25647 10931 25653
rect 20622 25644 20628 25696
rect 20680 25684 20686 25696
rect 47026 25684 47032 25696
rect 20680 25656 47032 25684
rect 20680 25644 20686 25656
rect 47026 25644 47032 25656
rect 47084 25644 47090 25696
rect 57974 25644 57980 25696
rect 58032 25684 58038 25696
rect 58253 25687 58311 25693
rect 58253 25684 58265 25687
rect 58032 25656 58265 25684
rect 58032 25644 58038 25656
rect 58253 25653 58265 25656
rect 58299 25653 58311 25687
rect 58253 25647 58311 25653
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 2869 25347 2927 25353
rect 2869 25344 2881 25347
rect 1596 25316 2881 25344
rect 1596 25285 1624 25316
rect 2869 25313 2881 25316
rect 2915 25313 2927 25347
rect 2869 25307 2927 25313
rect 1581 25279 1639 25285
rect 1581 25245 1593 25279
rect 1627 25245 1639 25279
rect 1581 25239 1639 25245
rect 2498 25236 2504 25288
rect 2556 25236 2562 25288
rect 2682 25285 2688 25288
rect 2655 25279 2688 25285
rect 2655 25245 2667 25279
rect 2655 25239 2688 25245
rect 2682 25236 2688 25239
rect 2740 25236 2746 25288
rect 52546 25236 52552 25288
rect 52604 25276 52610 25288
rect 57885 25279 57943 25285
rect 57885 25276 57897 25279
rect 52604 25248 57897 25276
rect 52604 25236 52610 25248
rect 57885 25245 57897 25248
rect 57931 25245 57943 25279
rect 57885 25239 57943 25245
rect 934 25168 940 25220
rect 992 25208 998 25220
rect 1857 25211 1915 25217
rect 1857 25208 1869 25211
rect 992 25180 1869 25208
rect 992 25168 998 25180
rect 1857 25177 1869 25180
rect 1903 25177 1915 25211
rect 1857 25171 1915 25177
rect 58158 25168 58164 25220
rect 58216 25168 58222 25220
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 47670 24828 47676 24880
rect 47728 24868 47734 24880
rect 48406 24868 48412 24880
rect 47728 24840 48412 24868
rect 47728 24828 47734 24840
rect 48406 24828 48412 24840
rect 48464 24828 48470 24880
rect 1581 24803 1639 24809
rect 1581 24769 1593 24803
rect 1627 24800 1639 24803
rect 2866 24800 2872 24812
rect 1627 24772 2872 24800
rect 1627 24769 1639 24772
rect 1581 24763 1639 24769
rect 2866 24760 2872 24772
rect 2924 24760 2930 24812
rect 58066 24760 58072 24812
rect 58124 24760 58130 24812
rect 934 24692 940 24744
rect 992 24732 998 24744
rect 1765 24735 1823 24741
rect 1765 24732 1777 24735
rect 992 24704 1777 24732
rect 992 24692 998 24704
rect 1765 24701 1777 24704
rect 1811 24701 1823 24735
rect 1765 24695 1823 24701
rect 38838 24556 38844 24608
rect 38896 24596 38902 24608
rect 58253 24599 58311 24605
rect 58253 24596 58265 24599
rect 38896 24568 58265 24596
rect 38896 24556 38902 24568
rect 58253 24565 58265 24568
rect 58299 24565 58311 24599
rect 58253 24559 58311 24565
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 2866 24352 2872 24404
rect 2924 24352 2930 24404
rect 24762 24352 24768 24404
rect 24820 24392 24826 24404
rect 42886 24392 42892 24404
rect 24820 24364 42892 24392
rect 24820 24352 24826 24364
rect 42886 24352 42892 24364
rect 42944 24352 42950 24404
rect 2682 24284 2688 24336
rect 2740 24324 2746 24336
rect 17678 24324 17684 24336
rect 2740 24296 17684 24324
rect 2740 24284 2746 24296
rect 17678 24284 17684 24296
rect 17736 24284 17742 24336
rect 18874 24284 18880 24336
rect 18932 24324 18938 24336
rect 39758 24324 39764 24336
rect 18932 24296 39764 24324
rect 18932 24284 18938 24296
rect 39758 24284 39764 24296
rect 39816 24284 39822 24336
rect 7926 24216 7932 24268
rect 7984 24256 7990 24268
rect 31570 24256 31576 24268
rect 7984 24228 31576 24256
rect 7984 24216 7990 24228
rect 31570 24216 31576 24228
rect 31628 24216 31634 24268
rect 36170 24216 36176 24268
rect 36228 24256 36234 24268
rect 54754 24256 54760 24268
rect 36228 24228 54760 24256
rect 36228 24216 36234 24228
rect 54754 24216 54760 24228
rect 54812 24216 54818 24268
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24188 1639 24191
rect 1627 24160 2636 24188
rect 1627 24157 1639 24160
rect 1581 24151 1639 24157
rect 934 24080 940 24132
rect 992 24120 998 24132
rect 1857 24123 1915 24129
rect 1857 24120 1869 24123
rect 992 24092 1869 24120
rect 992 24080 998 24092
rect 1857 24089 1869 24092
rect 1903 24089 1915 24123
rect 2608 24120 2636 24160
rect 2682 24148 2688 24200
rect 2740 24148 2746 24200
rect 2839 24191 2897 24197
rect 2839 24157 2851 24191
rect 2885 24188 2897 24191
rect 25590 24188 25596 24200
rect 2885 24160 25596 24188
rect 2885 24157 2897 24160
rect 2839 24151 2897 24157
rect 25590 24148 25596 24160
rect 25648 24148 25654 24200
rect 35526 24148 35532 24200
rect 35584 24188 35590 24200
rect 55858 24188 55864 24200
rect 35584 24160 55864 24188
rect 35584 24148 35590 24160
rect 55858 24148 55864 24160
rect 55916 24148 55922 24200
rect 12158 24120 12164 24132
rect 2608 24092 12164 24120
rect 1857 24083 1915 24089
rect 12158 24080 12164 24092
rect 12216 24080 12222 24132
rect 18966 24080 18972 24132
rect 19024 24120 19030 24132
rect 51810 24120 51816 24132
rect 19024 24092 51816 24120
rect 19024 24080 19030 24092
rect 51810 24080 51816 24092
rect 51868 24080 51874 24132
rect 2498 24012 2504 24064
rect 2556 24052 2562 24064
rect 2682 24052 2688 24064
rect 2556 24024 2688 24052
rect 2556 24012 2562 24024
rect 2682 24012 2688 24024
rect 2740 24052 2746 24064
rect 8938 24052 8944 24064
rect 2740 24024 8944 24052
rect 2740 24012 2746 24024
rect 8938 24012 8944 24024
rect 8996 24012 9002 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 12253 23715 12311 23721
rect 12253 23681 12265 23715
rect 12299 23712 12311 23715
rect 19426 23712 19432 23724
rect 12299 23684 19432 23712
rect 12299 23681 12311 23684
rect 12253 23675 12311 23681
rect 19426 23672 19432 23684
rect 19484 23672 19490 23724
rect 12802 23604 12808 23656
rect 12860 23644 12866 23656
rect 23566 23644 23572 23656
rect 12860 23616 23572 23644
rect 12860 23604 12866 23616
rect 23566 23604 23572 23616
rect 23624 23644 23630 23656
rect 24762 23644 24768 23656
rect 23624 23616 24768 23644
rect 23624 23604 23630 23616
rect 24762 23604 24768 23616
rect 24820 23604 24826 23656
rect 19426 23468 19432 23520
rect 19484 23508 19490 23520
rect 20438 23508 20444 23520
rect 19484 23480 20444 23508
rect 19484 23468 19490 23480
rect 20438 23468 20444 23480
rect 20496 23468 20502 23520
rect 27982 23468 27988 23520
rect 28040 23508 28046 23520
rect 34606 23508 34612 23520
rect 28040 23480 34612 23508
rect 28040 23468 28046 23480
rect 34606 23468 34612 23480
rect 34664 23468 34670 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 12158 23264 12164 23316
rect 12216 23264 12222 23316
rect 934 23128 940 23180
rect 992 23168 998 23180
rect 1765 23171 1823 23177
rect 1765 23168 1777 23171
rect 992 23140 1777 23168
rect 992 23128 998 23140
rect 1765 23137 1777 23140
rect 1811 23137 1823 23171
rect 11241 23171 11299 23177
rect 11241 23168 11253 23171
rect 1765 23131 1823 23137
rect 6886 23140 11253 23168
rect 1581 23103 1639 23109
rect 1581 23069 1593 23103
rect 1627 23100 1639 23103
rect 6886 23100 6914 23140
rect 11241 23137 11253 23140
rect 11287 23137 11299 23171
rect 11241 23131 11299 23137
rect 11900 23140 22094 23168
rect 1627 23072 6914 23100
rect 1627 23069 1639 23072
rect 1581 23063 1639 23069
rect 10134 23060 10140 23112
rect 10192 23100 10198 23112
rect 10686 23100 10692 23112
rect 10192 23072 10692 23100
rect 10192 23060 10198 23072
rect 10686 23060 10692 23072
rect 10744 23100 10750 23112
rect 10873 23103 10931 23109
rect 10873 23100 10885 23103
rect 10744 23072 10885 23100
rect 10744 23060 10750 23072
rect 10873 23069 10885 23072
rect 10919 23069 10931 23103
rect 10873 23063 10931 23069
rect 11027 23103 11085 23109
rect 11027 23069 11039 23103
rect 11073 23100 11085 23103
rect 11900 23100 11928 23140
rect 11073 23072 11928 23100
rect 11977 23103 12035 23109
rect 11073 23069 11085 23072
rect 11027 23063 11085 23069
rect 11977 23069 11989 23103
rect 12023 23069 12035 23103
rect 11977 23063 12035 23069
rect 12131 23103 12189 23109
rect 12131 23069 12143 23103
rect 12177 23100 12189 23103
rect 12802 23100 12808 23112
rect 12177 23072 12808 23100
rect 12177 23069 12189 23072
rect 12131 23063 12189 23069
rect 10888 23032 10916 23063
rect 11992 23032 12020 23063
rect 12802 23060 12808 23072
rect 12860 23060 12866 23112
rect 22066 23100 22094 23140
rect 25590 23128 25596 23180
rect 25648 23168 25654 23180
rect 29270 23168 29276 23180
rect 25648 23140 29276 23168
rect 25648 23128 25654 23140
rect 29270 23128 29276 23140
rect 29328 23128 29334 23180
rect 58161 23171 58219 23177
rect 58161 23137 58173 23171
rect 58207 23168 58219 23171
rect 58986 23168 58992 23180
rect 58207 23140 58992 23168
rect 58207 23137 58219 23140
rect 58161 23131 58219 23137
rect 58986 23128 58992 23140
rect 59044 23128 59050 23180
rect 24210 23100 24216 23112
rect 22066 23072 24216 23100
rect 24210 23060 24216 23072
rect 24268 23100 24274 23112
rect 25866 23100 25872 23112
rect 24268 23072 25872 23100
rect 24268 23060 24274 23072
rect 25866 23060 25872 23072
rect 25924 23060 25930 23112
rect 57882 23060 57888 23112
rect 57940 23060 57946 23112
rect 10888 23004 12020 23032
rect 22462 22992 22468 23044
rect 22520 23032 22526 23044
rect 33778 23032 33784 23044
rect 22520 23004 33784 23032
rect 22520 22992 22526 23004
rect 33778 22992 33784 23004
rect 33836 22992 33842 23044
rect 20898 22924 20904 22976
rect 20956 22964 20962 22976
rect 39482 22964 39488 22976
rect 20956 22936 39488 22964
rect 20956 22924 20962 22936
rect 39482 22924 39488 22936
rect 39540 22924 39546 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 33778 22720 33784 22772
rect 33836 22760 33842 22772
rect 59170 22760 59176 22772
rect 33836 22732 59176 22760
rect 33836 22720 33842 22732
rect 59170 22720 59176 22732
rect 59228 22720 59234 22772
rect 58158 22652 58164 22704
rect 58216 22652 58222 22704
rect 1581 22627 1639 22633
rect 1581 22593 1593 22627
rect 1627 22624 1639 22627
rect 9766 22624 9772 22636
rect 1627 22596 9772 22624
rect 1627 22593 1639 22596
rect 1581 22587 1639 22593
rect 9766 22584 9772 22596
rect 9824 22584 9830 22636
rect 17221 22627 17279 22633
rect 17221 22593 17233 22627
rect 17267 22593 17279 22627
rect 17221 22587 17279 22593
rect 17405 22627 17463 22633
rect 17405 22593 17417 22627
rect 17451 22624 17463 22627
rect 18046 22624 18052 22636
rect 17451 22596 18052 22624
rect 17451 22593 17463 22596
rect 17405 22587 17463 22593
rect 934 22516 940 22568
rect 992 22556 998 22568
rect 1765 22559 1823 22565
rect 1765 22556 1777 22559
rect 992 22528 1777 22556
rect 992 22516 998 22528
rect 1765 22525 1777 22528
rect 1811 22525 1823 22559
rect 17236 22556 17264 22587
rect 18046 22584 18052 22596
rect 18104 22584 18110 22636
rect 18782 22556 18788 22568
rect 17236 22528 18788 22556
rect 1765 22519 1823 22525
rect 18782 22516 18788 22528
rect 18840 22516 18846 22568
rect 16942 22380 16948 22432
rect 17000 22420 17006 22432
rect 17221 22423 17279 22429
rect 17221 22420 17233 22423
rect 17000 22392 17233 22420
rect 17000 22380 17006 22392
rect 17221 22389 17233 22392
rect 17267 22389 17279 22423
rect 17221 22383 17279 22389
rect 41966 22380 41972 22432
rect 42024 22420 42030 22432
rect 58253 22423 58311 22429
rect 58253 22420 58265 22423
rect 42024 22392 58265 22420
rect 42024 22380 42030 22392
rect 58253 22389 58265 22392
rect 58299 22389 58311 22423
rect 58253 22383 58311 22389
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 18874 22216 18880 22228
rect 9646 22188 18880 22216
rect 1581 22015 1639 22021
rect 1581 21981 1593 22015
rect 1627 22012 1639 22015
rect 6822 22012 6828 22024
rect 1627 21984 6828 22012
rect 1627 21981 1639 21984
rect 1581 21975 1639 21981
rect 6822 21972 6828 21984
rect 6880 21972 6886 22024
rect 9401 22015 9459 22021
rect 9401 21981 9413 22015
rect 9447 21981 9459 22015
rect 9401 21975 9459 21981
rect 9555 22015 9613 22021
rect 9555 21981 9567 22015
rect 9601 22012 9613 22015
rect 9646 22012 9674 22188
rect 18874 22176 18880 22188
rect 18932 22176 18938 22228
rect 17221 22151 17279 22157
rect 17221 22117 17233 22151
rect 17267 22117 17279 22151
rect 17221 22111 17279 22117
rect 9766 22040 9772 22092
rect 9824 22040 9830 22092
rect 9601 21984 9674 22012
rect 17037 22015 17095 22021
rect 9601 21981 9613 21984
rect 9555 21975 9613 21981
rect 17037 21981 17049 22015
rect 17083 21981 17095 22015
rect 17236 22012 17264 22111
rect 17954 22108 17960 22160
rect 18012 22108 18018 22160
rect 36630 22108 36636 22160
rect 36688 22148 36694 22160
rect 39574 22148 39580 22160
rect 36688 22120 39580 22148
rect 36688 22108 36694 22120
rect 39574 22108 39580 22120
rect 39632 22108 39638 22160
rect 17310 22040 17316 22092
rect 17368 22080 17374 22092
rect 21358 22080 21364 22092
rect 17368 22052 21364 22080
rect 17368 22040 17374 22052
rect 21358 22040 21364 22052
rect 21416 22040 21422 22092
rect 57054 22040 57060 22092
rect 57112 22080 57118 22092
rect 57422 22080 57428 22092
rect 57112 22052 57428 22080
rect 57112 22040 57118 22052
rect 57422 22040 57428 22052
rect 57480 22040 57486 22092
rect 17773 22015 17831 22021
rect 17773 22012 17785 22015
rect 17236 21984 17785 22012
rect 17037 21975 17095 21981
rect 17773 21981 17785 21984
rect 17819 21981 17831 22015
rect 17773 21975 17831 21981
rect 934 21904 940 21956
rect 992 21944 998 21956
rect 1857 21947 1915 21953
rect 1857 21944 1869 21947
rect 992 21916 1869 21944
rect 992 21904 998 21916
rect 1857 21913 1869 21916
rect 1903 21913 1915 21947
rect 9416 21944 9444 21975
rect 10134 21944 10140 21956
rect 9416 21916 10140 21944
rect 1857 21907 1915 21913
rect 10134 21904 10140 21916
rect 10192 21904 10198 21956
rect 17052 21944 17080 21975
rect 17862 21972 17868 22024
rect 17920 22012 17926 22024
rect 18509 22015 18567 22021
rect 17920 21984 18092 22012
rect 17920 21972 17926 21984
rect 17402 21944 17408 21956
rect 17052 21916 17408 21944
rect 17402 21904 17408 21916
rect 17460 21904 17466 21956
rect 18064 21876 18092 21984
rect 18509 21981 18521 22015
rect 18555 22012 18567 22015
rect 21082 22012 21088 22024
rect 18555 21984 21088 22012
rect 18555 21981 18567 21984
rect 18509 21975 18567 21981
rect 21082 21972 21088 21984
rect 21140 21972 21146 22024
rect 57146 21972 57152 22024
rect 57204 22012 57210 22024
rect 57885 22015 57943 22021
rect 57885 22012 57897 22015
rect 57204 21984 57897 22012
rect 57204 21972 57210 21984
rect 57885 21981 57897 21984
rect 57931 21981 57943 22015
rect 57885 21975 57943 21981
rect 18874 21904 18880 21956
rect 18932 21944 18938 21956
rect 22738 21944 22744 21956
rect 18932 21916 22744 21944
rect 18932 21904 18938 21916
rect 22738 21904 22744 21916
rect 22796 21944 22802 21956
rect 23290 21944 23296 21956
rect 22796 21916 23296 21944
rect 22796 21904 22802 21916
rect 23290 21904 23296 21916
rect 23348 21904 23354 21956
rect 58158 21904 58164 21956
rect 58216 21904 58222 21956
rect 18693 21879 18751 21885
rect 18693 21876 18705 21879
rect 18064 21848 18705 21876
rect 18693 21845 18705 21848
rect 18739 21845 18751 21879
rect 18693 21839 18751 21845
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 6822 21632 6828 21684
rect 6880 21672 6886 21684
rect 11057 21675 11115 21681
rect 11057 21672 11069 21675
rect 6880 21644 11069 21672
rect 6880 21632 6886 21644
rect 11057 21641 11069 21644
rect 11103 21641 11115 21675
rect 18509 21675 18567 21681
rect 18509 21672 18521 21675
rect 11057 21635 11115 21641
rect 18064 21644 18521 21672
rect 15654 21604 15660 21616
rect 12406 21576 15660 21604
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 6086 21536 6092 21548
rect 1719 21508 6092 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 6086 21496 6092 21508
rect 6144 21496 6150 21548
rect 10134 21496 10140 21548
rect 10192 21536 10198 21548
rect 10689 21539 10747 21545
rect 10689 21536 10701 21539
rect 10192 21508 10701 21536
rect 10192 21496 10198 21508
rect 10689 21505 10701 21508
rect 10735 21505 10747 21539
rect 10689 21499 10747 21505
rect 10843 21539 10901 21545
rect 10843 21505 10855 21539
rect 10889 21536 10901 21539
rect 12406 21536 12434 21576
rect 15654 21564 15660 21576
rect 15712 21564 15718 21616
rect 17862 21604 17868 21616
rect 16040 21576 17868 21604
rect 10889 21508 12434 21536
rect 10889 21505 10901 21508
rect 10843 21499 10901 21505
rect 14090 21496 14096 21548
rect 14148 21536 14154 21548
rect 16040 21545 16068 21576
rect 17862 21564 17868 21576
rect 17920 21564 17926 21616
rect 16025 21539 16083 21545
rect 16025 21536 16037 21539
rect 14148 21508 16037 21536
rect 14148 21496 14154 21508
rect 16025 21505 16037 21508
rect 16071 21505 16083 21539
rect 16025 21499 16083 21505
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21536 17095 21539
rect 18064 21536 18092 21644
rect 18509 21641 18521 21644
rect 18555 21672 18567 21675
rect 19245 21675 19303 21681
rect 18555 21644 19196 21672
rect 18555 21641 18567 21644
rect 18509 21635 18567 21641
rect 18230 21564 18236 21616
rect 18288 21604 18294 21616
rect 18288 21576 18644 21604
rect 18288 21564 18294 21576
rect 17083 21508 18092 21536
rect 17083 21505 17095 21508
rect 17037 21499 17095 21505
rect 18322 21496 18328 21548
rect 18380 21496 18386 21548
rect 18616 21545 18644 21576
rect 18601 21539 18659 21545
rect 18601 21505 18613 21539
rect 18647 21505 18659 21539
rect 18601 21499 18659 21505
rect 19061 21539 19119 21545
rect 19061 21505 19073 21539
rect 19107 21505 19119 21539
rect 19061 21499 19119 21505
rect 15378 21428 15384 21480
rect 15436 21468 15442 21480
rect 16945 21471 17003 21477
rect 16945 21468 16957 21471
rect 15436 21440 16957 21468
rect 15436 21428 15442 21440
rect 16945 21437 16957 21440
rect 16991 21437 17003 21471
rect 16945 21431 17003 21437
rect 16390 21360 16396 21412
rect 16448 21400 16454 21412
rect 16960 21400 16988 21431
rect 17402 21428 17408 21480
rect 17460 21428 17466 21480
rect 19076 21468 19104 21499
rect 18340 21440 19104 21468
rect 19168 21468 19196 21644
rect 19245 21641 19257 21675
rect 19291 21641 19303 21675
rect 19245 21635 19303 21641
rect 19260 21604 19288 21635
rect 21634 21632 21640 21684
rect 21692 21672 21698 21684
rect 23753 21675 23811 21681
rect 23753 21672 23765 21675
rect 21692 21644 23765 21672
rect 21692 21632 21698 21644
rect 23753 21641 23765 21644
rect 23799 21641 23811 21675
rect 23753 21635 23811 21641
rect 28813 21675 28871 21681
rect 28813 21641 28825 21675
rect 28859 21641 28871 21675
rect 28813 21635 28871 21641
rect 19260 21576 20024 21604
rect 19610 21496 19616 21548
rect 19668 21536 19674 21548
rect 19996 21545 20024 21576
rect 20898 21564 20904 21616
rect 20956 21604 20962 21616
rect 21818 21604 21824 21616
rect 20956 21576 21824 21604
rect 20956 21564 20962 21576
rect 21818 21564 21824 21576
rect 21876 21564 21882 21616
rect 28828 21604 28856 21635
rect 22848 21576 28856 21604
rect 19797 21539 19855 21545
rect 19797 21536 19809 21539
rect 19668 21508 19809 21536
rect 19668 21496 19674 21508
rect 19797 21505 19809 21508
rect 19843 21505 19855 21539
rect 19797 21499 19855 21505
rect 19981 21539 20039 21545
rect 19981 21505 19993 21539
rect 20027 21505 20039 21539
rect 19981 21499 20039 21505
rect 20254 21496 20260 21548
rect 20312 21536 20318 21548
rect 20717 21539 20775 21545
rect 20717 21536 20729 21539
rect 20312 21508 20729 21536
rect 20312 21496 20318 21508
rect 20717 21505 20729 21508
rect 20763 21505 20775 21539
rect 20717 21499 20775 21505
rect 20806 21496 20812 21548
rect 20864 21536 20870 21548
rect 22848 21545 22876 21576
rect 22833 21539 22891 21545
rect 22833 21536 22845 21539
rect 20864 21508 22845 21536
rect 20864 21496 20870 21508
rect 22833 21505 22845 21508
rect 22879 21505 22891 21539
rect 22833 21499 22891 21505
rect 23566 21496 23572 21548
rect 23624 21496 23630 21548
rect 24305 21539 24363 21545
rect 24305 21505 24317 21539
rect 24351 21505 24363 21539
rect 24305 21499 24363 21505
rect 19242 21468 19248 21480
rect 19168 21440 19248 21468
rect 18230 21400 18236 21412
rect 16448 21372 16896 21400
rect 16960 21372 18236 21400
rect 16448 21360 16454 21372
rect 934 21292 940 21344
rect 992 21332 998 21344
rect 1765 21335 1823 21341
rect 1765 21332 1777 21335
rect 992 21304 1777 21332
rect 992 21292 998 21304
rect 1765 21301 1777 21304
rect 1811 21301 1823 21335
rect 1765 21295 1823 21301
rect 13262 21292 13268 21344
rect 13320 21332 13326 21344
rect 16209 21335 16267 21341
rect 16209 21332 16221 21335
rect 13320 21304 16221 21332
rect 13320 21292 13326 21304
rect 16209 21301 16221 21304
rect 16255 21301 16267 21335
rect 16209 21295 16267 21301
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 16758 21332 16764 21344
rect 16632 21304 16764 21332
rect 16632 21292 16638 21304
rect 16758 21292 16764 21304
rect 16816 21292 16822 21344
rect 16868 21332 16896 21372
rect 18230 21360 18236 21372
rect 18288 21360 18294 21412
rect 18340 21409 18368 21440
rect 19242 21428 19248 21440
rect 19300 21468 19306 21480
rect 24320 21468 24348 21499
rect 25958 21496 25964 21548
rect 26016 21496 26022 21548
rect 28626 21496 28632 21548
rect 28684 21496 28690 21548
rect 34790 21496 34796 21548
rect 34848 21536 34854 21548
rect 38749 21539 38807 21545
rect 38749 21536 38761 21539
rect 34848 21508 38761 21536
rect 34848 21496 34854 21508
rect 38749 21505 38761 21508
rect 38795 21505 38807 21539
rect 38749 21499 38807 21505
rect 38841 21539 38899 21545
rect 38841 21505 38853 21539
rect 38887 21536 38899 21539
rect 39022 21536 39028 21548
rect 38887 21508 39028 21536
rect 38887 21505 38899 21508
rect 38841 21499 38899 21505
rect 28902 21468 28908 21480
rect 19300 21440 23060 21468
rect 24320 21440 28908 21468
rect 19300 21428 19306 21440
rect 18325 21403 18383 21409
rect 18325 21369 18337 21403
rect 18371 21369 18383 21403
rect 18325 21363 18383 21369
rect 21358 21360 21364 21412
rect 21416 21400 21422 21412
rect 23032 21409 23060 21440
rect 28902 21428 28908 21440
rect 28960 21428 28966 21480
rect 23017 21403 23075 21409
rect 21416 21372 22094 21400
rect 21416 21360 21422 21372
rect 19702 21332 19708 21344
rect 16868 21304 19708 21332
rect 19702 21292 19708 21304
rect 19760 21292 19766 21344
rect 19797 21335 19855 21341
rect 19797 21301 19809 21335
rect 19843 21332 19855 21335
rect 20162 21332 20168 21344
rect 19843 21304 20168 21332
rect 19843 21301 19855 21304
rect 19797 21295 19855 21301
rect 20162 21292 20168 21304
rect 20220 21292 20226 21344
rect 20714 21292 20720 21344
rect 20772 21332 20778 21344
rect 20901 21335 20959 21341
rect 20901 21332 20913 21335
rect 20772 21304 20913 21332
rect 20772 21292 20778 21304
rect 20901 21301 20913 21304
rect 20947 21301 20959 21335
rect 22066 21332 22094 21372
rect 23017 21369 23029 21403
rect 23063 21369 23075 21403
rect 24489 21403 24547 21409
rect 24489 21400 24501 21403
rect 23017 21363 23075 21369
rect 23124 21372 24501 21400
rect 23124 21332 23152 21372
rect 24489 21369 24501 21372
rect 24535 21369 24547 21403
rect 24489 21363 24547 21369
rect 26418 21360 26424 21412
rect 26476 21400 26482 21412
rect 38764 21400 38792 21499
rect 39022 21496 39028 21508
rect 39080 21496 39086 21548
rect 42797 21539 42855 21545
rect 42797 21505 42809 21539
rect 42843 21536 42855 21539
rect 43714 21536 43720 21548
rect 42843 21508 43720 21536
rect 42843 21505 42855 21508
rect 42797 21499 42855 21505
rect 43714 21496 43720 21508
rect 43772 21496 43778 21548
rect 58066 21496 58072 21548
rect 58124 21496 58130 21548
rect 38933 21471 38991 21477
rect 38933 21437 38945 21471
rect 38979 21468 38991 21471
rect 39206 21468 39212 21480
rect 38979 21440 39212 21468
rect 38979 21437 38991 21440
rect 38933 21431 38991 21437
rect 39206 21428 39212 21440
rect 39264 21468 39270 21480
rect 42242 21468 42248 21480
rect 39264 21440 42248 21468
rect 39264 21428 39270 21440
rect 42242 21428 42248 21440
rect 42300 21428 42306 21480
rect 42334 21428 42340 21480
rect 42392 21468 42398 21480
rect 42613 21471 42671 21477
rect 42613 21468 42625 21471
rect 42392 21440 42625 21468
rect 42392 21428 42398 21440
rect 42613 21437 42625 21440
rect 42659 21437 42671 21471
rect 42613 21431 42671 21437
rect 57698 21428 57704 21480
rect 57756 21468 57762 21480
rect 57882 21468 57888 21480
rect 57756 21440 57888 21468
rect 57756 21428 57762 21440
rect 57882 21428 57888 21440
rect 57940 21428 57946 21480
rect 40034 21400 40040 21412
rect 26476 21372 31754 21400
rect 38764 21372 40040 21400
rect 26476 21360 26482 21372
rect 22066 21304 23152 21332
rect 20901 21295 20959 21301
rect 23290 21292 23296 21344
rect 23348 21332 23354 21344
rect 26145 21335 26203 21341
rect 26145 21332 26157 21335
rect 23348 21304 26157 21332
rect 23348 21292 23354 21304
rect 26145 21301 26157 21304
rect 26191 21301 26203 21335
rect 31726 21332 31754 21372
rect 40034 21360 40040 21372
rect 40092 21360 40098 21412
rect 33318 21332 33324 21344
rect 31726 21304 33324 21332
rect 26145 21295 26203 21301
rect 33318 21292 33324 21304
rect 33376 21292 33382 21344
rect 38381 21335 38439 21341
rect 38381 21301 38393 21335
rect 38427 21332 38439 21335
rect 38562 21332 38568 21344
rect 38427 21304 38568 21332
rect 38427 21301 38439 21304
rect 38381 21295 38439 21301
rect 38562 21292 38568 21304
rect 38620 21292 38626 21344
rect 42978 21292 42984 21344
rect 43036 21292 43042 21344
rect 49050 21292 49056 21344
rect 49108 21332 49114 21344
rect 57882 21332 57888 21344
rect 49108 21304 57888 21332
rect 49108 21292 49114 21304
rect 57882 21292 57888 21304
rect 57940 21292 57946 21344
rect 58250 21292 58256 21344
rect 58308 21292 58314 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 13170 21088 13176 21140
rect 13228 21128 13234 21140
rect 17310 21128 17316 21140
rect 13228 21100 17316 21128
rect 13228 21088 13234 21100
rect 17310 21088 17316 21100
rect 17368 21088 17374 21140
rect 18230 21088 18236 21140
rect 18288 21128 18294 21140
rect 18417 21131 18475 21137
rect 18417 21128 18429 21131
rect 18288 21100 18429 21128
rect 18288 21088 18294 21100
rect 18417 21097 18429 21100
rect 18463 21097 18475 21131
rect 18417 21091 18475 21097
rect 19610 21088 19616 21140
rect 19668 21088 19674 21140
rect 19720 21100 20484 21128
rect 12253 21063 12311 21069
rect 12253 21029 12265 21063
rect 12299 21060 12311 21063
rect 12299 21032 12434 21060
rect 12299 21029 12311 21032
rect 12253 21023 12311 21029
rect 11882 20884 11888 20936
rect 11940 20924 11946 20936
rect 12069 20927 12127 20933
rect 12069 20924 12081 20927
rect 11940 20896 12081 20924
rect 11940 20884 11946 20896
rect 12069 20893 12081 20896
rect 12115 20893 12127 20927
rect 12406 20924 12434 21032
rect 15194 21020 15200 21072
rect 15252 21060 15258 21072
rect 16761 21063 16819 21069
rect 16761 21060 16773 21063
rect 15252 21032 16773 21060
rect 15252 21020 15258 21032
rect 16761 21029 16773 21032
rect 16807 21029 16819 21063
rect 16761 21023 16819 21029
rect 18138 21020 18144 21072
rect 18196 21060 18202 21072
rect 19720 21060 19748 21100
rect 18196 21032 19748 21060
rect 20349 21063 20407 21069
rect 18196 21020 18202 21032
rect 20349 21029 20361 21063
rect 20395 21029 20407 21063
rect 20456 21060 20484 21100
rect 21082 21088 21088 21140
rect 21140 21088 21146 21140
rect 23566 21088 23572 21140
rect 23624 21128 23630 21140
rect 26053 21131 26111 21137
rect 26053 21128 26065 21131
rect 23624 21100 26065 21128
rect 23624 21088 23630 21100
rect 26053 21097 26065 21100
rect 26099 21097 26111 21131
rect 26053 21091 26111 21097
rect 26142 21088 26148 21140
rect 26200 21128 26206 21140
rect 26200 21100 28120 21128
rect 26200 21088 26206 21100
rect 23937 21063 23995 21069
rect 23937 21060 23949 21063
rect 20456 21032 22094 21060
rect 20349 21023 20407 21029
rect 20364 20992 20392 21023
rect 17328 20964 20392 20992
rect 12805 20927 12863 20933
rect 12805 20924 12817 20927
rect 12406 20896 12817 20924
rect 12069 20887 12127 20893
rect 12805 20893 12817 20896
rect 12851 20893 12863 20927
rect 12805 20887 12863 20893
rect 14274 20884 14280 20936
rect 14332 20884 14338 20936
rect 15197 20927 15255 20933
rect 15197 20893 15209 20927
rect 15243 20893 15255 20927
rect 15197 20887 15255 20893
rect 15212 20856 15240 20887
rect 15378 20884 15384 20936
rect 15436 20884 15442 20936
rect 15841 20927 15899 20933
rect 15841 20893 15853 20927
rect 15887 20924 15899 20927
rect 16577 20927 16635 20933
rect 15887 20896 16528 20924
rect 15887 20893 15899 20896
rect 15841 20887 15899 20893
rect 16206 20856 16212 20868
rect 15212 20828 16212 20856
rect 16206 20816 16212 20828
rect 16264 20816 16270 20868
rect 16500 20856 16528 20896
rect 16577 20893 16589 20927
rect 16623 20924 16635 20927
rect 17218 20924 17224 20936
rect 16623 20896 17224 20924
rect 16623 20893 16635 20896
rect 16577 20887 16635 20893
rect 17218 20884 17224 20896
rect 17276 20884 17282 20936
rect 17328 20933 17356 20964
rect 17313 20927 17371 20933
rect 17313 20893 17325 20927
rect 17359 20893 17371 20927
rect 17313 20887 17371 20893
rect 18138 20884 18144 20936
rect 18196 20884 18202 20936
rect 18233 20927 18291 20933
rect 18233 20893 18245 20927
rect 18279 20924 18291 20927
rect 18782 20924 18788 20936
rect 18279 20896 18788 20924
rect 18279 20893 18291 20896
rect 18233 20887 18291 20893
rect 18782 20884 18788 20896
rect 18840 20884 18846 20936
rect 19426 20884 19432 20936
rect 19484 20884 19490 20936
rect 20162 20884 20168 20936
rect 20220 20884 20226 20936
rect 20898 20884 20904 20936
rect 20956 20884 20962 20936
rect 21634 20884 21640 20936
rect 21692 20884 21698 20936
rect 22066 20924 22094 21032
rect 23584 21032 23949 21060
rect 23584 20924 23612 21032
rect 23937 21029 23949 21032
rect 23983 21029 23995 21063
rect 25682 21060 25688 21072
rect 23937 21023 23995 21029
rect 24504 21032 25688 21060
rect 22066 20896 23612 20924
rect 23753 20927 23811 20933
rect 23753 20893 23765 20927
rect 23799 20924 23811 20927
rect 23842 20924 23848 20936
rect 23799 20896 23848 20924
rect 23799 20893 23811 20896
rect 23753 20887 23811 20893
rect 23842 20884 23848 20896
rect 23900 20884 23906 20936
rect 24504 20924 24532 21032
rect 25682 21020 25688 21032
rect 25740 21020 25746 21072
rect 27433 21063 27491 21069
rect 27433 21060 27445 21063
rect 26712 21032 27445 21060
rect 26418 20952 26424 21004
rect 26476 20952 26482 21004
rect 24581 20927 24639 20933
rect 24581 20924 24593 20927
rect 24504 20896 24593 20924
rect 24581 20893 24593 20896
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20924 24823 20927
rect 25590 20924 25596 20936
rect 24811 20896 25596 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 25590 20884 25596 20896
rect 25648 20884 25654 20936
rect 25774 20884 25780 20936
rect 25832 20924 25838 20936
rect 25869 20927 25927 20933
rect 25869 20924 25881 20927
rect 25832 20896 25881 20924
rect 25832 20884 25838 20896
rect 25869 20893 25881 20896
rect 25915 20893 25927 20927
rect 25869 20887 25927 20893
rect 26605 20927 26663 20933
rect 26605 20893 26617 20927
rect 26651 20924 26663 20927
rect 26712 20924 26740 21032
rect 27433 21029 27445 21032
rect 27479 21029 27491 21063
rect 27433 21023 27491 21029
rect 27985 20995 28043 21001
rect 27985 20961 27997 20995
rect 28031 20961 28043 20995
rect 28092 20992 28120 21100
rect 28626 21088 28632 21140
rect 28684 21128 28690 21140
rect 34977 21131 35035 21137
rect 34977 21128 34989 21131
rect 28684 21100 34989 21128
rect 28684 21088 28690 21100
rect 34977 21097 34989 21100
rect 35023 21097 35035 21131
rect 34977 21091 35035 21097
rect 38470 21088 38476 21140
rect 38528 21128 38534 21140
rect 42334 21128 42340 21140
rect 38528 21100 42340 21128
rect 38528 21088 38534 21100
rect 42334 21088 42340 21100
rect 42392 21088 42398 21140
rect 57974 21128 57980 21140
rect 51046 21100 57980 21128
rect 29178 21020 29184 21072
rect 29236 21060 29242 21072
rect 31573 21063 31631 21069
rect 31573 21060 31585 21063
rect 29236 21032 31585 21060
rect 29236 21020 29242 21032
rect 31573 21029 31585 21032
rect 31619 21029 31631 21063
rect 31573 21023 31631 21029
rect 31662 21020 31668 21072
rect 31720 21060 31726 21072
rect 51046 21060 51074 21100
rect 57974 21088 57980 21100
rect 58032 21088 58038 21140
rect 31720 21032 51074 21060
rect 31720 21020 31726 21032
rect 53374 21020 53380 21072
rect 53432 21020 53438 21072
rect 59262 21060 59268 21072
rect 53484 21032 59268 21060
rect 36357 20995 36415 21001
rect 28092 20964 36308 20992
rect 27985 20955 28043 20961
rect 26651 20896 26740 20924
rect 26651 20893 26663 20896
rect 26605 20887 26663 20893
rect 26786 20884 26792 20936
rect 26844 20924 26850 20936
rect 27798 20924 27804 20936
rect 26844 20896 27804 20924
rect 26844 20884 26850 20896
rect 27798 20884 27804 20896
rect 27856 20884 27862 20936
rect 28000 20924 28028 20955
rect 28626 20924 28632 20936
rect 28000 20896 28632 20924
rect 28626 20884 28632 20896
rect 28684 20884 28690 20936
rect 30650 20884 30656 20936
rect 30708 20884 30714 20936
rect 30742 20884 30748 20936
rect 30800 20884 30806 20936
rect 30926 20884 30932 20936
rect 30984 20884 30990 20936
rect 31386 20884 31392 20936
rect 31444 20884 31450 20936
rect 34790 20884 34796 20936
rect 34848 20884 34854 20936
rect 35437 20927 35495 20933
rect 35437 20893 35449 20927
rect 35483 20924 35495 20927
rect 35618 20924 35624 20936
rect 35483 20896 35624 20924
rect 35483 20893 35495 20896
rect 35437 20887 35495 20893
rect 35618 20884 35624 20896
rect 35676 20924 35682 20936
rect 36280 20924 36308 20964
rect 36357 20961 36369 20995
rect 36403 20992 36415 20995
rect 36538 20992 36544 21004
rect 36403 20964 36544 20992
rect 36403 20961 36415 20964
rect 36357 20955 36415 20961
rect 36538 20952 36544 20964
rect 36596 20952 36602 21004
rect 41874 20992 41880 21004
rect 36924 20964 41880 20992
rect 36924 20933 36952 20964
rect 41874 20952 41880 20964
rect 41932 20952 41938 21004
rect 42242 20952 42248 21004
rect 42300 20952 42306 21004
rect 53484 20992 53512 21032
rect 59262 21020 59268 21032
rect 59320 21020 59326 21072
rect 43272 20964 53512 20992
rect 36909 20927 36967 20933
rect 36909 20924 36921 20927
rect 35676 20896 36216 20924
rect 36280 20896 36921 20924
rect 35676 20884 35682 20896
rect 17954 20856 17960 20868
rect 16500 20828 17960 20856
rect 17954 20816 17960 20828
rect 18012 20816 18018 20868
rect 18506 20816 18512 20868
rect 18564 20856 18570 20868
rect 34808 20856 34836 20884
rect 18564 20828 21956 20856
rect 18564 20816 18570 20828
rect 11974 20748 11980 20800
rect 12032 20788 12038 20800
rect 12989 20791 13047 20797
rect 12989 20788 13001 20791
rect 12032 20760 13001 20788
rect 12032 20748 12038 20760
rect 12989 20757 13001 20760
rect 13035 20757 13047 20791
rect 12989 20751 13047 20757
rect 13998 20748 14004 20800
rect 14056 20788 14062 20800
rect 14461 20791 14519 20797
rect 14461 20788 14473 20791
rect 14056 20760 14473 20788
rect 14056 20748 14062 20760
rect 14461 20757 14473 20760
rect 14507 20757 14519 20791
rect 14461 20751 14519 20757
rect 15286 20748 15292 20800
rect 15344 20748 15350 20800
rect 16025 20791 16083 20797
rect 16025 20757 16037 20791
rect 16071 20788 16083 20791
rect 17126 20788 17132 20800
rect 16071 20760 17132 20788
rect 16071 20757 16083 20760
rect 16025 20751 16083 20757
rect 17126 20748 17132 20760
rect 17184 20748 17190 20800
rect 17494 20748 17500 20800
rect 17552 20748 17558 20800
rect 18322 20748 18328 20800
rect 18380 20788 18386 20800
rect 18966 20788 18972 20800
rect 18380 20760 18972 20788
rect 18380 20748 18386 20760
rect 18966 20748 18972 20760
rect 19024 20788 19030 20800
rect 21821 20791 21879 20797
rect 21821 20788 21833 20791
rect 19024 20760 21833 20788
rect 19024 20748 19030 20760
rect 21821 20757 21833 20760
rect 21867 20757 21879 20791
rect 21928 20788 21956 20828
rect 24780 20828 34836 20856
rect 24780 20788 24808 20828
rect 21928 20760 24808 20788
rect 21821 20751 21879 20757
rect 24946 20748 24952 20800
rect 25004 20748 25010 20800
rect 26786 20748 26792 20800
rect 26844 20748 26850 20800
rect 27157 20791 27215 20797
rect 27157 20757 27169 20791
rect 27203 20788 27215 20791
rect 27614 20788 27620 20800
rect 27203 20760 27620 20788
rect 27203 20757 27215 20760
rect 27157 20751 27215 20757
rect 27614 20748 27620 20760
rect 27672 20788 27678 20800
rect 27893 20791 27951 20797
rect 27893 20788 27905 20791
rect 27672 20760 27905 20788
rect 27672 20748 27678 20760
rect 27893 20757 27905 20760
rect 27939 20788 27951 20791
rect 31662 20788 31668 20800
rect 27939 20760 31668 20788
rect 27939 20757 27951 20760
rect 27893 20751 27951 20757
rect 31662 20748 31668 20760
rect 31720 20748 31726 20800
rect 35710 20748 35716 20800
rect 35768 20748 35774 20800
rect 35986 20748 35992 20800
rect 36044 20788 36050 20800
rect 36188 20797 36216 20896
rect 36909 20893 36921 20896
rect 36955 20893 36967 20927
rect 36909 20887 36967 20893
rect 38470 20884 38476 20936
rect 38528 20884 38534 20936
rect 38562 20884 38568 20936
rect 38620 20884 38626 20936
rect 41966 20884 41972 20936
rect 42024 20924 42030 20936
rect 42153 20927 42211 20933
rect 42153 20924 42165 20927
rect 42024 20896 42165 20924
rect 42024 20884 42030 20896
rect 42153 20893 42165 20896
rect 42199 20893 42211 20927
rect 42153 20887 42211 20893
rect 43272 20856 43300 20964
rect 53834 20952 53840 21004
rect 53892 20992 53898 21004
rect 53892 20964 54064 20992
rect 53892 20952 53898 20964
rect 45554 20884 45560 20936
rect 45612 20924 45618 20936
rect 47489 20927 47547 20933
rect 47489 20924 47501 20927
rect 45612 20896 47501 20924
rect 45612 20884 45618 20896
rect 47489 20893 47501 20896
rect 47535 20893 47547 20927
rect 47489 20887 47547 20893
rect 47854 20884 47860 20936
rect 47912 20884 47918 20936
rect 52825 20927 52883 20933
rect 52825 20924 52837 20927
rect 52656 20896 52837 20924
rect 37016 20828 43300 20856
rect 36081 20791 36139 20797
rect 36081 20788 36093 20791
rect 36044 20760 36093 20788
rect 36044 20748 36050 20760
rect 36081 20757 36093 20760
rect 36127 20757 36139 20791
rect 36081 20751 36139 20757
rect 36173 20791 36231 20797
rect 36173 20757 36185 20791
rect 36219 20788 36231 20791
rect 37016 20788 37044 20828
rect 43346 20816 43352 20868
rect 43404 20856 43410 20868
rect 43806 20856 43812 20868
rect 43404 20828 43812 20856
rect 43404 20816 43410 20828
rect 43806 20816 43812 20828
rect 43864 20816 43870 20868
rect 47670 20816 47676 20868
rect 47728 20816 47734 20868
rect 47765 20859 47823 20865
rect 47765 20825 47777 20859
rect 47811 20856 47823 20859
rect 48958 20856 48964 20868
rect 47811 20828 48964 20856
rect 47811 20825 47823 20828
rect 47765 20819 47823 20825
rect 48958 20816 48964 20828
rect 49016 20856 49022 20868
rect 49602 20856 49608 20868
rect 49016 20828 49608 20856
rect 49016 20816 49022 20828
rect 49602 20816 49608 20828
rect 49660 20816 49666 20868
rect 52656 20800 52684 20896
rect 52825 20893 52837 20896
rect 52871 20893 52883 20927
rect 52825 20887 52883 20893
rect 52914 20884 52920 20936
rect 52972 20924 52978 20936
rect 53193 20927 53251 20933
rect 53193 20924 53205 20927
rect 52972 20896 53205 20924
rect 52972 20884 52978 20896
rect 53193 20893 53205 20896
rect 53239 20893 53251 20927
rect 53193 20887 53251 20893
rect 53926 20884 53932 20936
rect 53984 20884 53990 20936
rect 54036 20933 54064 20964
rect 54021 20927 54079 20933
rect 54021 20893 54033 20927
rect 54067 20893 54079 20927
rect 54021 20887 54079 20893
rect 55674 20884 55680 20936
rect 55732 20924 55738 20936
rect 55861 20927 55919 20933
rect 55861 20924 55873 20927
rect 55732 20896 55873 20924
rect 55732 20884 55738 20896
rect 55861 20893 55873 20896
rect 55907 20893 55919 20927
rect 55861 20887 55919 20893
rect 56042 20884 56048 20936
rect 56100 20884 56106 20936
rect 57882 20884 57888 20936
rect 57940 20884 57946 20936
rect 53009 20859 53067 20865
rect 53009 20825 53021 20859
rect 53055 20825 53067 20859
rect 53009 20819 53067 20825
rect 53101 20859 53159 20865
rect 53101 20825 53113 20859
rect 53147 20856 53159 20859
rect 54478 20856 54484 20868
rect 53147 20828 54484 20856
rect 53147 20825 53159 20828
rect 53101 20819 53159 20825
rect 36219 20760 37044 20788
rect 36219 20757 36231 20760
rect 36173 20751 36231 20757
rect 37090 20748 37096 20800
rect 37148 20748 37154 20800
rect 38746 20748 38752 20800
rect 38804 20748 38810 20800
rect 41598 20748 41604 20800
rect 41656 20788 41662 20800
rect 41693 20791 41751 20797
rect 41693 20788 41705 20791
rect 41656 20760 41705 20788
rect 41656 20748 41662 20760
rect 41693 20757 41705 20760
rect 41739 20757 41751 20791
rect 41693 20751 41751 20757
rect 41874 20748 41880 20800
rect 41932 20788 41938 20800
rect 42061 20791 42119 20797
rect 42061 20788 42073 20791
rect 41932 20760 42073 20788
rect 41932 20748 41938 20760
rect 42061 20757 42073 20760
rect 42107 20788 42119 20791
rect 42702 20788 42708 20800
rect 42107 20760 42708 20788
rect 42107 20757 42119 20760
rect 42061 20751 42119 20757
rect 42702 20748 42708 20760
rect 42760 20748 42766 20800
rect 43622 20748 43628 20800
rect 43680 20748 43686 20800
rect 48041 20791 48099 20797
rect 48041 20757 48053 20791
rect 48087 20788 48099 20791
rect 48314 20788 48320 20800
rect 48087 20760 48320 20788
rect 48087 20757 48099 20760
rect 48041 20751 48099 20757
rect 48314 20748 48320 20760
rect 48372 20748 48378 20800
rect 52549 20791 52607 20797
rect 52549 20757 52561 20791
rect 52595 20788 52607 20791
rect 52638 20788 52644 20800
rect 52595 20760 52644 20788
rect 52595 20757 52607 20760
rect 52549 20751 52607 20757
rect 52638 20748 52644 20760
rect 52696 20748 52702 20800
rect 53024 20788 53052 20819
rect 54478 20816 54484 20828
rect 54536 20816 54542 20868
rect 58161 20859 58219 20865
rect 58161 20825 58173 20859
rect 58207 20856 58219 20859
rect 58986 20856 58992 20868
rect 58207 20828 58992 20856
rect 58207 20825 58219 20828
rect 58161 20819 58219 20825
rect 58986 20816 58992 20828
rect 59044 20816 59050 20868
rect 53834 20788 53840 20800
rect 53024 20760 53840 20788
rect 53834 20748 53840 20760
rect 53892 20748 53898 20800
rect 54202 20748 54208 20800
rect 54260 20748 54266 20800
rect 56229 20791 56287 20797
rect 56229 20757 56241 20791
rect 56275 20788 56287 20791
rect 56962 20788 56968 20800
rect 56275 20760 56968 20788
rect 56275 20757 56287 20760
rect 56229 20751 56287 20757
rect 56962 20748 56968 20760
rect 57020 20748 57026 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 16206 20544 16212 20596
rect 16264 20544 16270 20596
rect 18230 20544 18236 20596
rect 18288 20584 18294 20596
rect 19169 20587 19227 20593
rect 19169 20584 19181 20587
rect 18288 20556 19181 20584
rect 18288 20544 18294 20556
rect 19169 20553 19181 20556
rect 19215 20553 19227 20587
rect 19169 20547 19227 20553
rect 19337 20587 19395 20593
rect 19337 20553 19349 20587
rect 19383 20584 19395 20587
rect 19426 20584 19432 20596
rect 19383 20556 19432 20584
rect 19383 20553 19395 20556
rect 19337 20547 19395 20553
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 19812 20556 22094 20584
rect 11514 20476 11520 20528
rect 11572 20516 11578 20528
rect 15194 20516 15200 20528
rect 11572 20488 15200 20516
rect 11572 20476 11578 20488
rect 15194 20476 15200 20488
rect 15252 20476 15258 20528
rect 16942 20516 16948 20528
rect 16040 20488 16948 20516
rect 1581 20451 1639 20457
rect 1581 20417 1593 20451
rect 1627 20448 1639 20451
rect 3510 20448 3516 20460
rect 1627 20420 3516 20448
rect 1627 20417 1639 20420
rect 1581 20411 1639 20417
rect 3510 20408 3516 20420
rect 3568 20408 3574 20460
rect 8021 20451 8079 20457
rect 8021 20417 8033 20451
rect 8067 20448 8079 20451
rect 9306 20448 9312 20460
rect 8067 20420 9312 20448
rect 8067 20417 8079 20420
rect 8021 20411 8079 20417
rect 9306 20408 9312 20420
rect 9364 20408 9370 20460
rect 10226 20408 10232 20460
rect 10284 20408 10290 20460
rect 11977 20451 12035 20457
rect 11977 20417 11989 20451
rect 12023 20448 12035 20451
rect 12023 20420 12434 20448
rect 12023 20417 12035 20420
rect 11977 20411 12035 20417
rect 934 20340 940 20392
rect 992 20380 998 20392
rect 1765 20383 1823 20389
rect 1765 20380 1777 20383
rect 992 20352 1777 20380
rect 992 20340 998 20352
rect 1765 20349 1777 20352
rect 1811 20349 1823 20383
rect 12406 20380 12434 20420
rect 13170 20408 13176 20460
rect 13228 20408 13234 20460
rect 13262 20408 13268 20460
rect 13320 20408 13326 20460
rect 13998 20408 14004 20460
rect 14056 20408 14062 20460
rect 15286 20408 15292 20460
rect 15344 20408 15350 20460
rect 16040 20457 16068 20488
rect 16942 20476 16948 20488
rect 17000 20476 17006 20528
rect 18506 20476 18512 20528
rect 18564 20476 18570 20528
rect 18966 20476 18972 20528
rect 19024 20476 19030 20528
rect 19812 20525 19840 20556
rect 19797 20519 19855 20525
rect 19797 20485 19809 20519
rect 19843 20485 19855 20519
rect 19797 20479 19855 20485
rect 20013 20519 20071 20525
rect 20013 20485 20025 20519
rect 20059 20516 20071 20519
rect 20162 20516 20168 20528
rect 20059 20488 20168 20516
rect 20059 20485 20071 20488
rect 20013 20479 20071 20485
rect 16025 20451 16083 20457
rect 16025 20417 16037 20451
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 16850 20408 16856 20460
rect 16908 20408 16914 20460
rect 17126 20408 17132 20460
rect 17184 20408 17190 20460
rect 19150 20408 19156 20460
rect 19208 20448 19214 20460
rect 19812 20448 19840 20479
rect 20162 20476 20168 20488
rect 20220 20476 20226 20528
rect 22066 20516 22094 20556
rect 22462 20544 22468 20596
rect 22520 20544 22526 20596
rect 25590 20544 25596 20596
rect 25648 20544 25654 20596
rect 27798 20544 27804 20596
rect 27856 20584 27862 20596
rect 28442 20584 28448 20596
rect 27856 20556 28448 20584
rect 27856 20544 27862 20556
rect 28442 20544 28448 20556
rect 28500 20584 28506 20596
rect 28537 20587 28595 20593
rect 28537 20584 28549 20587
rect 28500 20556 28549 20584
rect 28500 20544 28506 20556
rect 28537 20553 28549 20556
rect 28583 20553 28595 20587
rect 28537 20547 28595 20553
rect 28902 20544 28908 20596
rect 28960 20584 28966 20596
rect 30101 20587 30159 20593
rect 30101 20584 30113 20587
rect 28960 20556 30113 20584
rect 28960 20544 28966 20556
rect 30101 20553 30113 20556
rect 30147 20553 30159 20587
rect 30101 20547 30159 20553
rect 30653 20587 30711 20593
rect 30653 20553 30665 20587
rect 30699 20584 30711 20587
rect 30742 20584 30748 20596
rect 30699 20556 30748 20584
rect 30699 20553 30711 20556
rect 30653 20547 30711 20553
rect 30742 20544 30748 20556
rect 30800 20544 30806 20596
rect 31018 20544 31024 20596
rect 31076 20544 31082 20596
rect 37090 20584 37096 20596
rect 31726 20556 37096 20584
rect 24020 20519 24078 20525
rect 22066 20488 23888 20516
rect 23860 20460 23888 20488
rect 24020 20485 24032 20519
rect 24066 20516 24078 20519
rect 24946 20516 24952 20528
rect 24066 20488 24952 20516
rect 24066 20485 24078 20488
rect 24020 20479 24078 20485
rect 24946 20476 24952 20488
rect 25004 20476 25010 20528
rect 25130 20476 25136 20528
rect 25188 20516 25194 20528
rect 25961 20519 26019 20525
rect 25961 20516 25973 20519
rect 25188 20488 25973 20516
rect 25188 20476 25194 20488
rect 25961 20485 25973 20488
rect 26007 20485 26019 20519
rect 25961 20479 26019 20485
rect 26786 20476 26792 20528
rect 26844 20516 26850 20528
rect 27402 20519 27460 20525
rect 27402 20516 27414 20519
rect 26844 20488 27414 20516
rect 26844 20476 26850 20488
rect 27402 20485 27414 20488
rect 27448 20485 27460 20519
rect 31726 20516 31754 20556
rect 37090 20544 37096 20556
rect 37148 20544 37154 20596
rect 37274 20544 37280 20596
rect 37332 20584 37338 20596
rect 37332 20556 39436 20584
rect 37332 20544 37338 20556
rect 27402 20479 27460 20485
rect 29196 20488 31754 20516
rect 34793 20519 34851 20525
rect 19208 20420 19840 20448
rect 21177 20451 21235 20457
rect 19208 20408 19214 20420
rect 21177 20417 21189 20451
rect 21223 20448 21235 20451
rect 21223 20420 22048 20448
rect 21223 20417 21235 20420
rect 21177 20411 21235 20417
rect 12805 20383 12863 20389
rect 12805 20380 12817 20383
rect 12406 20352 12817 20380
rect 1765 20343 1823 20349
rect 12805 20349 12817 20352
rect 12851 20349 12863 20383
rect 12805 20343 12863 20349
rect 12894 20340 12900 20392
rect 12952 20380 12958 20392
rect 12989 20383 13047 20389
rect 12989 20380 13001 20383
rect 12952 20352 13001 20380
rect 12952 20340 12958 20352
rect 12989 20349 13001 20352
rect 13035 20349 13047 20383
rect 12989 20343 13047 20349
rect 13078 20340 13084 20392
rect 13136 20340 13142 20392
rect 13722 20340 13728 20392
rect 13780 20380 13786 20392
rect 20898 20380 20904 20392
rect 13780 20352 20904 20380
rect 13780 20340 13786 20352
rect 20898 20340 20904 20352
rect 20956 20340 20962 20392
rect 20990 20340 20996 20392
rect 21048 20340 21054 20392
rect 11698 20272 11704 20324
rect 11756 20312 11762 20324
rect 11756 20284 16896 20312
rect 11756 20272 11762 20284
rect 8110 20204 8116 20256
rect 8168 20244 8174 20256
rect 8205 20247 8263 20253
rect 8205 20244 8217 20247
rect 8168 20216 8217 20244
rect 8168 20204 8174 20216
rect 8205 20213 8217 20216
rect 8251 20213 8263 20247
rect 8205 20207 8263 20213
rect 10318 20204 10324 20256
rect 10376 20244 10382 20256
rect 10413 20247 10471 20253
rect 10413 20244 10425 20247
rect 10376 20216 10425 20244
rect 10376 20204 10382 20216
rect 10413 20213 10425 20216
rect 10459 20213 10471 20247
rect 10413 20207 10471 20213
rect 10962 20204 10968 20256
rect 11020 20244 11026 20256
rect 12161 20247 12219 20253
rect 12161 20244 12173 20247
rect 11020 20216 12173 20244
rect 11020 20204 11026 20216
rect 12161 20213 12173 20216
rect 12207 20213 12219 20247
rect 12161 20207 12219 20213
rect 14182 20204 14188 20256
rect 14240 20204 14246 20256
rect 15470 20204 15476 20256
rect 15528 20204 15534 20256
rect 16868 20244 16896 20284
rect 18874 20272 18880 20324
rect 18932 20312 18938 20324
rect 20530 20312 20536 20324
rect 18932 20284 20536 20312
rect 18932 20272 18938 20284
rect 18782 20244 18788 20256
rect 16868 20216 18788 20244
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 19153 20247 19211 20253
rect 19153 20213 19165 20247
rect 19199 20244 19211 20247
rect 19242 20244 19248 20256
rect 19199 20216 19248 20244
rect 19199 20213 19211 20216
rect 19153 20207 19211 20213
rect 19242 20204 19248 20216
rect 19300 20204 19306 20256
rect 19996 20253 20024 20284
rect 20530 20272 20536 20284
rect 20588 20272 20594 20324
rect 20916 20312 20944 20340
rect 21726 20312 21732 20324
rect 20916 20284 21732 20312
rect 21726 20272 21732 20284
rect 21784 20272 21790 20324
rect 22020 20321 22048 20420
rect 22094 20408 22100 20460
rect 22152 20448 22158 20460
rect 22373 20451 22431 20457
rect 22373 20448 22385 20451
rect 22152 20420 22385 20448
rect 22152 20408 22158 20420
rect 22373 20417 22385 20420
rect 22419 20417 22431 20451
rect 22373 20411 22431 20417
rect 23842 20408 23848 20460
rect 23900 20448 23906 20460
rect 26053 20451 26111 20457
rect 23900 20420 25268 20448
rect 23900 20408 23906 20420
rect 22649 20383 22707 20389
rect 22649 20349 22661 20383
rect 22695 20380 22707 20383
rect 22695 20352 23336 20380
rect 22695 20349 22707 20352
rect 22649 20343 22707 20349
rect 22005 20315 22063 20321
rect 22005 20281 22017 20315
rect 22051 20281 22063 20315
rect 22005 20275 22063 20281
rect 19981 20247 20039 20253
rect 19981 20213 19993 20247
rect 20027 20213 20039 20247
rect 19981 20207 20039 20213
rect 20165 20247 20223 20253
rect 20165 20213 20177 20247
rect 20211 20244 20223 20247
rect 20346 20244 20352 20256
rect 20211 20216 20352 20244
rect 20211 20213 20223 20216
rect 20165 20207 20223 20213
rect 20346 20204 20352 20216
rect 20404 20204 20410 20256
rect 21358 20204 21364 20256
rect 21416 20204 21422 20256
rect 22830 20204 22836 20256
rect 22888 20244 22894 20256
rect 23198 20244 23204 20256
rect 22888 20216 23204 20244
rect 22888 20204 22894 20216
rect 23198 20204 23204 20216
rect 23256 20204 23262 20256
rect 23308 20244 23336 20352
rect 23382 20340 23388 20392
rect 23440 20380 23446 20392
rect 23753 20383 23811 20389
rect 23753 20380 23765 20383
rect 23440 20352 23765 20380
rect 23440 20340 23446 20352
rect 23753 20349 23765 20352
rect 23799 20349 23811 20383
rect 23753 20343 23811 20349
rect 24854 20244 24860 20256
rect 23308 20216 24860 20244
rect 24854 20204 24860 20216
rect 24912 20204 24918 20256
rect 25130 20204 25136 20256
rect 25188 20204 25194 20256
rect 25240 20244 25268 20420
rect 26053 20417 26065 20451
rect 26099 20448 26111 20451
rect 28994 20448 29000 20460
rect 26099 20420 29000 20448
rect 26099 20417 26111 20420
rect 26053 20411 26111 20417
rect 28994 20408 29000 20420
rect 29052 20408 29058 20460
rect 29196 20457 29224 20488
rect 34793 20485 34805 20519
rect 34839 20516 34851 20519
rect 35498 20519 35556 20525
rect 35498 20516 35510 20519
rect 34839 20488 35510 20516
rect 34839 20485 34851 20488
rect 34793 20479 34851 20485
rect 35498 20485 35510 20488
rect 35544 20485 35556 20519
rect 35498 20479 35556 20485
rect 35710 20476 35716 20528
rect 35768 20476 35774 20528
rect 36078 20476 36084 20528
rect 36136 20516 36142 20528
rect 37829 20519 37887 20525
rect 37829 20516 37841 20519
rect 36136 20488 37841 20516
rect 36136 20476 36142 20488
rect 37829 20485 37841 20488
rect 37875 20485 37887 20519
rect 39408 20516 39436 20556
rect 40034 20544 40040 20596
rect 40092 20584 40098 20596
rect 40678 20584 40684 20596
rect 40092 20556 40684 20584
rect 40092 20544 40098 20556
rect 40678 20544 40684 20556
rect 40736 20544 40742 20596
rect 44450 20584 44456 20596
rect 43732 20556 44456 20584
rect 42889 20519 42947 20525
rect 42889 20516 42901 20519
rect 39408 20488 42901 20516
rect 37829 20479 37887 20485
rect 42889 20485 42901 20488
rect 42935 20485 42947 20519
rect 42889 20479 42947 20485
rect 43119 20519 43177 20525
rect 43119 20485 43131 20519
rect 43165 20516 43177 20519
rect 43732 20516 43760 20556
rect 44218 20525 44246 20556
rect 44450 20544 44456 20556
rect 44508 20544 44514 20596
rect 49602 20544 49608 20596
rect 49660 20544 49666 20596
rect 56318 20544 56324 20596
rect 56376 20544 56382 20596
rect 43165 20488 43760 20516
rect 44203 20519 44261 20525
rect 43165 20485 43177 20488
rect 43119 20479 43177 20485
rect 44203 20485 44215 20519
rect 44249 20485 44261 20519
rect 44726 20516 44732 20528
rect 44203 20479 44261 20485
rect 44376 20488 44732 20516
rect 29181 20451 29239 20457
rect 29181 20417 29193 20451
rect 29227 20417 29239 20451
rect 29181 20411 29239 20417
rect 29917 20451 29975 20457
rect 29917 20417 29929 20451
rect 29963 20417 29975 20451
rect 29917 20411 29975 20417
rect 25498 20340 25504 20392
rect 25556 20380 25562 20392
rect 26145 20383 26203 20389
rect 26145 20380 26157 20383
rect 25556 20352 26157 20380
rect 25556 20340 25562 20352
rect 26145 20349 26157 20352
rect 26191 20349 26203 20383
rect 26145 20343 26203 20349
rect 26510 20340 26516 20392
rect 26568 20380 26574 20392
rect 27157 20383 27215 20389
rect 27157 20380 27169 20383
rect 26568 20352 27169 20380
rect 26568 20340 26574 20352
rect 27157 20349 27169 20352
rect 27203 20349 27215 20383
rect 27157 20343 27215 20349
rect 29086 20340 29092 20392
rect 29144 20380 29150 20392
rect 29932 20380 29960 20411
rect 30190 20408 30196 20460
rect 30248 20448 30254 20460
rect 30650 20448 30656 20460
rect 30248 20420 30656 20448
rect 30248 20408 30254 20420
rect 30650 20408 30656 20420
rect 30708 20448 30714 20460
rect 33229 20451 33287 20457
rect 33229 20448 33241 20451
rect 30708 20420 33241 20448
rect 30708 20408 30714 20420
rect 33229 20417 33241 20420
rect 33275 20417 33287 20451
rect 33229 20411 33287 20417
rect 33410 20408 33416 20460
rect 33468 20408 33474 20460
rect 33594 20408 33600 20460
rect 33652 20408 33658 20460
rect 34609 20451 34667 20457
rect 34609 20417 34621 20451
rect 34655 20448 34667 20451
rect 35728 20448 35756 20476
rect 34655 20420 35756 20448
rect 34655 20417 34667 20420
rect 34609 20411 34667 20417
rect 35894 20408 35900 20460
rect 35952 20448 35958 20460
rect 37645 20451 37703 20457
rect 37645 20448 37657 20451
rect 35952 20420 37657 20448
rect 35952 20408 35958 20420
rect 37645 20417 37657 20420
rect 37691 20417 37703 20451
rect 37645 20411 37703 20417
rect 38746 20408 38752 20460
rect 38804 20408 38810 20460
rect 41598 20408 41604 20460
rect 41656 20408 41662 20460
rect 42794 20408 42800 20460
rect 42852 20408 42858 20460
rect 42981 20451 43039 20457
rect 42981 20417 42993 20451
rect 43027 20417 43039 20451
rect 42981 20411 43039 20417
rect 30742 20380 30748 20392
rect 29144 20352 30748 20380
rect 29144 20340 29150 20352
rect 30742 20340 30748 20352
rect 30800 20340 30806 20392
rect 31110 20340 31116 20392
rect 31168 20340 31174 20392
rect 31205 20383 31263 20389
rect 31205 20349 31217 20383
rect 31251 20380 31263 20383
rect 31478 20380 31484 20392
rect 31251 20352 31484 20380
rect 31251 20349 31263 20352
rect 31205 20343 31263 20349
rect 31478 20340 31484 20352
rect 31536 20340 31542 20392
rect 33318 20340 33324 20392
rect 33376 20380 33382 20392
rect 34425 20383 34483 20389
rect 34425 20380 34437 20383
rect 33376 20352 34437 20380
rect 33376 20340 33382 20352
rect 34425 20349 34437 20352
rect 34471 20349 34483 20383
rect 34425 20343 34483 20349
rect 35253 20383 35311 20389
rect 35253 20349 35265 20383
rect 35299 20349 35311 20383
rect 35253 20343 35311 20349
rect 37461 20383 37519 20389
rect 37461 20349 37473 20383
rect 37507 20380 37519 20383
rect 38378 20380 38384 20392
rect 37507 20352 38384 20380
rect 37507 20349 37519 20352
rect 37461 20343 37519 20349
rect 28092 20284 28672 20312
rect 28092 20244 28120 20284
rect 25240 20216 28120 20244
rect 28644 20244 28672 20284
rect 32858 20272 32864 20324
rect 32916 20312 32922 20324
rect 35268 20312 35296 20343
rect 38378 20340 38384 20352
rect 38436 20340 38442 20392
rect 38473 20383 38531 20389
rect 38473 20349 38485 20383
rect 38519 20349 38531 20383
rect 38473 20343 38531 20349
rect 41417 20383 41475 20389
rect 41417 20349 41429 20383
rect 41463 20380 41475 20383
rect 41690 20380 41696 20392
rect 41463 20352 41696 20380
rect 41463 20349 41475 20352
rect 41417 20343 41475 20349
rect 32916 20284 35296 20312
rect 32916 20272 32922 20284
rect 37182 20272 37188 20324
rect 37240 20312 37246 20324
rect 38488 20312 38516 20343
rect 41690 20340 41696 20352
rect 41748 20340 41754 20392
rect 37240 20284 38516 20312
rect 37240 20272 37246 20284
rect 39666 20272 39672 20324
rect 39724 20312 39730 20324
rect 42996 20312 43024 20411
rect 43714 20408 43720 20460
rect 43772 20408 43778 20460
rect 43898 20408 43904 20460
rect 43956 20408 43962 20460
rect 43990 20408 43996 20460
rect 44048 20408 44054 20460
rect 44376 20457 44404 20488
rect 44726 20476 44732 20488
rect 44784 20516 44790 20528
rect 57698 20516 57704 20528
rect 44784 20488 57704 20516
rect 44784 20476 44790 20488
rect 57698 20476 57704 20488
rect 57756 20476 57762 20528
rect 44085 20451 44143 20457
rect 44085 20417 44097 20451
rect 44131 20417 44143 20451
rect 44085 20411 44143 20417
rect 44361 20451 44419 20457
rect 44361 20417 44373 20451
rect 44407 20417 44419 20451
rect 44361 20411 44419 20417
rect 46017 20451 46075 20457
rect 46017 20417 46029 20451
rect 46063 20448 46075 20451
rect 46750 20448 46756 20460
rect 46063 20420 46756 20448
rect 46063 20417 46075 20420
rect 46017 20411 46075 20417
rect 43257 20383 43315 20389
rect 43257 20349 43269 20383
rect 43303 20380 43315 20383
rect 43346 20380 43352 20392
rect 43303 20352 43352 20380
rect 43303 20349 43315 20352
rect 43257 20343 43315 20349
rect 43346 20340 43352 20352
rect 43404 20340 43410 20392
rect 44100 20380 44128 20411
rect 46750 20408 46756 20420
rect 46808 20408 46814 20460
rect 48498 20457 48504 20460
rect 48492 20411 48504 20457
rect 48498 20408 48504 20411
rect 48556 20408 48562 20460
rect 50154 20408 50160 20460
rect 50212 20448 50218 20460
rect 50433 20451 50491 20457
rect 50433 20448 50445 20451
rect 50212 20420 50445 20448
rect 50212 20408 50218 20420
rect 50433 20417 50445 20420
rect 50479 20417 50491 20451
rect 50433 20411 50491 20417
rect 51626 20408 51632 20460
rect 51684 20408 51690 20460
rect 53101 20451 53159 20457
rect 53101 20417 53113 20451
rect 53147 20417 53159 20451
rect 53101 20411 53159 20417
rect 53368 20451 53426 20457
rect 53368 20417 53380 20451
rect 53414 20448 53426 20451
rect 54202 20448 54208 20460
rect 53414 20420 54208 20448
rect 53414 20417 53426 20420
rect 53368 20411 53426 20417
rect 46934 20380 46940 20392
rect 44100 20352 46940 20380
rect 44100 20312 44128 20352
rect 46934 20340 46940 20352
rect 46992 20380 46998 20392
rect 47670 20380 47676 20392
rect 46992 20352 47676 20380
rect 46992 20340 46998 20352
rect 47670 20340 47676 20352
rect 47728 20340 47734 20392
rect 48222 20340 48228 20392
rect 48280 20340 48286 20392
rect 49234 20340 49240 20392
rect 49292 20380 49298 20392
rect 50249 20383 50307 20389
rect 50249 20380 50261 20383
rect 49292 20352 50261 20380
rect 49292 20340 49298 20352
rect 50249 20349 50261 20352
rect 50295 20380 50307 20383
rect 51442 20380 51448 20392
rect 50295 20352 51448 20380
rect 50295 20349 50307 20352
rect 50249 20343 50307 20349
rect 51442 20340 51448 20352
rect 51500 20340 51506 20392
rect 39724 20284 42748 20312
rect 42996 20284 44128 20312
rect 39724 20272 39730 20284
rect 29365 20247 29423 20253
rect 29365 20244 29377 20247
rect 28644 20216 29377 20244
rect 29365 20213 29377 20216
rect 29411 20213 29423 20247
rect 29365 20207 29423 20213
rect 30742 20204 30748 20256
rect 30800 20244 30806 20256
rect 35986 20244 35992 20256
rect 30800 20216 35992 20244
rect 30800 20204 30806 20216
rect 35986 20204 35992 20216
rect 36044 20244 36050 20256
rect 36633 20247 36691 20253
rect 36633 20244 36645 20247
rect 36044 20216 36645 20244
rect 36044 20204 36050 20216
rect 36633 20213 36645 20216
rect 36679 20244 36691 20247
rect 37090 20244 37096 20256
rect 36679 20216 37096 20244
rect 36679 20213 36691 20216
rect 36633 20207 36691 20213
rect 37090 20204 37096 20216
rect 37148 20204 37154 20256
rect 41782 20204 41788 20256
rect 41840 20204 41846 20256
rect 41874 20204 41880 20256
rect 41932 20244 41938 20256
rect 42613 20247 42671 20253
rect 42613 20244 42625 20247
rect 41932 20216 42625 20244
rect 41932 20204 41938 20216
rect 42613 20213 42625 20216
rect 42659 20213 42671 20247
rect 42720 20244 42748 20284
rect 52362 20272 52368 20324
rect 52420 20312 52426 20324
rect 53116 20312 53144 20411
rect 54202 20408 54208 20420
rect 54260 20408 54266 20460
rect 55030 20408 55036 20460
rect 55088 20448 55094 20460
rect 55197 20451 55255 20457
rect 55197 20448 55209 20451
rect 55088 20420 55209 20448
rect 55088 20408 55094 20420
rect 55197 20417 55209 20420
rect 55243 20417 55255 20451
rect 55197 20411 55255 20417
rect 54941 20383 54999 20389
rect 54941 20349 54953 20383
rect 54987 20349 54999 20383
rect 54941 20343 54999 20349
rect 52420 20284 53144 20312
rect 52420 20272 52426 20284
rect 43990 20244 43996 20256
rect 42720 20216 43996 20244
rect 42613 20207 42671 20213
rect 43990 20204 43996 20216
rect 44048 20204 44054 20256
rect 45370 20204 45376 20256
rect 45428 20244 45434 20256
rect 46293 20247 46351 20253
rect 46293 20244 46305 20247
rect 45428 20216 46305 20244
rect 45428 20204 45434 20216
rect 46293 20213 46305 20216
rect 46339 20244 46351 20247
rect 48406 20244 48412 20256
rect 46339 20216 48412 20244
rect 46339 20213 46351 20216
rect 46293 20207 46351 20213
rect 48406 20204 48412 20216
rect 48464 20204 48470 20256
rect 50522 20204 50528 20256
rect 50580 20244 50586 20256
rect 50617 20247 50675 20253
rect 50617 20244 50629 20247
rect 50580 20216 50629 20244
rect 50580 20204 50586 20216
rect 50617 20213 50629 20216
rect 50663 20213 50675 20247
rect 50617 20207 50675 20213
rect 51813 20247 51871 20253
rect 51813 20213 51825 20247
rect 51859 20244 51871 20247
rect 52454 20244 52460 20256
rect 51859 20216 52460 20244
rect 51859 20213 51871 20216
rect 51813 20207 51871 20213
rect 52454 20204 52460 20216
rect 52512 20204 52518 20256
rect 53116 20244 53144 20284
rect 54478 20272 54484 20324
rect 54536 20272 54542 20324
rect 54956 20244 54984 20343
rect 55858 20244 55864 20256
rect 53116 20216 55864 20244
rect 55858 20204 55864 20216
rect 55916 20204 55922 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 2746 20012 8248 20040
rect 1581 19839 1639 19845
rect 1581 19805 1593 19839
rect 1627 19836 1639 19839
rect 2746 19836 2774 20012
rect 8110 19932 8116 19984
rect 8168 19932 8174 19984
rect 8220 19972 8248 20012
rect 9306 20000 9312 20052
rect 9364 20000 9370 20052
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 17954 20040 17960 20052
rect 10192 20012 17960 20040
rect 10192 20000 10198 20012
rect 17954 20000 17960 20012
rect 18012 20000 18018 20052
rect 18325 20043 18383 20049
rect 18325 20009 18337 20043
rect 18371 20040 18383 20043
rect 20070 20040 20076 20052
rect 18371 20012 20076 20040
rect 18371 20009 18383 20012
rect 18325 20003 18383 20009
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 20162 20000 20168 20052
rect 20220 20000 20226 20052
rect 23382 20040 23388 20052
rect 20732 20012 23388 20040
rect 8220 19944 11744 19972
rect 8205 19907 8263 19913
rect 8205 19904 8217 19907
rect 7024 19876 8217 19904
rect 7024 19845 7052 19876
rect 8205 19873 8217 19876
rect 8251 19873 8263 19907
rect 11238 19904 11244 19916
rect 8205 19867 8263 19873
rect 8312 19876 11244 19904
rect 1627 19808 2774 19836
rect 7009 19839 7067 19845
rect 1627 19805 1639 19808
rect 1581 19799 1639 19805
rect 7009 19805 7021 19839
rect 7055 19805 7067 19839
rect 7009 19799 7067 19805
rect 7558 19796 7564 19848
rect 7616 19836 7622 19848
rect 8312 19836 8340 19876
rect 11238 19864 11244 19876
rect 11296 19864 11302 19916
rect 11606 19864 11612 19916
rect 11664 19864 11670 19916
rect 11716 19904 11744 19944
rect 11882 19932 11888 19984
rect 11940 19932 11946 19984
rect 13722 19932 13728 19984
rect 13780 19932 13786 19984
rect 16390 19932 16396 19984
rect 16448 19932 16454 19984
rect 19613 19975 19671 19981
rect 19613 19941 19625 19975
rect 19659 19972 19671 19975
rect 20254 19972 20260 19984
rect 19659 19944 20260 19972
rect 19659 19941 19671 19944
rect 19613 19935 19671 19941
rect 20254 19932 20260 19944
rect 20312 19932 20318 19984
rect 11716 19876 12480 19904
rect 7616 19808 8340 19836
rect 7616 19796 7622 19808
rect 8386 19796 8392 19848
rect 8444 19836 8450 19848
rect 9125 19839 9183 19845
rect 9125 19836 9137 19839
rect 8444 19808 9137 19836
rect 8444 19796 8450 19808
rect 9125 19805 9137 19808
rect 9171 19805 9183 19839
rect 9125 19799 9183 19805
rect 9858 19796 9864 19848
rect 9916 19796 9922 19848
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19836 10655 19839
rect 11146 19836 11152 19848
rect 10643 19808 11152 19836
rect 10643 19805 10655 19808
rect 10597 19799 10655 19805
rect 11146 19796 11152 19808
rect 11204 19796 11210 19848
rect 11514 19796 11520 19848
rect 11572 19796 11578 19848
rect 12342 19796 12348 19848
rect 12400 19796 12406 19848
rect 12452 19836 12480 19876
rect 16850 19864 16856 19916
rect 16908 19904 16914 19916
rect 16945 19907 17003 19913
rect 16945 19904 16957 19907
rect 16908 19876 16957 19904
rect 16908 19864 16914 19876
rect 16945 19873 16957 19876
rect 16991 19873 17003 19907
rect 16945 19867 17003 19873
rect 20070 19864 20076 19916
rect 20128 19904 20134 19916
rect 20732 19913 20760 20012
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 24946 20040 24952 20052
rect 24504 20012 24952 20040
rect 21726 19932 21732 19984
rect 21784 19972 21790 19984
rect 24504 19972 24532 20012
rect 24946 20000 24952 20012
rect 25004 20040 25010 20052
rect 25130 20040 25136 20052
rect 25004 20012 25136 20040
rect 25004 20000 25010 20012
rect 25130 20000 25136 20012
rect 25188 20000 25194 20052
rect 26142 20000 26148 20052
rect 26200 20040 26206 20052
rect 31018 20040 31024 20052
rect 26200 20012 31024 20040
rect 26200 20000 26206 20012
rect 31018 20000 31024 20012
rect 31076 20040 31082 20052
rect 32033 20043 32091 20049
rect 32033 20040 32045 20043
rect 31076 20012 32045 20040
rect 31076 20000 31082 20012
rect 32033 20009 32045 20012
rect 32079 20009 32091 20043
rect 32033 20003 32091 20009
rect 40865 20043 40923 20049
rect 40865 20009 40877 20043
rect 40911 20040 40923 20043
rect 42794 20040 42800 20052
rect 40911 20012 42800 20040
rect 40911 20009 40923 20012
rect 40865 20003 40923 20009
rect 42794 20000 42800 20012
rect 42852 20000 42858 20052
rect 43438 20040 43444 20052
rect 42904 20012 43444 20040
rect 21784 19944 24532 19972
rect 24581 19975 24639 19981
rect 21784 19932 21790 19944
rect 24581 19941 24593 19975
rect 24627 19972 24639 19975
rect 24627 19944 26004 19972
rect 24627 19941 24639 19944
rect 24581 19935 24639 19941
rect 20717 19907 20775 19913
rect 20717 19904 20729 19907
rect 20128 19876 20729 19904
rect 20128 19864 20134 19876
rect 20717 19873 20729 19876
rect 20763 19873 20775 19907
rect 20717 19867 20775 19873
rect 23198 19864 23204 19916
rect 23256 19904 23262 19916
rect 23256 19876 23428 19904
rect 23256 19864 23262 19876
rect 13538 19836 13544 19848
rect 12452 19808 13544 19836
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 14277 19839 14335 19845
rect 14277 19805 14289 19839
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 934 19728 940 19780
rect 992 19768 998 19780
rect 1857 19771 1915 19777
rect 1857 19768 1869 19771
rect 992 19740 1869 19768
rect 992 19728 998 19740
rect 1857 19737 1869 19740
rect 1903 19737 1915 19771
rect 1857 19731 1915 19737
rect 6914 19728 6920 19780
rect 6972 19768 6978 19780
rect 7745 19771 7803 19777
rect 7745 19768 7757 19771
rect 6972 19740 7757 19768
rect 6972 19728 6978 19740
rect 7745 19737 7757 19740
rect 7791 19737 7803 19771
rect 12590 19771 12648 19777
rect 12590 19768 12602 19771
rect 7745 19731 7803 19737
rect 10796 19740 12602 19768
rect 7098 19660 7104 19712
rect 7156 19700 7162 19712
rect 7193 19703 7251 19709
rect 7193 19700 7205 19703
rect 7156 19672 7205 19700
rect 7156 19660 7162 19672
rect 7193 19669 7205 19672
rect 7239 19669 7251 19703
rect 7193 19663 7251 19669
rect 10042 19660 10048 19712
rect 10100 19660 10106 19712
rect 10796 19709 10824 19740
rect 12590 19737 12602 19740
rect 12636 19737 12648 19771
rect 14292 19768 14320 19799
rect 14366 19796 14372 19848
rect 14424 19836 14430 19848
rect 15013 19839 15071 19845
rect 15013 19836 15025 19839
rect 14424 19808 15025 19836
rect 14424 19796 14430 19808
rect 15013 19805 15025 19808
rect 15059 19836 15071 19839
rect 16868 19836 16896 19864
rect 15059 19808 16896 19836
rect 17212 19839 17270 19845
rect 15059 19805 15071 19808
rect 15013 19799 15071 19805
rect 17212 19805 17224 19839
rect 17258 19836 17270 19839
rect 17494 19836 17500 19848
rect 17258 19808 17500 19836
rect 17258 19805 17270 19808
rect 17212 19799 17270 19805
rect 17494 19796 17500 19808
rect 17552 19796 17558 19848
rect 19981 19839 20039 19845
rect 19981 19805 19993 19839
rect 20027 19836 20039 19839
rect 20806 19836 20812 19848
rect 20027 19808 20812 19836
rect 20027 19805 20039 19808
rect 19981 19799 20039 19805
rect 20806 19796 20812 19808
rect 20864 19796 20870 19848
rect 20984 19839 21042 19845
rect 20984 19805 20996 19839
rect 21030 19836 21042 19839
rect 21358 19836 21364 19848
rect 21030 19808 21364 19836
rect 21030 19805 21042 19808
rect 20984 19799 21042 19805
rect 21358 19796 21364 19808
rect 21416 19796 21422 19848
rect 21726 19796 21732 19848
rect 21784 19836 21790 19848
rect 23400 19845 23428 19876
rect 24026 19864 24032 19916
rect 24084 19864 24090 19916
rect 24854 19864 24860 19916
rect 24912 19904 24918 19916
rect 25225 19907 25283 19913
rect 25225 19904 25237 19907
rect 24912 19876 25237 19904
rect 24912 19864 24918 19876
rect 25225 19873 25237 19876
rect 25271 19904 25283 19907
rect 25498 19904 25504 19916
rect 25271 19876 25504 19904
rect 25271 19873 25283 19876
rect 25225 19867 25283 19873
rect 25498 19864 25504 19876
rect 25556 19864 25562 19916
rect 23293 19839 23351 19845
rect 23293 19836 23305 19839
rect 21784 19808 23305 19836
rect 21784 19796 21790 19808
rect 23293 19805 23305 19808
rect 23339 19805 23351 19839
rect 23293 19799 23351 19805
rect 23385 19839 23443 19845
rect 23385 19805 23397 19839
rect 23431 19805 23443 19839
rect 23385 19799 23443 19805
rect 23569 19839 23627 19845
rect 23569 19805 23581 19839
rect 23615 19836 23627 19839
rect 24486 19836 24492 19848
rect 23615 19808 24492 19836
rect 23615 19805 23627 19808
rect 23569 19799 23627 19805
rect 15280 19771 15338 19777
rect 14292 19740 15240 19768
rect 12590 19731 12648 19737
rect 10781 19703 10839 19709
rect 10781 19669 10793 19703
rect 10827 19669 10839 19703
rect 10781 19663 10839 19669
rect 14461 19703 14519 19709
rect 14461 19669 14473 19703
rect 14507 19700 14519 19703
rect 15102 19700 15108 19712
rect 14507 19672 15108 19700
rect 14507 19669 14519 19672
rect 14461 19663 14519 19669
rect 15102 19660 15108 19672
rect 15160 19660 15166 19712
rect 15212 19700 15240 19740
rect 15280 19737 15292 19771
rect 15326 19768 15338 19771
rect 15470 19768 15476 19780
rect 15326 19740 15476 19768
rect 15326 19737 15338 19740
rect 15280 19731 15338 19737
rect 15470 19728 15476 19740
rect 15528 19728 15534 19780
rect 15562 19728 15568 19780
rect 15620 19768 15626 19780
rect 19334 19768 19340 19780
rect 15620 19740 19340 19768
rect 15620 19728 15626 19740
rect 19334 19728 19340 19740
rect 19392 19728 19398 19780
rect 19797 19771 19855 19777
rect 19797 19737 19809 19771
rect 19843 19768 19855 19771
rect 21450 19768 21456 19780
rect 19843 19740 21456 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 21450 19728 21456 19740
rect 21508 19728 21514 19780
rect 23308 19768 23336 19799
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 25774 19796 25780 19848
rect 25832 19796 25838 19848
rect 25976 19845 26004 19944
rect 42702 19932 42708 19984
rect 42760 19972 42766 19984
rect 42904 19972 42932 20012
rect 43438 20000 43444 20012
rect 43496 20000 43502 20052
rect 44637 20043 44695 20049
rect 44637 20009 44649 20043
rect 44683 20040 44695 20043
rect 44726 20040 44732 20052
rect 44683 20012 44732 20040
rect 44683 20009 44695 20012
rect 44637 20003 44695 20009
rect 44726 20000 44732 20012
rect 44784 20000 44790 20052
rect 47578 20000 47584 20052
rect 47636 20000 47642 20052
rect 48498 20000 48504 20052
rect 48556 20000 48562 20052
rect 50614 20000 50620 20052
rect 50672 20040 50678 20052
rect 51813 20043 51871 20049
rect 51813 20040 51825 20043
rect 50672 20012 51825 20040
rect 50672 20000 50678 20012
rect 51813 20009 51825 20012
rect 51859 20040 51871 20043
rect 51859 20012 53328 20040
rect 51859 20009 51871 20012
rect 51813 20003 51871 20009
rect 48406 19972 48412 19984
rect 42760 19944 42932 19972
rect 48148 19944 48412 19972
rect 42760 19932 42766 19944
rect 26789 19907 26847 19913
rect 26789 19873 26801 19907
rect 26835 19904 26847 19907
rect 28261 19907 28319 19913
rect 26835 19876 28212 19904
rect 26835 19873 26847 19876
rect 26789 19867 26847 19873
rect 25961 19839 26019 19845
rect 25961 19805 25973 19839
rect 26007 19805 26019 19839
rect 25961 19799 26019 19805
rect 26973 19839 27031 19845
rect 26973 19805 26985 19839
rect 27019 19836 27031 19839
rect 27019 19808 27660 19836
rect 27019 19805 27031 19808
rect 26973 19799 27031 19805
rect 24762 19768 24768 19780
rect 23308 19740 24768 19768
rect 24762 19728 24768 19740
rect 24820 19768 24826 19780
rect 24949 19771 25007 19777
rect 24949 19768 24961 19771
rect 24820 19740 24961 19768
rect 24820 19728 24826 19740
rect 24949 19737 24961 19740
rect 24995 19737 25007 19771
rect 24949 19731 25007 19737
rect 25041 19771 25099 19777
rect 25041 19737 25053 19771
rect 25087 19768 25099 19771
rect 27522 19768 27528 19780
rect 25087 19740 27528 19768
rect 25087 19737 25099 19740
rect 25041 19731 25099 19737
rect 27522 19728 27528 19740
rect 27580 19728 27586 19780
rect 15378 19700 15384 19712
rect 15212 19672 15384 19700
rect 15378 19660 15384 19672
rect 15436 19660 15442 19712
rect 18874 19660 18880 19712
rect 18932 19700 18938 19712
rect 19242 19700 19248 19712
rect 18932 19672 19248 19700
rect 18932 19660 18938 19672
rect 19242 19660 19248 19672
rect 19300 19660 19306 19712
rect 19889 19703 19947 19709
rect 19889 19669 19901 19703
rect 19935 19700 19947 19703
rect 21634 19700 21640 19712
rect 19935 19672 21640 19700
rect 19935 19669 19947 19672
rect 19889 19663 19947 19669
rect 21634 19660 21640 19672
rect 21692 19660 21698 19712
rect 22094 19660 22100 19712
rect 22152 19660 22158 19712
rect 25130 19660 25136 19712
rect 25188 19700 25194 19712
rect 26145 19703 26203 19709
rect 26145 19700 26157 19703
rect 25188 19672 26157 19700
rect 25188 19660 25194 19672
rect 26145 19669 26157 19672
rect 26191 19669 26203 19703
rect 26145 19663 26203 19669
rect 27157 19703 27215 19709
rect 27157 19669 27169 19703
rect 27203 19700 27215 19703
rect 27430 19700 27436 19712
rect 27203 19672 27436 19700
rect 27203 19669 27215 19672
rect 27157 19663 27215 19669
rect 27430 19660 27436 19672
rect 27488 19660 27494 19712
rect 27632 19709 27660 19808
rect 27982 19796 27988 19848
rect 28040 19836 28046 19848
rect 28077 19839 28135 19845
rect 28077 19836 28089 19839
rect 28040 19808 28089 19836
rect 28040 19796 28046 19808
rect 28077 19805 28089 19808
rect 28123 19805 28135 19839
rect 28184 19836 28212 19876
rect 28261 19873 28273 19907
rect 28307 19904 28319 19907
rect 28626 19904 28632 19916
rect 28307 19876 28632 19904
rect 28307 19873 28319 19876
rect 28261 19867 28319 19873
rect 28626 19864 28632 19876
rect 28684 19864 28690 19916
rect 32858 19904 32864 19916
rect 31726 19876 32864 19904
rect 30190 19836 30196 19848
rect 28184 19808 30196 19836
rect 28077 19799 28135 19805
rect 30190 19796 30196 19808
rect 30248 19796 30254 19848
rect 30282 19796 30288 19848
rect 30340 19836 30346 19848
rect 30653 19839 30711 19845
rect 30653 19836 30665 19839
rect 30340 19808 30665 19836
rect 30340 19796 30346 19808
rect 30653 19805 30665 19808
rect 30699 19836 30711 19839
rect 31726 19836 31754 19876
rect 32858 19864 32864 19876
rect 32916 19864 32922 19916
rect 37366 19864 37372 19916
rect 37424 19904 37430 19916
rect 38381 19907 38439 19913
rect 38381 19904 38393 19907
rect 37424 19876 38393 19904
rect 37424 19864 37430 19876
rect 38381 19873 38393 19876
rect 38427 19904 38439 19907
rect 45462 19904 45468 19916
rect 38427 19876 39712 19904
rect 38427 19873 38439 19876
rect 38381 19867 38439 19873
rect 30699 19808 31754 19836
rect 33128 19839 33186 19845
rect 30699 19805 30711 19808
rect 30653 19799 30711 19805
rect 33128 19805 33140 19839
rect 33174 19836 33186 19839
rect 33594 19836 33600 19848
rect 33174 19808 33600 19836
rect 33174 19805 33186 19808
rect 33128 19799 33186 19805
rect 33594 19796 33600 19808
rect 33652 19796 33658 19848
rect 35805 19839 35863 19845
rect 35805 19805 35817 19839
rect 35851 19836 35863 19839
rect 37182 19836 37188 19848
rect 35851 19808 37188 19836
rect 35851 19805 35863 19808
rect 35805 19799 35863 19805
rect 37182 19796 37188 19808
rect 37240 19796 37246 19848
rect 38105 19839 38163 19845
rect 38105 19836 38117 19839
rect 37292 19808 38117 19836
rect 30926 19777 30932 19780
rect 30920 19768 30932 19777
rect 30887 19740 30932 19768
rect 30920 19731 30932 19740
rect 30926 19728 30932 19731
rect 30984 19728 30990 19780
rect 36078 19777 36084 19780
rect 36072 19768 36084 19777
rect 36039 19740 36084 19768
rect 36072 19731 36084 19740
rect 36078 19728 36084 19731
rect 36136 19728 36142 19780
rect 27617 19703 27675 19709
rect 27617 19669 27629 19703
rect 27663 19669 27675 19703
rect 27617 19663 27675 19669
rect 27985 19703 28043 19709
rect 27985 19669 27997 19703
rect 28031 19700 28043 19703
rect 28074 19700 28080 19712
rect 28031 19672 28080 19700
rect 28031 19669 28043 19672
rect 27985 19663 28043 19669
rect 28074 19660 28080 19672
rect 28132 19660 28138 19712
rect 33962 19660 33968 19712
rect 34020 19700 34026 19712
rect 34241 19703 34299 19709
rect 34241 19700 34253 19703
rect 34020 19672 34253 19700
rect 34020 19660 34026 19672
rect 34241 19669 34253 19672
rect 34287 19669 34299 19703
rect 34241 19663 34299 19669
rect 34330 19660 34336 19712
rect 34388 19700 34394 19712
rect 36170 19700 36176 19712
rect 34388 19672 36176 19700
rect 34388 19660 34394 19672
rect 36170 19660 36176 19672
rect 36228 19660 36234 19712
rect 36262 19660 36268 19712
rect 36320 19700 36326 19712
rect 37185 19703 37243 19709
rect 37185 19700 37197 19703
rect 36320 19672 37197 19700
rect 36320 19660 36326 19672
rect 37185 19669 37197 19672
rect 37231 19700 37243 19703
rect 37292 19700 37320 19808
rect 38105 19805 38117 19808
rect 38151 19805 38163 19839
rect 38105 19799 38163 19805
rect 39684 19768 39712 19876
rect 44284 19876 45468 19904
rect 40218 19796 40224 19848
rect 40276 19836 40282 19848
rect 41325 19839 41383 19845
rect 41325 19836 41337 19839
rect 40276 19808 41337 19836
rect 40276 19796 40282 19808
rect 41325 19805 41337 19808
rect 41371 19836 41383 19839
rect 42886 19836 42892 19848
rect 41371 19808 42892 19836
rect 41371 19805 41383 19808
rect 41325 19799 41383 19805
rect 42886 19796 42892 19808
rect 42944 19836 42950 19848
rect 43257 19839 43315 19845
rect 43257 19836 43269 19839
rect 42944 19808 43269 19836
rect 42944 19796 42950 19808
rect 43257 19805 43269 19808
rect 43303 19836 43315 19839
rect 44284 19836 44312 19876
rect 45462 19864 45468 19876
rect 45520 19904 45526 19916
rect 48148 19913 48176 19944
rect 48406 19932 48412 19944
rect 48464 19972 48470 19984
rect 49234 19972 49240 19984
rect 48464 19944 49240 19972
rect 48464 19932 48470 19944
rect 49234 19932 49240 19944
rect 49292 19932 49298 19984
rect 53300 19972 53328 20012
rect 53558 20000 53564 20052
rect 53616 20040 53622 20052
rect 53745 20043 53803 20049
rect 53745 20040 53757 20043
rect 53616 20012 53757 20040
rect 53616 20000 53622 20012
rect 53745 20009 53757 20012
rect 53791 20009 53803 20043
rect 53745 20003 53803 20009
rect 53834 20000 53840 20052
rect 53892 20040 53898 20052
rect 55122 20040 55128 20052
rect 53892 20012 55128 20040
rect 53892 20000 53898 20012
rect 55122 20000 55128 20012
rect 55180 20000 55186 20052
rect 56042 20000 56048 20052
rect 56100 20000 56106 20052
rect 54938 19972 54944 19984
rect 53300 19944 54944 19972
rect 54938 19932 54944 19944
rect 54996 19932 55002 19984
rect 46201 19907 46259 19913
rect 46201 19904 46213 19907
rect 45520 19876 46213 19904
rect 45520 19864 45526 19876
rect 46201 19873 46213 19876
rect 46247 19873 46259 19907
rect 46201 19867 46259 19873
rect 48133 19907 48191 19913
rect 48133 19873 48145 19907
rect 48179 19873 48191 19907
rect 48133 19867 48191 19873
rect 48222 19864 48228 19916
rect 48280 19904 48286 19916
rect 50433 19907 50491 19913
rect 50433 19904 50445 19907
rect 48280 19876 50445 19904
rect 48280 19864 48286 19876
rect 50433 19873 50445 19876
rect 50479 19873 50491 19907
rect 50433 19867 50491 19873
rect 43303 19808 44312 19836
rect 43303 19805 43315 19808
rect 43257 19799 43315 19805
rect 45370 19796 45376 19848
rect 45428 19796 45434 19848
rect 45557 19839 45615 19845
rect 45557 19805 45569 19839
rect 45603 19836 45615 19839
rect 46290 19836 46296 19848
rect 45603 19808 46296 19836
rect 45603 19805 45615 19808
rect 45557 19799 45615 19805
rect 46290 19796 46296 19808
rect 46348 19796 46354 19848
rect 48314 19796 48320 19848
rect 48372 19796 48378 19848
rect 50448 19836 50476 19867
rect 52362 19864 52368 19916
rect 52420 19864 52426 19916
rect 56318 19904 56324 19916
rect 54588 19876 56324 19904
rect 50632 19836 50844 19838
rect 52380 19836 52408 19864
rect 50448 19810 52408 19836
rect 50448 19808 50660 19810
rect 50816 19808 52408 19810
rect 52454 19796 52460 19848
rect 52512 19836 52518 19848
rect 52621 19839 52679 19845
rect 52621 19836 52633 19839
rect 52512 19808 52633 19836
rect 52512 19796 52518 19808
rect 52621 19805 52633 19808
rect 52667 19805 52679 19839
rect 52621 19799 52679 19805
rect 54294 19796 54300 19848
rect 54352 19796 54358 19848
rect 54588 19845 54616 19876
rect 56318 19864 56324 19876
rect 56376 19864 56382 19916
rect 54573 19839 54631 19845
rect 54573 19805 54585 19839
rect 54619 19805 54631 19839
rect 54573 19799 54631 19805
rect 54665 19839 54723 19845
rect 54665 19805 54677 19839
rect 54711 19836 54723 19839
rect 55306 19836 55312 19848
rect 54711 19808 55312 19836
rect 54711 19805 54723 19808
rect 54665 19799 54723 19805
rect 55306 19796 55312 19808
rect 55364 19796 55370 19848
rect 55490 19796 55496 19848
rect 55548 19796 55554 19848
rect 55861 19839 55919 19845
rect 55861 19836 55873 19839
rect 55600 19808 55873 19836
rect 40494 19768 40500 19780
rect 38028 19740 39620 19768
rect 39684 19740 40500 19768
rect 37231 19672 37320 19700
rect 37737 19703 37795 19709
rect 37231 19669 37243 19672
rect 37185 19663 37243 19669
rect 37737 19669 37749 19703
rect 37783 19700 37795 19703
rect 38028 19700 38056 19740
rect 37783 19672 38056 19700
rect 37783 19669 37795 19672
rect 37737 19663 37795 19669
rect 38194 19660 38200 19712
rect 38252 19660 38258 19712
rect 39592 19700 39620 19740
rect 40494 19728 40500 19740
rect 40552 19728 40558 19780
rect 40678 19728 40684 19780
rect 40736 19728 40742 19780
rect 41592 19771 41650 19777
rect 40788 19740 41414 19768
rect 40788 19700 40816 19740
rect 39592 19672 40816 19700
rect 41386 19700 41414 19740
rect 41592 19737 41604 19771
rect 41638 19768 41650 19771
rect 41782 19768 41788 19780
rect 41638 19740 41788 19768
rect 41638 19737 41650 19740
rect 41592 19731 41650 19737
rect 41782 19728 41788 19740
rect 41840 19728 41846 19780
rect 41892 19740 42932 19768
rect 41892 19700 41920 19740
rect 41386 19672 41920 19700
rect 42904 19700 42932 19740
rect 42978 19728 42984 19780
rect 43036 19768 43042 19780
rect 43502 19771 43560 19777
rect 43502 19768 43514 19771
rect 43036 19740 43514 19768
rect 43036 19728 43042 19740
rect 43502 19737 43514 19740
rect 43548 19737 43560 19771
rect 43502 19731 43560 19737
rect 45741 19771 45799 19777
rect 45741 19737 45753 19771
rect 45787 19768 45799 19771
rect 46446 19771 46504 19777
rect 46446 19768 46458 19771
rect 45787 19740 46458 19768
rect 45787 19737 45799 19740
rect 45741 19731 45799 19737
rect 46446 19737 46458 19740
rect 46492 19737 46504 19771
rect 46446 19731 46504 19737
rect 50522 19728 50528 19780
rect 50580 19768 50586 19780
rect 50678 19771 50736 19777
rect 50678 19768 50690 19771
rect 50580 19740 50690 19768
rect 50580 19728 50586 19740
rect 50678 19737 50690 19740
rect 50724 19737 50736 19771
rect 52362 19768 52368 19780
rect 50678 19731 50736 19737
rect 51046 19740 52368 19768
rect 45554 19700 45560 19712
rect 42904 19672 45560 19700
rect 45554 19660 45560 19672
rect 45612 19660 45618 19712
rect 45922 19660 45928 19712
rect 45980 19700 45986 19712
rect 51046 19700 51074 19740
rect 52362 19728 52368 19740
rect 52420 19728 52426 19780
rect 54481 19771 54539 19777
rect 54481 19737 54493 19771
rect 54527 19737 54539 19771
rect 55324 19768 55352 19796
rect 55600 19768 55628 19808
rect 55861 19805 55873 19808
rect 55907 19805 55919 19839
rect 55861 19799 55919 19805
rect 55950 19796 55956 19848
rect 56008 19836 56014 19848
rect 56873 19839 56931 19845
rect 56873 19836 56885 19839
rect 56008 19808 56885 19836
rect 56008 19796 56014 19808
rect 56873 19805 56885 19808
rect 56919 19805 56931 19839
rect 56873 19799 56931 19805
rect 56962 19796 56968 19848
rect 57020 19836 57026 19848
rect 57129 19839 57187 19845
rect 57129 19836 57141 19839
rect 57020 19808 57141 19836
rect 57020 19796 57026 19808
rect 57129 19805 57141 19808
rect 57175 19805 57187 19839
rect 57129 19799 57187 19805
rect 55324 19740 55628 19768
rect 55677 19771 55735 19777
rect 54481 19731 54539 19737
rect 55677 19737 55689 19771
rect 55723 19737 55735 19771
rect 55677 19731 55735 19737
rect 55769 19771 55827 19777
rect 55769 19737 55781 19771
rect 55815 19768 55827 19771
rect 55815 19740 58296 19768
rect 55815 19737 55827 19740
rect 55769 19731 55827 19737
rect 45980 19672 51074 19700
rect 54496 19700 54524 19731
rect 54662 19700 54668 19712
rect 54496 19672 54668 19700
rect 45980 19660 45986 19672
rect 54662 19660 54668 19672
rect 54720 19660 54726 19712
rect 54754 19660 54760 19712
rect 54812 19700 54818 19712
rect 54849 19703 54907 19709
rect 54849 19700 54861 19703
rect 54812 19672 54861 19700
rect 54812 19660 54818 19672
rect 54849 19669 54861 19672
rect 54895 19669 54907 19703
rect 54849 19663 54907 19669
rect 55122 19660 55128 19712
rect 55180 19700 55186 19712
rect 55692 19700 55720 19731
rect 57072 19712 57100 19740
rect 55180 19672 55720 19700
rect 55180 19660 55186 19672
rect 57054 19660 57060 19712
rect 57112 19660 57118 19712
rect 58268 19709 58296 19740
rect 58253 19703 58311 19709
rect 58253 19669 58265 19703
rect 58299 19669 58311 19703
rect 58253 19663 58311 19669
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 7558 19496 7564 19508
rect 2746 19468 7564 19496
rect 934 19388 940 19440
rect 992 19428 998 19440
rect 1857 19431 1915 19437
rect 1857 19428 1869 19431
rect 992 19400 1869 19428
rect 992 19388 998 19400
rect 1857 19397 1869 19400
rect 1903 19397 1915 19431
rect 1857 19391 1915 19397
rect 1581 19363 1639 19369
rect 1581 19329 1593 19363
rect 1627 19360 1639 19363
rect 2746 19360 2774 19468
rect 7558 19456 7564 19468
rect 7616 19456 7622 19508
rect 8205 19499 8263 19505
rect 8205 19465 8217 19499
rect 8251 19496 8263 19499
rect 9674 19496 9680 19508
rect 8251 19468 9680 19496
rect 8251 19465 8263 19468
rect 8205 19459 8263 19465
rect 9674 19456 9680 19468
rect 9732 19456 9738 19508
rect 10134 19456 10140 19508
rect 10192 19456 10198 19508
rect 10612 19468 11100 19496
rect 10612 19428 10640 19468
rect 11072 19440 11100 19468
rect 11146 19456 11152 19508
rect 11204 19456 11210 19508
rect 13817 19499 13875 19505
rect 13817 19465 13829 19499
rect 13863 19496 13875 19499
rect 15749 19499 15807 19505
rect 13863 19468 15700 19496
rect 13863 19465 13875 19468
rect 13817 19459 13875 19465
rect 1627 19332 2774 19360
rect 6840 19400 10640 19428
rect 1627 19329 1639 19332
rect 1581 19323 1639 19329
rect 6086 19252 6092 19304
rect 6144 19292 6150 19304
rect 6840 19301 6868 19400
rect 7098 19369 7104 19372
rect 7092 19360 7104 19369
rect 7059 19332 7104 19360
rect 7092 19323 7104 19332
rect 7098 19320 7104 19323
rect 7156 19320 7162 19372
rect 8772 19369 8800 19400
rect 10686 19388 10692 19440
rect 10744 19388 10750 19440
rect 11054 19388 11060 19440
rect 11112 19428 11118 19440
rect 12066 19428 12072 19440
rect 11112 19400 12072 19428
rect 11112 19388 11118 19400
rect 12066 19388 12072 19400
rect 12124 19428 12130 19440
rect 12342 19428 12348 19440
rect 12124 19400 12348 19428
rect 12124 19388 12130 19400
rect 12342 19388 12348 19400
rect 12400 19428 12406 19440
rect 15562 19428 15568 19440
rect 12400 19400 14412 19428
rect 12400 19388 12406 19400
rect 8757 19363 8815 19369
rect 8757 19329 8769 19363
rect 8803 19329 8815 19363
rect 8757 19323 8815 19329
rect 9024 19363 9082 19369
rect 9024 19329 9036 19363
rect 9070 19360 9082 19363
rect 10042 19360 10048 19372
rect 9070 19332 10048 19360
rect 9070 19329 9082 19332
rect 9024 19323 9082 19329
rect 10042 19320 10048 19332
rect 10100 19320 10106 19372
rect 11698 19320 11704 19372
rect 11756 19320 11762 19372
rect 12452 19369 12480 19400
rect 14384 19372 14412 19400
rect 14476 19400 15568 19428
rect 12437 19363 12495 19369
rect 12437 19329 12449 19363
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 12704 19363 12762 19369
rect 12704 19329 12716 19363
rect 12750 19360 12762 19363
rect 14182 19360 14188 19372
rect 12750 19332 14188 19360
rect 12750 19329 12762 19332
rect 12704 19323 12762 19329
rect 14182 19320 14188 19332
rect 14240 19320 14246 19372
rect 14366 19320 14372 19372
rect 14424 19320 14430 19372
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6144 19264 6837 19292
rect 6144 19252 6150 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 14476 19292 14504 19400
rect 15562 19388 15568 19400
rect 15620 19388 15626 19440
rect 15672 19428 15700 19468
rect 15749 19465 15761 19499
rect 15795 19496 15807 19499
rect 18138 19496 18144 19508
rect 15795 19468 18144 19496
rect 15795 19465 15807 19468
rect 15749 19459 15807 19465
rect 18138 19456 18144 19468
rect 18196 19456 18202 19508
rect 19061 19499 19119 19505
rect 19061 19465 19073 19499
rect 19107 19496 19119 19499
rect 19150 19496 19156 19508
rect 19107 19468 19156 19496
rect 19107 19465 19119 19468
rect 19061 19459 19119 19465
rect 19150 19456 19156 19468
rect 19208 19456 19214 19508
rect 21634 19496 21640 19508
rect 20180 19468 21640 19496
rect 20180 19428 20208 19468
rect 21634 19456 21640 19468
rect 21692 19456 21698 19508
rect 24762 19456 24768 19508
rect 24820 19456 24826 19508
rect 25590 19456 25596 19508
rect 25648 19496 25654 19508
rect 25648 19468 30696 19496
rect 25648 19456 25654 19468
rect 26510 19428 26516 19440
rect 15672 19400 20208 19428
rect 23584 19400 26516 19428
rect 14636 19363 14694 19369
rect 14636 19329 14648 19363
rect 14682 19360 14694 19363
rect 15194 19360 15200 19372
rect 14682 19332 15200 19360
rect 14682 19329 14694 19332
rect 14636 19323 14694 19329
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 16574 19320 16580 19372
rect 16632 19360 16638 19372
rect 17293 19363 17351 19369
rect 17293 19360 17305 19363
rect 16632 19332 17305 19360
rect 16632 19320 16638 19332
rect 17293 19329 17305 19332
rect 17339 19329 17351 19363
rect 17293 19323 17351 19329
rect 19150 19320 19156 19372
rect 19208 19320 19214 19372
rect 19245 19363 19303 19369
rect 19245 19329 19257 19363
rect 19291 19360 19303 19363
rect 19291 19332 20024 19360
rect 19291 19329 19303 19332
rect 19245 19323 19303 19329
rect 6825 19255 6883 19261
rect 13464 19264 14504 19292
rect 10962 19184 10968 19236
rect 11020 19184 11026 19236
rect 11422 19184 11428 19236
rect 11480 19224 11486 19236
rect 11480 19196 12020 19224
rect 11480 19184 11486 19196
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 11885 19159 11943 19165
rect 11885 19156 11897 19159
rect 9732 19128 11897 19156
rect 9732 19116 9738 19128
rect 11885 19125 11897 19128
rect 11931 19125 11943 19159
rect 11992 19156 12020 19196
rect 12802 19156 12808 19168
rect 11992 19128 12808 19156
rect 11885 19119 11943 19125
rect 12802 19116 12808 19128
rect 12860 19156 12866 19168
rect 13354 19156 13360 19168
rect 12860 19128 13360 19156
rect 12860 19116 12866 19128
rect 13354 19116 13360 19128
rect 13412 19156 13418 19168
rect 13464 19156 13492 19264
rect 17034 19252 17040 19304
rect 17092 19252 17098 19304
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19429 19295 19487 19301
rect 19429 19292 19441 19295
rect 19392 19264 19441 19292
rect 19392 19252 19398 19264
rect 19429 19261 19441 19264
rect 19475 19261 19487 19295
rect 19996 19292 20024 19332
rect 20070 19320 20076 19372
rect 20128 19320 20134 19372
rect 20162 19320 20168 19372
rect 20220 19320 20226 19372
rect 20340 19363 20398 19369
rect 20340 19329 20352 19363
rect 20386 19360 20398 19363
rect 20898 19360 20904 19372
rect 20386 19332 20904 19360
rect 20386 19329 20398 19332
rect 20340 19323 20398 19329
rect 20898 19320 20904 19332
rect 20956 19320 20962 19372
rect 21174 19320 21180 19372
rect 21232 19360 21238 19372
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 21232 19332 22017 19360
rect 21232 19320 21238 19332
rect 22005 19329 22017 19332
rect 22051 19360 22063 19363
rect 22094 19360 22100 19372
rect 22051 19332 22100 19360
rect 22051 19329 22063 19332
rect 22005 19323 22063 19329
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 23382 19320 23388 19372
rect 23440 19360 23446 19372
rect 23584 19360 23612 19400
rect 26510 19388 26516 19400
rect 26568 19428 26574 19440
rect 26568 19400 27476 19428
rect 26568 19388 26574 19400
rect 23440 19332 23612 19360
rect 23652 19363 23710 19369
rect 23440 19320 23446 19332
rect 23652 19329 23664 19363
rect 23698 19360 23710 19363
rect 25130 19360 25136 19372
rect 23698 19332 25136 19360
rect 23698 19329 23710 19332
rect 23652 19323 23710 19329
rect 25130 19320 25136 19332
rect 25188 19320 25194 19372
rect 25590 19320 25596 19372
rect 25648 19320 25654 19372
rect 25774 19320 25780 19372
rect 25832 19360 25838 19372
rect 25958 19360 25964 19372
rect 25832 19332 25964 19360
rect 25832 19320 25838 19332
rect 25958 19320 25964 19332
rect 26016 19320 26022 19372
rect 26142 19320 26148 19372
rect 26200 19360 26206 19372
rect 27448 19369 27476 19400
rect 27522 19388 27528 19440
rect 27580 19428 27586 19440
rect 27678 19431 27736 19437
rect 27678 19428 27690 19431
rect 27580 19400 27690 19428
rect 27580 19388 27586 19400
rect 27678 19397 27690 19400
rect 27724 19397 27736 19431
rect 27678 19391 27736 19397
rect 26329 19363 26387 19369
rect 26329 19360 26341 19363
rect 26200 19332 26341 19360
rect 26200 19320 26206 19332
rect 26329 19329 26341 19332
rect 26375 19329 26387 19363
rect 26329 19323 26387 19329
rect 27433 19363 27491 19369
rect 27433 19329 27445 19363
rect 27479 19329 27491 19363
rect 27433 19323 27491 19329
rect 30282 19320 30288 19372
rect 30340 19320 30346 19372
rect 30558 19369 30564 19372
rect 30552 19323 30564 19369
rect 30558 19320 30564 19323
rect 30616 19320 30622 19372
rect 30668 19360 30696 19468
rect 31662 19456 31668 19508
rect 31720 19456 31726 19508
rect 33410 19456 33416 19508
rect 33468 19496 33474 19508
rect 33597 19499 33655 19505
rect 33597 19496 33609 19499
rect 33468 19468 33609 19496
rect 33468 19456 33474 19468
rect 33597 19465 33609 19468
rect 33643 19465 33655 19499
rect 33597 19459 33655 19465
rect 33962 19456 33968 19508
rect 34020 19456 34026 19508
rect 34054 19456 34060 19508
rect 34112 19456 34118 19508
rect 35894 19456 35900 19508
rect 35952 19456 35958 19508
rect 40494 19456 40500 19508
rect 40552 19496 40558 19508
rect 41322 19496 41328 19508
rect 40552 19468 41328 19496
rect 40552 19456 40558 19468
rect 41322 19456 41328 19468
rect 41380 19496 41386 19508
rect 41380 19468 43300 19496
rect 41380 19456 41386 19468
rect 31386 19388 31392 19440
rect 31444 19428 31450 19440
rect 36262 19428 36268 19440
rect 31444 19400 36268 19428
rect 31444 19388 31450 19400
rect 36262 19388 36268 19400
rect 36320 19388 36326 19440
rect 42061 19431 42119 19437
rect 42061 19397 42073 19431
rect 42107 19428 42119 19431
rect 43134 19431 43192 19437
rect 43134 19428 43146 19431
rect 42107 19400 43146 19428
rect 42107 19397 42119 19400
rect 42061 19391 42119 19397
rect 43134 19397 43146 19400
rect 43180 19397 43192 19431
rect 43272 19428 43300 19468
rect 43346 19456 43352 19508
rect 43404 19496 43410 19508
rect 44269 19499 44327 19505
rect 44269 19496 44281 19499
rect 43404 19468 44281 19496
rect 43404 19456 43410 19468
rect 44269 19465 44281 19468
rect 44315 19496 44327 19499
rect 45922 19496 45928 19508
rect 44315 19468 45928 19496
rect 44315 19465 44327 19468
rect 44269 19459 44327 19465
rect 45922 19456 45928 19468
rect 45980 19456 45986 19508
rect 46842 19456 46848 19508
rect 46900 19456 46906 19508
rect 46934 19456 46940 19508
rect 46992 19496 46998 19508
rect 49694 19496 49700 19508
rect 46992 19468 49700 19496
rect 46992 19456 46998 19468
rect 49694 19456 49700 19468
rect 49752 19496 49758 19508
rect 49752 19468 49924 19496
rect 49752 19456 49758 19468
rect 43622 19428 43628 19440
rect 43272 19400 43628 19428
rect 43134 19391 43192 19397
rect 43622 19388 43628 19400
rect 43680 19388 43686 19440
rect 47854 19388 47860 19440
rect 47912 19428 47918 19440
rect 48041 19431 48099 19437
rect 48041 19428 48053 19431
rect 47912 19400 48053 19428
rect 47912 19388 47918 19400
rect 48041 19397 48053 19400
rect 48087 19428 48099 19431
rect 48130 19428 48136 19440
rect 48087 19400 48136 19428
rect 48087 19397 48099 19400
rect 48041 19391 48099 19397
rect 48130 19388 48136 19400
rect 48188 19388 48194 19440
rect 32490 19360 32496 19372
rect 30668 19332 32496 19360
rect 32490 19320 32496 19332
rect 32548 19360 32554 19372
rect 33962 19360 33968 19372
rect 32548 19332 33968 19360
rect 32548 19320 32554 19332
rect 33962 19320 33968 19332
rect 34020 19320 34026 19372
rect 36354 19320 36360 19372
rect 36412 19320 36418 19372
rect 39206 19360 39212 19372
rect 37568 19332 39212 19360
rect 20180 19292 20208 19320
rect 19996 19264 20208 19292
rect 19429 19255 19487 19261
rect 21358 19252 21364 19304
rect 21416 19292 21422 19304
rect 22462 19292 22468 19304
rect 21416 19264 22468 19292
rect 21416 19252 21422 19264
rect 22462 19252 22468 19264
rect 22520 19252 22526 19304
rect 25406 19252 25412 19304
rect 25464 19292 25470 19304
rect 34241 19295 34299 19301
rect 25464 19264 27476 19292
rect 25464 19252 25470 19264
rect 27448 19236 27476 19264
rect 34241 19261 34253 19295
rect 34287 19292 34299 19295
rect 36538 19292 36544 19304
rect 34287 19264 36544 19292
rect 34287 19261 34299 19264
rect 34241 19255 34299 19261
rect 36538 19252 36544 19264
rect 36596 19292 36602 19304
rect 37568 19292 37596 19332
rect 39206 19320 39212 19332
rect 39264 19320 39270 19372
rect 41690 19360 41696 19372
rect 41386 19334 41696 19360
rect 41340 19332 41696 19334
rect 41340 19306 41414 19332
rect 41690 19320 41696 19332
rect 41748 19320 41754 19372
rect 41874 19320 41880 19372
rect 41932 19320 41938 19372
rect 42886 19320 42892 19372
rect 42944 19320 42950 19372
rect 45462 19320 45468 19372
rect 45520 19320 45526 19372
rect 45738 19369 45744 19372
rect 45732 19323 45744 19369
rect 45738 19320 45744 19323
rect 45796 19320 45802 19372
rect 47670 19320 47676 19372
rect 47728 19360 47734 19372
rect 47765 19363 47823 19369
rect 47765 19360 47777 19363
rect 47728 19332 47777 19360
rect 47728 19320 47734 19332
rect 47765 19329 47777 19332
rect 47811 19329 47823 19363
rect 47765 19323 47823 19329
rect 49786 19320 49792 19372
rect 49844 19320 49850 19372
rect 49896 19366 49924 19468
rect 51626 19456 51632 19508
rect 51684 19456 51690 19508
rect 54941 19499 54999 19505
rect 54941 19465 54953 19499
rect 54987 19496 54999 19499
rect 55030 19496 55036 19508
rect 54987 19468 55036 19496
rect 54987 19465 54999 19468
rect 54941 19459 54999 19465
rect 55030 19456 55036 19468
rect 55088 19456 55094 19508
rect 50522 19388 50528 19440
rect 50580 19428 50586 19440
rect 50580 19400 51120 19428
rect 50580 19388 50586 19400
rect 51092 19369 51120 19400
rect 51258 19388 51264 19440
rect 51316 19388 51322 19440
rect 51353 19431 51411 19437
rect 51353 19397 51365 19431
rect 51399 19428 51411 19431
rect 53558 19428 53564 19440
rect 51399 19400 53564 19428
rect 51399 19397 51411 19400
rect 51353 19391 51411 19397
rect 53558 19388 53564 19400
rect 53616 19388 53622 19440
rect 49973 19366 50031 19369
rect 49896 19363 50031 19366
rect 49896 19338 49985 19363
rect 49973 19329 49985 19338
rect 50019 19329 50031 19363
rect 49973 19323 50031 19329
rect 50065 19363 50123 19369
rect 50065 19329 50077 19363
rect 50111 19329 50123 19363
rect 50065 19323 50123 19329
rect 50181 19363 50239 19369
rect 50181 19329 50193 19363
rect 50227 19360 50239 19363
rect 51077 19363 51135 19369
rect 50227 19358 50246 19360
rect 50356 19358 51028 19360
rect 50227 19332 51028 19358
rect 50227 19330 50384 19332
rect 50227 19329 50239 19330
rect 50181 19323 50239 19329
rect 40034 19292 40040 19304
rect 36596 19264 37596 19292
rect 37624 19264 40040 19292
rect 36596 19252 36602 19264
rect 18322 19184 18328 19236
rect 18380 19224 18386 19236
rect 18877 19227 18935 19233
rect 18877 19224 18889 19227
rect 18380 19196 18889 19224
rect 18380 19184 18386 19196
rect 18877 19193 18889 19196
rect 18923 19224 18935 19227
rect 18923 19196 20116 19224
rect 18923 19193 18935 19196
rect 18877 19187 18935 19193
rect 13412 19128 13492 19156
rect 13412 19116 13418 19128
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 17310 19156 17316 19168
rect 13964 19128 17316 19156
rect 13964 19116 13970 19128
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 18417 19159 18475 19165
rect 18417 19125 18429 19159
rect 18463 19156 18475 19159
rect 19886 19156 19892 19168
rect 18463 19128 19892 19156
rect 18463 19125 18475 19128
rect 18417 19119 18475 19125
rect 19886 19116 19892 19128
rect 19944 19116 19950 19168
rect 20088 19156 20116 19196
rect 21910 19184 21916 19236
rect 21968 19224 21974 19236
rect 26513 19227 26571 19233
rect 26513 19224 26525 19227
rect 21968 19196 23428 19224
rect 21968 19184 21974 19196
rect 21082 19156 21088 19168
rect 20088 19128 21088 19156
rect 21082 19116 21088 19128
rect 21140 19116 21146 19168
rect 21174 19116 21180 19168
rect 21232 19156 21238 19168
rect 21453 19159 21511 19165
rect 21453 19156 21465 19159
rect 21232 19128 21465 19156
rect 21232 19116 21238 19128
rect 21453 19125 21465 19128
rect 21499 19125 21511 19159
rect 21453 19119 21511 19125
rect 21542 19116 21548 19168
rect 21600 19156 21606 19168
rect 22189 19159 22247 19165
rect 22189 19156 22201 19159
rect 21600 19128 22201 19156
rect 21600 19116 21606 19128
rect 22189 19125 22201 19128
rect 22235 19125 22247 19159
rect 23400 19156 23428 19196
rect 24320 19196 26525 19224
rect 24320 19156 24348 19196
rect 26513 19193 26525 19196
rect 26559 19193 26571 19227
rect 26513 19187 26571 19193
rect 27430 19184 27436 19236
rect 27488 19184 27494 19236
rect 23400 19128 24348 19156
rect 22189 19119 22247 19125
rect 24486 19116 24492 19168
rect 24544 19156 24550 19168
rect 25222 19156 25228 19168
rect 24544 19128 25228 19156
rect 24544 19116 24550 19128
rect 25222 19116 25228 19128
rect 25280 19116 25286 19168
rect 25774 19116 25780 19168
rect 25832 19116 25838 19168
rect 28074 19116 28080 19168
rect 28132 19156 28138 19168
rect 28813 19159 28871 19165
rect 28813 19156 28825 19159
rect 28132 19128 28825 19156
rect 28132 19116 28138 19128
rect 28813 19125 28825 19128
rect 28859 19125 28871 19159
rect 28813 19119 28871 19125
rect 29270 19116 29276 19168
rect 29328 19156 29334 19168
rect 37624 19156 37652 19264
rect 40034 19252 40040 19264
rect 40092 19252 40098 19304
rect 40494 19252 40500 19304
rect 40552 19292 40558 19304
rect 41340 19292 41368 19306
rect 40552 19264 41368 19292
rect 41708 19292 41736 19320
rect 42334 19292 42340 19304
rect 41708 19264 42340 19292
rect 40552 19252 40558 19264
rect 42334 19252 42340 19264
rect 42392 19252 42398 19304
rect 50080 19292 50108 19323
rect 51000 19304 51028 19332
rect 51077 19329 51089 19363
rect 51123 19329 51135 19363
rect 51077 19323 51135 19329
rect 51445 19363 51503 19369
rect 51445 19329 51457 19363
rect 51491 19329 51503 19363
rect 51445 19323 51503 19329
rect 50614 19292 50620 19304
rect 50080 19264 50620 19292
rect 50614 19252 50620 19264
rect 50672 19252 50678 19304
rect 50982 19252 50988 19304
rect 51040 19292 51046 19304
rect 51460 19292 51488 19323
rect 54754 19320 54760 19372
rect 54812 19320 54818 19372
rect 51040 19264 51488 19292
rect 54573 19295 54631 19301
rect 51040 19252 51046 19264
rect 54573 19261 54585 19295
rect 54619 19261 54631 19295
rect 54573 19255 54631 19261
rect 49694 19224 49700 19236
rect 44192 19196 44404 19224
rect 29328 19128 37652 19156
rect 29328 19116 29334 19128
rect 37826 19116 37832 19168
rect 37884 19156 37890 19168
rect 40954 19156 40960 19168
rect 37884 19128 40960 19156
rect 37884 19116 37890 19128
rect 40954 19116 40960 19128
rect 41012 19156 41018 19168
rect 44192 19156 44220 19196
rect 41012 19128 44220 19156
rect 44376 19156 44404 19196
rect 46400 19196 49700 19224
rect 46400 19156 46428 19196
rect 49694 19184 49700 19196
rect 49752 19184 49758 19236
rect 51442 19184 51448 19236
rect 51500 19224 51506 19236
rect 54588 19224 54616 19255
rect 55490 19224 55496 19236
rect 51500 19196 55496 19224
rect 51500 19184 51506 19196
rect 55490 19184 55496 19196
rect 55548 19224 55554 19236
rect 55674 19224 55680 19236
rect 55548 19196 55680 19224
rect 55548 19184 55554 19196
rect 55674 19184 55680 19196
rect 55732 19184 55738 19236
rect 44376 19128 46428 19156
rect 41012 19116 41018 19128
rect 50154 19116 50160 19168
rect 50212 19156 50218 19168
rect 50341 19159 50399 19165
rect 50341 19156 50353 19159
rect 50212 19128 50353 19156
rect 50212 19116 50218 19128
rect 50341 19125 50353 19128
rect 50387 19125 50399 19159
rect 50341 19119 50399 19125
rect 50430 19116 50436 19168
rect 50488 19156 50494 19168
rect 58618 19156 58624 19168
rect 50488 19128 58624 19156
rect 50488 19116 50494 19128
rect 58618 19116 58624 19128
rect 58676 19116 58682 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 8021 18955 8079 18961
rect 8021 18921 8033 18955
rect 8067 18952 8079 18955
rect 8386 18952 8392 18964
rect 8067 18924 8392 18952
rect 8067 18921 8079 18924
rect 8021 18915 8079 18921
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 9582 18952 9588 18964
rect 9140 18924 9588 18952
rect 7469 18887 7527 18893
rect 7469 18853 7481 18887
rect 7515 18884 7527 18887
rect 9030 18884 9036 18896
rect 7515 18856 9036 18884
rect 7515 18853 7527 18856
rect 7469 18847 7527 18853
rect 9030 18844 9036 18856
rect 9088 18844 9094 18896
rect 9140 18893 9168 18924
rect 9582 18912 9588 18924
rect 9640 18912 9646 18964
rect 10226 18912 10232 18964
rect 10284 18952 10290 18964
rect 10597 18955 10655 18961
rect 10597 18952 10609 18955
rect 10284 18924 10609 18952
rect 10284 18912 10290 18924
rect 10597 18921 10609 18924
rect 10643 18921 10655 18955
rect 10597 18915 10655 18921
rect 11517 18955 11575 18961
rect 11517 18921 11529 18955
rect 11563 18952 11575 18955
rect 11606 18952 11612 18964
rect 11563 18924 11612 18952
rect 11563 18921 11575 18924
rect 11517 18915 11575 18921
rect 11606 18912 11612 18924
rect 11664 18912 11670 18964
rect 13449 18955 13507 18961
rect 13449 18921 13461 18955
rect 13495 18952 13507 18955
rect 13906 18952 13912 18964
rect 13495 18924 13912 18952
rect 13495 18921 13507 18924
rect 13449 18915 13507 18921
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 16574 18912 16580 18964
rect 16632 18912 16638 18964
rect 18782 18912 18788 18964
rect 18840 18912 18846 18964
rect 20898 18912 20904 18964
rect 20956 18952 20962 18964
rect 20993 18955 21051 18961
rect 20993 18952 21005 18955
rect 20956 18924 21005 18952
rect 20956 18912 20962 18924
rect 20993 18921 21005 18924
rect 21039 18921 21051 18955
rect 20993 18915 21051 18921
rect 21082 18912 21088 18964
rect 21140 18952 21146 18964
rect 22373 18955 22431 18961
rect 22373 18952 22385 18955
rect 21140 18924 22385 18952
rect 21140 18912 21146 18924
rect 22373 18921 22385 18924
rect 22419 18921 22431 18955
rect 25774 18952 25780 18964
rect 22373 18915 22431 18921
rect 23952 18924 25780 18952
rect 9125 18887 9183 18893
rect 9125 18853 9137 18887
rect 9171 18853 9183 18887
rect 9125 18847 9183 18853
rect 9306 18844 9312 18896
rect 9364 18884 9370 18896
rect 11882 18884 11888 18896
rect 9364 18856 11888 18884
rect 9364 18844 9370 18856
rect 11882 18844 11888 18856
rect 11940 18844 11946 18896
rect 15841 18887 15899 18893
rect 15841 18884 15853 18887
rect 14476 18856 15853 18884
rect 6086 18776 6092 18828
rect 6144 18776 6150 18828
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 8128 18788 9689 18816
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18748 1639 18751
rect 5258 18748 5264 18760
rect 1627 18720 5264 18748
rect 1627 18717 1639 18720
rect 1581 18711 1639 18717
rect 5258 18708 5264 18720
rect 5316 18708 5322 18760
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18748 5411 18751
rect 7098 18748 7104 18760
rect 5399 18720 7104 18748
rect 5399 18717 5411 18720
rect 5353 18711 5411 18717
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 934 18640 940 18692
rect 992 18680 998 18692
rect 1857 18683 1915 18689
rect 1857 18680 1869 18683
rect 992 18652 1869 18680
rect 992 18640 998 18652
rect 1857 18649 1869 18652
rect 1903 18649 1915 18683
rect 1857 18643 1915 18649
rect 6356 18683 6414 18689
rect 6356 18649 6368 18683
rect 6402 18680 6414 18683
rect 6730 18680 6736 18692
rect 6402 18652 6736 18680
rect 6402 18649 6414 18652
rect 6356 18643 6414 18649
rect 6730 18640 6736 18652
rect 6788 18640 6794 18692
rect 6914 18640 6920 18692
rect 6972 18680 6978 18692
rect 8128 18680 8156 18788
rect 9677 18785 9689 18788
rect 9723 18785 9735 18819
rect 9677 18779 9735 18785
rect 10226 18776 10232 18828
rect 10284 18776 10290 18828
rect 12066 18776 12072 18828
rect 12124 18776 12130 18828
rect 8202 18708 8208 18760
rect 8260 18708 8266 18760
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18717 8355 18751
rect 8297 18711 8355 18717
rect 6972 18652 8156 18680
rect 8312 18680 8340 18711
rect 8386 18708 8392 18760
rect 8444 18708 8450 18760
rect 8481 18751 8539 18757
rect 8481 18717 8493 18751
rect 8527 18748 8539 18751
rect 10134 18748 10140 18760
rect 8527 18720 10140 18748
rect 8527 18717 8539 18720
rect 8481 18711 8539 18717
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18717 10379 18751
rect 10321 18711 10379 18717
rect 9401 18683 9459 18689
rect 9401 18680 9413 18683
rect 8312 18652 9413 18680
rect 6972 18640 6978 18652
rect 9401 18649 9413 18652
rect 9447 18680 9459 18683
rect 10042 18680 10048 18692
rect 9447 18652 10048 18680
rect 9447 18649 9459 18652
rect 9401 18643 9459 18649
rect 10042 18640 10048 18652
rect 10100 18640 10106 18692
rect 10336 18680 10364 18711
rect 11422 18708 11428 18760
rect 11480 18708 11486 18760
rect 11609 18751 11667 18757
rect 11609 18717 11621 18751
rect 11655 18748 11667 18751
rect 13170 18748 13176 18760
rect 11655 18720 13176 18748
rect 11655 18717 11667 18720
rect 11609 18711 11667 18717
rect 13170 18708 13176 18720
rect 13228 18708 13234 18760
rect 14476 18757 14504 18856
rect 15841 18853 15853 18856
rect 15887 18853 15899 18887
rect 18049 18887 18107 18893
rect 18049 18884 18061 18887
rect 15841 18847 15899 18853
rect 15948 18856 18061 18884
rect 14553 18819 14611 18825
rect 14553 18785 14565 18819
rect 14599 18785 14611 18819
rect 14553 18779 14611 18785
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18717 14519 18751
rect 14568 18748 14596 18779
rect 14826 18776 14832 18828
rect 14884 18776 14890 18828
rect 15562 18748 15568 18760
rect 14568 18720 15568 18748
rect 14461 18711 14519 18717
rect 15562 18708 15568 18720
rect 15620 18708 15626 18760
rect 15657 18751 15715 18757
rect 15657 18717 15669 18751
rect 15703 18748 15715 18751
rect 15948 18748 15976 18856
rect 18049 18853 18061 18856
rect 18095 18853 18107 18887
rect 23952 18884 23980 18924
rect 25774 18912 25780 18924
rect 25832 18912 25838 18964
rect 29178 18952 29184 18964
rect 26436 18924 29184 18952
rect 18049 18847 18107 18853
rect 19536 18856 23980 18884
rect 19429 18819 19487 18825
rect 19429 18816 19441 18819
rect 17144 18788 19441 18816
rect 15703 18720 15976 18748
rect 16393 18751 16451 18757
rect 15703 18717 15715 18720
rect 15657 18711 15715 18717
rect 16393 18717 16405 18751
rect 16439 18748 16451 18751
rect 16942 18748 16948 18760
rect 16439 18720 16948 18748
rect 16439 18717 16451 18720
rect 16393 18711 16451 18717
rect 10336 18652 12112 18680
rect 5537 18615 5595 18621
rect 5537 18581 5549 18615
rect 5583 18612 5595 18615
rect 5718 18612 5724 18624
rect 5583 18584 5724 18612
rect 5583 18581 5595 18584
rect 5537 18575 5595 18581
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 8386 18572 8392 18624
rect 8444 18612 8450 18624
rect 9306 18612 9312 18624
rect 8444 18584 9312 18612
rect 8444 18572 8450 18584
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 9493 18615 9551 18621
rect 9493 18581 9505 18615
rect 9539 18612 9551 18615
rect 9950 18612 9956 18624
rect 9539 18584 9956 18612
rect 9539 18581 9551 18584
rect 9493 18575 9551 18581
rect 9950 18572 9956 18584
rect 10008 18612 10014 18624
rect 10686 18612 10692 18624
rect 10008 18584 10692 18612
rect 10008 18572 10014 18584
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 12084 18612 12112 18652
rect 12158 18640 12164 18692
rect 12216 18680 12222 18692
rect 12314 18683 12372 18689
rect 12314 18680 12326 18683
rect 12216 18652 12326 18680
rect 12216 18640 12222 18652
rect 12314 18649 12326 18652
rect 12360 18649 12372 18683
rect 15470 18680 15476 18692
rect 12314 18643 12372 18649
rect 13096 18652 15476 18680
rect 13096 18612 13124 18652
rect 15470 18640 15476 18652
rect 15528 18640 15534 18692
rect 12084 18584 13124 18612
rect 13170 18572 13176 18624
rect 13228 18612 13234 18624
rect 15672 18612 15700 18711
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 17144 18757 17172 18788
rect 19429 18785 19441 18788
rect 19475 18785 19487 18819
rect 19429 18779 19487 18785
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 17865 18751 17923 18757
rect 17865 18717 17877 18751
rect 17911 18748 17923 18751
rect 18506 18748 18512 18760
rect 17911 18720 18512 18748
rect 17911 18717 17923 18720
rect 17865 18711 17923 18717
rect 18506 18708 18512 18720
rect 18564 18708 18570 18760
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18748 18659 18751
rect 19536 18748 19564 18856
rect 24670 18844 24676 18896
rect 24728 18844 24734 18896
rect 25961 18887 26019 18893
rect 25961 18853 25973 18887
rect 26007 18853 26019 18887
rect 25961 18847 26019 18853
rect 20346 18816 20352 18828
rect 19628 18788 20352 18816
rect 19628 18757 19656 18788
rect 20346 18776 20352 18788
rect 20404 18776 20410 18828
rect 21637 18819 21695 18825
rect 21637 18785 21649 18819
rect 21683 18816 21695 18819
rect 22646 18816 22652 18828
rect 21683 18788 22652 18816
rect 21683 18785 21695 18788
rect 21637 18779 21695 18785
rect 22646 18776 22652 18788
rect 22704 18776 22710 18828
rect 25976 18816 26004 18847
rect 22848 18788 26004 18816
rect 18647 18720 19564 18748
rect 19613 18751 19671 18757
rect 18647 18717 18659 18720
rect 18601 18711 18659 18717
rect 19613 18717 19625 18751
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 19889 18751 19947 18757
rect 19889 18717 19901 18751
rect 19935 18717 19947 18751
rect 19889 18711 19947 18717
rect 20073 18751 20131 18757
rect 20073 18717 20085 18751
rect 20119 18748 20131 18751
rect 20714 18748 20720 18760
rect 20119 18720 20720 18748
rect 20119 18717 20131 18720
rect 20073 18711 20131 18717
rect 19334 18640 19340 18692
rect 19392 18680 19398 18692
rect 19904 18680 19932 18711
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 21358 18708 21364 18760
rect 21416 18708 21422 18760
rect 22189 18751 22247 18757
rect 22189 18717 22201 18751
rect 22235 18748 22247 18751
rect 22848 18748 22876 18788
rect 22235 18720 22876 18748
rect 22925 18751 22983 18757
rect 22235 18717 22247 18720
rect 22189 18711 22247 18717
rect 22925 18717 22937 18751
rect 22971 18748 22983 18751
rect 23198 18748 23204 18760
rect 22971 18720 23204 18748
rect 22971 18717 22983 18720
rect 22925 18711 22983 18717
rect 23198 18708 23204 18720
rect 23256 18708 23262 18760
rect 23753 18751 23811 18757
rect 23753 18717 23765 18751
rect 23799 18748 23811 18751
rect 25682 18748 25688 18760
rect 23799 18720 25688 18748
rect 23799 18717 23811 18720
rect 23753 18711 23811 18717
rect 25682 18708 25688 18720
rect 25740 18708 25746 18760
rect 25777 18751 25835 18757
rect 25777 18717 25789 18751
rect 25823 18748 25835 18751
rect 26436 18748 26464 18924
rect 29178 18912 29184 18924
rect 29236 18912 29242 18964
rect 30469 18955 30527 18961
rect 30469 18921 30481 18955
rect 30515 18952 30527 18955
rect 30558 18952 30564 18964
rect 30515 18924 30564 18952
rect 30515 18921 30527 18924
rect 30469 18915 30527 18921
rect 30558 18912 30564 18924
rect 30616 18912 30622 18964
rect 36725 18955 36783 18961
rect 36725 18921 36737 18955
rect 36771 18952 36783 18955
rect 43714 18952 43720 18964
rect 36771 18924 43720 18952
rect 36771 18921 36783 18924
rect 36725 18915 36783 18921
rect 43714 18912 43720 18924
rect 43772 18912 43778 18964
rect 43898 18912 43904 18964
rect 43956 18952 43962 18964
rect 43993 18955 44051 18961
rect 43993 18952 44005 18955
rect 43956 18924 44005 18952
rect 43956 18912 43962 18924
rect 43993 18921 44005 18924
rect 44039 18921 44051 18955
rect 43993 18915 44051 18921
rect 45649 18955 45707 18961
rect 45649 18921 45661 18955
rect 45695 18952 45707 18955
rect 45738 18952 45744 18964
rect 45695 18924 45744 18952
rect 45695 18921 45707 18924
rect 45649 18915 45707 18921
rect 45738 18912 45744 18924
rect 45796 18912 45802 18964
rect 46290 18912 46296 18964
rect 46348 18952 46354 18964
rect 46661 18955 46719 18961
rect 46661 18952 46673 18955
rect 46348 18924 46673 18952
rect 46348 18912 46354 18924
rect 46661 18921 46673 18924
rect 46707 18921 46719 18955
rect 46661 18915 46719 18921
rect 48498 18912 48504 18964
rect 48556 18952 48562 18964
rect 50522 18952 50528 18964
rect 48556 18924 50528 18952
rect 48556 18912 48562 18924
rect 50522 18912 50528 18924
rect 50580 18912 50586 18964
rect 28905 18887 28963 18893
rect 28905 18853 28917 18887
rect 28951 18884 28963 18887
rect 54294 18884 54300 18896
rect 28951 18856 54300 18884
rect 28951 18853 28963 18856
rect 28905 18847 28963 18853
rect 54294 18844 54300 18856
rect 54352 18844 54358 18896
rect 26510 18776 26516 18828
rect 26568 18776 26574 18828
rect 27522 18776 27528 18828
rect 27580 18816 27586 18828
rect 29454 18816 29460 18828
rect 27580 18788 29460 18816
rect 27580 18776 27586 18788
rect 29454 18776 29460 18788
rect 29512 18776 29518 18828
rect 29730 18776 29736 18828
rect 29788 18816 29794 18828
rect 29788 18788 30696 18816
rect 29788 18776 29794 18788
rect 25823 18720 26464 18748
rect 25823 18717 25835 18720
rect 25777 18711 25835 18717
rect 27798 18708 27804 18760
rect 27856 18748 27862 18760
rect 28353 18751 28411 18757
rect 28353 18748 28365 18751
rect 27856 18720 28365 18748
rect 27856 18708 27862 18720
rect 28353 18717 28365 18720
rect 28399 18717 28411 18751
rect 28353 18711 28411 18717
rect 28442 18708 28448 18760
rect 28500 18748 28506 18760
rect 28810 18757 28816 18760
rect 28629 18751 28687 18757
rect 28629 18748 28641 18751
rect 28500 18720 28641 18748
rect 28500 18708 28506 18720
rect 28629 18717 28641 18720
rect 28675 18717 28687 18751
rect 28629 18711 28687 18717
rect 28773 18751 28816 18757
rect 28773 18717 28785 18751
rect 28773 18711 28816 18717
rect 28810 18708 28816 18711
rect 28868 18708 28874 18760
rect 30190 18708 30196 18760
rect 30248 18708 30254 18760
rect 30285 18751 30343 18757
rect 30285 18717 30297 18751
rect 30331 18717 30343 18751
rect 30285 18711 30343 18717
rect 19392 18652 19932 18680
rect 19392 18640 19398 18652
rect 20162 18640 20168 18692
rect 20220 18680 20226 18692
rect 20220 18652 23152 18680
rect 20220 18640 20226 18652
rect 13228 18584 15700 18612
rect 17313 18615 17371 18621
rect 13228 18572 13234 18584
rect 17313 18581 17325 18615
rect 17359 18612 17371 18615
rect 17954 18612 17960 18624
rect 17359 18584 17960 18612
rect 17359 18581 17371 18584
rect 17313 18575 17371 18581
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 19242 18572 19248 18624
rect 19300 18612 19306 18624
rect 21174 18612 21180 18624
rect 19300 18584 21180 18612
rect 19300 18572 19306 18584
rect 21174 18572 21180 18584
rect 21232 18612 21238 18624
rect 23124 18621 23152 18652
rect 21453 18615 21511 18621
rect 21453 18612 21465 18615
rect 21232 18584 21465 18612
rect 21232 18572 21238 18584
rect 21453 18581 21465 18584
rect 21499 18581 21511 18615
rect 21453 18575 21511 18581
rect 23109 18615 23167 18621
rect 23109 18581 23121 18615
rect 23155 18581 23167 18615
rect 23216 18612 23244 18708
rect 24946 18640 24952 18692
rect 25004 18640 25010 18692
rect 25222 18640 25228 18692
rect 25280 18680 25286 18692
rect 26780 18683 26838 18689
rect 25280 18652 25360 18680
rect 25280 18640 25286 18652
rect 23937 18615 23995 18621
rect 23937 18612 23949 18615
rect 23216 18584 23949 18612
rect 23109 18575 23167 18581
rect 23937 18581 23949 18584
rect 23983 18581 23995 18615
rect 23937 18575 23995 18581
rect 24854 18572 24860 18624
rect 24912 18612 24918 18624
rect 25133 18615 25191 18621
rect 25133 18612 25145 18615
rect 24912 18584 25145 18612
rect 24912 18572 24918 18584
rect 25133 18581 25145 18584
rect 25179 18581 25191 18615
rect 25332 18612 25360 18652
rect 26780 18649 26792 18683
rect 26826 18680 26838 18683
rect 27246 18680 27252 18692
rect 26826 18652 27252 18680
rect 26826 18649 26838 18652
rect 26780 18643 26838 18649
rect 27246 18640 27252 18652
rect 27304 18640 27310 18692
rect 27356 18652 28028 18680
rect 27356 18612 27384 18652
rect 25332 18584 27384 18612
rect 25133 18575 25191 18581
rect 27706 18572 27712 18624
rect 27764 18612 27770 18624
rect 27893 18615 27951 18621
rect 27893 18612 27905 18615
rect 27764 18584 27905 18612
rect 27764 18572 27770 18584
rect 27893 18581 27905 18584
rect 27939 18581 27951 18615
rect 28000 18612 28028 18652
rect 28534 18640 28540 18692
rect 28592 18640 28598 18692
rect 30006 18612 30012 18624
rect 28000 18584 30012 18612
rect 27893 18575 27951 18581
rect 30006 18572 30012 18584
rect 30064 18572 30070 18624
rect 30300 18612 30328 18711
rect 30668 18680 30696 18788
rect 30742 18776 30748 18828
rect 30800 18816 30806 18828
rect 30800 18788 31340 18816
rect 30800 18776 30806 18788
rect 31312 18757 31340 18788
rect 31386 18776 31392 18828
rect 31444 18776 31450 18828
rect 31478 18776 31484 18828
rect 31536 18776 31542 18828
rect 37366 18776 37372 18828
rect 37424 18776 37430 18828
rect 38749 18819 38807 18825
rect 38749 18785 38761 18819
rect 38795 18816 38807 18819
rect 40494 18816 40500 18828
rect 38795 18788 40500 18816
rect 38795 18785 38807 18788
rect 38749 18779 38807 18785
rect 40494 18776 40500 18788
rect 40552 18776 40558 18828
rect 41230 18776 41236 18828
rect 41288 18776 41294 18828
rect 49786 18816 49792 18828
rect 41386 18788 46152 18816
rect 31297 18751 31355 18757
rect 31297 18717 31309 18751
rect 31343 18748 31355 18751
rect 31662 18748 31668 18760
rect 31343 18720 31668 18748
rect 31343 18717 31355 18720
rect 31297 18711 31355 18717
rect 31662 18708 31668 18720
rect 31720 18708 31726 18760
rect 32398 18708 32404 18760
rect 32456 18708 32462 18760
rect 37090 18708 37096 18760
rect 37148 18708 37154 18760
rect 38838 18708 38844 18760
rect 38896 18748 38902 18760
rect 38933 18751 38991 18757
rect 38933 18748 38945 18751
rect 38896 18720 38945 18748
rect 38896 18708 38902 18720
rect 38933 18717 38945 18720
rect 38979 18717 38991 18751
rect 38933 18711 38991 18717
rect 40954 18708 40960 18760
rect 41012 18708 41018 18760
rect 30668 18652 31754 18680
rect 30929 18615 30987 18621
rect 30929 18612 30941 18615
rect 30300 18584 30941 18612
rect 30929 18581 30941 18584
rect 30975 18581 30987 18615
rect 31726 18612 31754 18652
rect 32950 18640 32956 18692
rect 33008 18680 33014 18692
rect 41386 18680 41414 18788
rect 42518 18708 42524 18760
rect 42576 18708 42582 18760
rect 42614 18751 42672 18757
rect 42614 18717 42626 18751
rect 42660 18717 42672 18751
rect 42614 18711 42672 18717
rect 33008 18652 41414 18680
rect 33008 18640 33014 18652
rect 32585 18615 32643 18621
rect 32585 18612 32597 18615
rect 31726 18584 32597 18612
rect 30929 18575 30987 18581
rect 32585 18581 32597 18584
rect 32631 18581 32643 18615
rect 32585 18575 32643 18581
rect 37090 18572 37096 18624
rect 37148 18612 37154 18624
rect 37185 18615 37243 18621
rect 37185 18612 37197 18615
rect 37148 18584 37197 18612
rect 37148 18572 37154 18584
rect 37185 18581 37197 18584
rect 37231 18581 37243 18615
rect 37185 18575 37243 18581
rect 39114 18572 39120 18624
rect 39172 18572 39178 18624
rect 40494 18572 40500 18624
rect 40552 18612 40558 18624
rect 40589 18615 40647 18621
rect 40589 18612 40601 18615
rect 40552 18584 40601 18612
rect 40552 18572 40558 18584
rect 40589 18581 40601 18584
rect 40635 18581 40647 18615
rect 40589 18575 40647 18581
rect 41049 18615 41107 18621
rect 41049 18581 41061 18615
rect 41095 18612 41107 18615
rect 41138 18612 41144 18624
rect 41095 18584 41144 18612
rect 41095 18581 41107 18584
rect 41049 18575 41107 18581
rect 41138 18572 41144 18584
rect 41196 18572 41202 18624
rect 42629 18612 42657 18711
rect 42702 18708 42708 18760
rect 42760 18748 42766 18760
rect 42986 18751 43044 18757
rect 42986 18748 42998 18751
rect 42760 18720 42998 18748
rect 42760 18708 42766 18720
rect 42986 18717 42998 18720
rect 43032 18717 43044 18751
rect 42986 18711 43044 18717
rect 43714 18708 43720 18760
rect 43772 18748 43778 18760
rect 43772 18720 43944 18748
rect 43772 18708 43778 18720
rect 42794 18640 42800 18692
rect 42852 18640 42858 18692
rect 42886 18640 42892 18692
rect 42944 18640 42950 18692
rect 43622 18640 43628 18692
rect 43680 18640 43686 18692
rect 43809 18683 43867 18689
rect 43809 18649 43821 18683
rect 43855 18649 43867 18683
rect 43916 18680 43944 18720
rect 45370 18708 45376 18760
rect 45428 18708 45434 18760
rect 45465 18751 45523 18757
rect 45465 18717 45477 18751
rect 45511 18748 45523 18751
rect 46014 18748 46020 18760
rect 45511 18720 46020 18748
rect 45511 18717 45523 18720
rect 45465 18711 45523 18717
rect 46014 18708 46020 18720
rect 46072 18708 46078 18760
rect 46124 18757 46152 18788
rect 46216 18788 49792 18816
rect 46109 18751 46167 18757
rect 46109 18717 46121 18751
rect 46155 18717 46167 18751
rect 46109 18711 46167 18717
rect 46216 18680 46244 18788
rect 49786 18776 49792 18788
rect 49844 18776 49850 18828
rect 55490 18776 55496 18828
rect 55548 18776 55554 18828
rect 46477 18751 46535 18757
rect 46477 18717 46489 18751
rect 46523 18748 46535 18751
rect 46566 18748 46572 18760
rect 46523 18720 46572 18748
rect 46523 18717 46535 18720
rect 46477 18711 46535 18717
rect 46566 18708 46572 18720
rect 46624 18708 46630 18760
rect 46658 18708 46664 18760
rect 46716 18748 46722 18760
rect 47213 18751 47271 18757
rect 47213 18748 47225 18751
rect 46716 18720 47225 18748
rect 46716 18708 46722 18720
rect 47213 18717 47225 18720
rect 47259 18717 47271 18751
rect 47213 18711 47271 18717
rect 48406 18708 48412 18760
rect 48464 18748 48470 18760
rect 48501 18751 48559 18757
rect 48501 18748 48513 18751
rect 48464 18720 48513 18748
rect 48464 18708 48470 18720
rect 48501 18717 48513 18720
rect 48547 18717 48559 18751
rect 48501 18711 48559 18717
rect 48682 18708 48688 18760
rect 48740 18708 48746 18760
rect 55674 18708 55680 18760
rect 55732 18708 55738 18760
rect 56965 18751 57023 18757
rect 56965 18717 56977 18751
rect 57011 18717 57023 18751
rect 56965 18711 57023 18717
rect 57977 18751 58035 18757
rect 57977 18717 57989 18751
rect 58023 18748 58035 18751
rect 58986 18748 58992 18760
rect 58023 18720 58992 18748
rect 58023 18717 58035 18720
rect 57977 18711 58035 18717
rect 43916 18652 46244 18680
rect 46293 18683 46351 18689
rect 43809 18643 43867 18649
rect 46293 18649 46305 18683
rect 46339 18649 46351 18683
rect 46293 18643 46351 18649
rect 46385 18683 46443 18689
rect 46385 18649 46397 18683
rect 46431 18680 46443 18683
rect 47578 18680 47584 18692
rect 46431 18652 47584 18680
rect 46431 18649 46443 18652
rect 46385 18643 46443 18649
rect 42702 18612 42708 18624
rect 42629 18584 42708 18612
rect 42702 18572 42708 18584
rect 42760 18572 42766 18624
rect 43162 18572 43168 18624
rect 43220 18572 43226 18624
rect 43438 18572 43444 18624
rect 43496 18612 43502 18624
rect 43824 18612 43852 18643
rect 43496 18584 43852 18612
rect 43496 18572 43502 18584
rect 46106 18572 46112 18624
rect 46164 18612 46170 18624
rect 46308 18612 46336 18643
rect 47578 18640 47584 18652
rect 47636 18640 47642 18692
rect 47762 18640 47768 18692
rect 47820 18680 47826 18692
rect 50062 18680 50068 18692
rect 47820 18652 50068 18680
rect 47820 18640 47826 18652
rect 50062 18640 50068 18652
rect 50120 18640 50126 18692
rect 52362 18640 52368 18692
rect 52420 18680 52426 18692
rect 56980 18680 57008 18711
rect 58986 18708 58992 18720
rect 59044 18708 59050 18760
rect 52420 18652 57008 18680
rect 57241 18683 57299 18689
rect 52420 18640 52426 18652
rect 57241 18649 57253 18683
rect 57287 18680 57299 18683
rect 57287 18652 59032 18680
rect 57287 18649 57299 18652
rect 57241 18643 57299 18649
rect 59004 18624 59032 18652
rect 46934 18612 46940 18624
rect 46164 18584 46940 18612
rect 46164 18572 46170 18584
rect 46934 18572 46940 18584
rect 46992 18572 46998 18624
rect 47489 18615 47547 18621
rect 47489 18581 47501 18615
rect 47535 18612 47547 18615
rect 47670 18612 47676 18624
rect 47535 18584 47676 18612
rect 47535 18581 47547 18584
rect 47489 18575 47547 18581
rect 47670 18572 47676 18584
rect 47728 18572 47734 18624
rect 48869 18615 48927 18621
rect 48869 18581 48881 18615
rect 48915 18612 48927 18615
rect 48958 18612 48964 18624
rect 48915 18584 48964 18612
rect 48915 18581 48927 18584
rect 48869 18575 48927 18581
rect 48958 18572 48964 18584
rect 49016 18572 49022 18624
rect 55861 18615 55919 18621
rect 55861 18581 55873 18615
rect 55907 18612 55919 18615
rect 56134 18612 56140 18624
rect 55907 18584 56140 18612
rect 55907 18581 55919 18584
rect 55861 18575 55919 18581
rect 56134 18572 56140 18584
rect 56192 18572 56198 18624
rect 58066 18572 58072 18624
rect 58124 18572 58130 18624
rect 58986 18572 58992 18624
rect 59044 18572 59050 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 8110 18368 8116 18420
rect 8168 18408 8174 18420
rect 8168 18380 9168 18408
rect 8168 18368 8174 18380
rect 6086 18300 6092 18352
rect 6144 18340 6150 18352
rect 9140 18340 9168 18380
rect 9858 18368 9864 18420
rect 9916 18408 9922 18420
rect 10505 18411 10563 18417
rect 10505 18408 10517 18411
rect 9916 18380 10517 18408
rect 9916 18368 9922 18380
rect 10505 18377 10517 18380
rect 10551 18377 10563 18411
rect 10505 18371 10563 18377
rect 12158 18368 12164 18420
rect 12216 18368 12222 18420
rect 14645 18411 14703 18417
rect 14645 18408 14657 18411
rect 12406 18380 14657 18408
rect 9950 18340 9956 18352
rect 6144 18312 8248 18340
rect 9140 18312 9956 18340
rect 6144 18300 6150 18312
rect 5718 18232 5724 18284
rect 5776 18232 5782 18284
rect 8220 18281 8248 18312
rect 9950 18300 9956 18312
rect 10008 18300 10014 18352
rect 10134 18300 10140 18352
rect 10192 18340 10198 18352
rect 12406 18340 12434 18380
rect 14645 18377 14657 18380
rect 14691 18377 14703 18411
rect 14645 18371 14703 18377
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 16209 18411 16267 18417
rect 16209 18408 16221 18411
rect 15528 18380 16221 18408
rect 15528 18368 15534 18380
rect 16209 18377 16221 18380
rect 16255 18377 16267 18411
rect 16209 18371 16267 18377
rect 16390 18368 16396 18420
rect 16448 18408 16454 18420
rect 18322 18408 18328 18420
rect 16448 18380 18328 18408
rect 16448 18368 16454 18380
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 18509 18411 18567 18417
rect 18509 18377 18521 18411
rect 18555 18408 18567 18411
rect 25590 18408 25596 18420
rect 18555 18380 25596 18408
rect 18555 18377 18567 18380
rect 18509 18371 18567 18377
rect 25590 18368 25596 18380
rect 25648 18368 25654 18420
rect 25682 18368 25688 18420
rect 25740 18408 25746 18420
rect 26513 18411 26571 18417
rect 26513 18408 26525 18411
rect 25740 18380 26525 18408
rect 25740 18368 25746 18380
rect 26513 18377 26525 18380
rect 26559 18377 26571 18411
rect 26513 18371 26571 18377
rect 27246 18368 27252 18420
rect 27304 18368 27310 18420
rect 27614 18368 27620 18420
rect 27672 18368 27678 18420
rect 29730 18368 29736 18420
rect 29788 18368 29794 18420
rect 43162 18408 43168 18420
rect 29840 18380 43168 18408
rect 10192 18312 12434 18340
rect 13081 18343 13139 18349
rect 10192 18300 10198 18312
rect 13081 18309 13093 18343
rect 13127 18340 13139 18343
rect 13354 18340 13360 18352
rect 13127 18312 13360 18340
rect 13127 18309 13139 18312
rect 13081 18303 13139 18309
rect 13354 18300 13360 18312
rect 13412 18300 13418 18352
rect 21542 18340 21548 18352
rect 14384 18312 20383 18340
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18272 6791 18275
rect 8205 18275 8263 18281
rect 6779 18244 8156 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18204 6883 18207
rect 6914 18204 6920 18216
rect 6871 18176 6920 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 7098 18164 7104 18216
rect 7156 18164 7162 18216
rect 8128 18204 8156 18244
rect 8205 18241 8217 18275
rect 8251 18241 8263 18275
rect 9674 18272 9680 18284
rect 8205 18235 8263 18241
rect 8312 18244 9680 18272
rect 8312 18204 8340 18244
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 10318 18232 10324 18284
rect 10376 18232 10382 18284
rect 11974 18232 11980 18284
rect 12032 18232 12038 18284
rect 12894 18232 12900 18284
rect 12952 18232 12958 18284
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18272 13047 18275
rect 13170 18272 13176 18284
rect 13035 18244 13176 18272
rect 13035 18241 13047 18244
rect 12989 18235 13047 18241
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 13262 18232 13268 18284
rect 13320 18232 13326 18284
rect 8128 18176 8340 18204
rect 8478 18164 8484 18216
rect 8536 18164 8542 18216
rect 9306 18164 9312 18216
rect 9364 18204 9370 18216
rect 14384 18204 14412 18312
rect 14458 18232 14464 18284
rect 14516 18232 14522 18284
rect 16040 18281 16068 18312
rect 15289 18275 15347 18281
rect 15289 18241 15301 18275
rect 15335 18241 15347 18275
rect 15289 18235 15347 18241
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18241 16083 18275
rect 16025 18235 16083 18241
rect 9364 18176 14412 18204
rect 15304 18204 15332 18235
rect 17034 18232 17040 18284
rect 17092 18272 17098 18284
rect 17129 18275 17187 18281
rect 17129 18272 17141 18275
rect 17092 18244 17141 18272
rect 17092 18232 17098 18244
rect 17129 18241 17141 18244
rect 17175 18241 17187 18275
rect 17129 18235 17187 18241
rect 17396 18275 17454 18281
rect 17396 18241 17408 18275
rect 17442 18272 17454 18275
rect 17954 18272 17960 18284
rect 17442 18244 17960 18272
rect 17442 18241 17454 18244
rect 17396 18235 17454 18241
rect 17954 18232 17960 18244
rect 18012 18232 18018 18284
rect 19518 18232 19524 18284
rect 19576 18232 19582 18284
rect 16758 18204 16764 18216
rect 15304 18176 16764 18204
rect 9364 18164 9370 18176
rect 16758 18164 16764 18176
rect 16816 18164 16822 18216
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18204 19395 18207
rect 19610 18204 19616 18216
rect 19383 18176 19616 18204
rect 19383 18173 19395 18176
rect 19337 18167 19395 18173
rect 19610 18164 19616 18176
rect 19668 18204 19674 18216
rect 20162 18204 20168 18216
rect 19668 18176 20168 18204
rect 19668 18164 19674 18176
rect 20162 18164 20168 18176
rect 20220 18164 20226 18216
rect 20355 18204 20383 18312
rect 20456 18312 21548 18340
rect 20456 18281 20484 18312
rect 21542 18300 21548 18312
rect 21600 18300 21606 18352
rect 29748 18340 29776 18368
rect 24320 18312 29776 18340
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 20714 18272 20720 18284
rect 20441 18235 20499 18241
rect 20548 18244 20720 18272
rect 20548 18204 20576 18244
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 21177 18275 21235 18281
rect 21177 18241 21189 18275
rect 21223 18241 21235 18275
rect 21177 18235 21235 18241
rect 21192 18204 21220 18235
rect 21634 18232 21640 18284
rect 21692 18272 21698 18284
rect 22005 18275 22063 18281
rect 22005 18272 22017 18275
rect 21692 18244 22017 18272
rect 21692 18232 21698 18244
rect 22005 18241 22017 18244
rect 22051 18241 22063 18275
rect 22005 18235 22063 18241
rect 22094 18232 22100 18284
rect 22152 18272 22158 18284
rect 23109 18275 23167 18281
rect 23109 18272 23121 18275
rect 22152 18244 23121 18272
rect 22152 18232 22158 18244
rect 23109 18241 23121 18244
rect 23155 18241 23167 18275
rect 23109 18235 23167 18241
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18272 23351 18275
rect 24210 18272 24216 18284
rect 23339 18244 24216 18272
rect 23339 18241 23351 18244
rect 23293 18235 23351 18241
rect 24210 18232 24216 18244
rect 24268 18232 24274 18284
rect 24320 18281 24348 18312
rect 24305 18275 24363 18281
rect 24305 18241 24317 18275
rect 24351 18241 24363 18275
rect 24305 18235 24363 18241
rect 25590 18232 25596 18284
rect 25648 18272 25654 18284
rect 26329 18275 26387 18281
rect 26329 18272 26341 18275
rect 25648 18244 26341 18272
rect 25648 18232 25654 18244
rect 26329 18241 26341 18244
rect 26375 18272 26387 18275
rect 28074 18272 28080 18284
rect 26375 18244 28080 18272
rect 26375 18241 26387 18244
rect 26329 18235 26387 18241
rect 28074 18232 28080 18244
rect 28132 18232 28138 18284
rect 29454 18232 29460 18284
rect 29512 18232 29518 18284
rect 29546 18232 29552 18284
rect 29604 18232 29610 18284
rect 29730 18232 29736 18284
rect 29788 18232 29794 18284
rect 29840 18281 29868 18380
rect 43162 18368 43168 18380
rect 43220 18368 43226 18420
rect 46014 18368 46020 18420
rect 46072 18408 46078 18420
rect 46477 18411 46535 18417
rect 46477 18408 46489 18411
rect 46072 18380 46489 18408
rect 46072 18368 46078 18380
rect 46477 18377 46489 18380
rect 46523 18377 46535 18411
rect 46477 18371 46535 18377
rect 48314 18368 48320 18420
rect 48372 18408 48378 18420
rect 48372 18380 48728 18408
rect 48372 18368 48378 18380
rect 30837 18343 30895 18349
rect 30837 18340 30849 18343
rect 29932 18312 30849 18340
rect 29825 18275 29883 18281
rect 29825 18241 29837 18275
rect 29871 18241 29883 18275
rect 29825 18235 29883 18241
rect 21910 18204 21916 18216
rect 20355 18176 20576 18204
rect 20640 18176 20852 18204
rect 21192 18176 21916 18204
rect 9769 18139 9827 18145
rect 9769 18105 9781 18139
rect 9815 18136 9827 18139
rect 12618 18136 12624 18148
rect 9815 18108 12624 18136
rect 9815 18105 9827 18108
rect 9769 18099 9827 18105
rect 12618 18096 12624 18108
rect 12676 18096 12682 18148
rect 12713 18139 12771 18145
rect 12713 18105 12725 18139
rect 12759 18136 12771 18139
rect 14090 18136 14096 18148
rect 12759 18108 14096 18136
rect 12759 18105 12771 18108
rect 12713 18099 12771 18105
rect 14090 18096 14096 18108
rect 14148 18096 14154 18148
rect 14550 18096 14556 18148
rect 14608 18136 14614 18148
rect 14608 18108 17172 18136
rect 14608 18096 14614 18108
rect 5905 18071 5963 18077
rect 5905 18037 5917 18071
rect 5951 18068 5963 18071
rect 6546 18068 6552 18080
rect 5951 18040 6552 18068
rect 5951 18037 5963 18040
rect 5905 18031 5963 18037
rect 6546 18028 6552 18040
rect 6604 18028 6610 18080
rect 9582 18028 9588 18080
rect 9640 18068 9646 18080
rect 14458 18068 14464 18080
rect 9640 18040 14464 18068
rect 9640 18028 9646 18040
rect 14458 18028 14464 18040
rect 14516 18028 14522 18080
rect 15286 18028 15292 18080
rect 15344 18068 15350 18080
rect 15473 18071 15531 18077
rect 15473 18068 15485 18071
rect 15344 18040 15485 18068
rect 15344 18028 15350 18040
rect 15473 18037 15485 18040
rect 15519 18037 15531 18071
rect 17144 18068 17172 18108
rect 18506 18096 18512 18148
rect 18564 18136 18570 18148
rect 20640 18136 20668 18176
rect 18564 18108 20668 18136
rect 20824 18136 20852 18176
rect 21910 18164 21916 18176
rect 21968 18164 21974 18216
rect 26142 18164 26148 18216
rect 26200 18204 26206 18216
rect 27706 18204 27712 18216
rect 26200 18176 27712 18204
rect 26200 18164 26206 18176
rect 27706 18164 27712 18176
rect 27764 18164 27770 18216
rect 27893 18207 27951 18213
rect 27893 18173 27905 18207
rect 27939 18173 27951 18207
rect 27893 18167 27951 18173
rect 22189 18139 22247 18145
rect 22189 18136 22201 18139
rect 20824 18108 22201 18136
rect 18564 18096 18570 18108
rect 22189 18105 22201 18108
rect 22235 18105 22247 18139
rect 22189 18099 22247 18105
rect 23477 18139 23535 18145
rect 23477 18105 23489 18139
rect 23523 18136 23535 18139
rect 24302 18136 24308 18148
rect 23523 18108 24308 18136
rect 23523 18105 23535 18108
rect 23477 18099 23535 18105
rect 24302 18096 24308 18108
rect 24360 18096 24366 18148
rect 24486 18096 24492 18148
rect 24544 18096 24550 18148
rect 25130 18096 25136 18148
rect 25188 18136 25194 18148
rect 25958 18136 25964 18148
rect 25188 18108 25964 18136
rect 25188 18096 25194 18108
rect 25958 18096 25964 18108
rect 26016 18096 26022 18148
rect 19242 18068 19248 18080
rect 17144 18040 19248 18068
rect 15473 18031 15531 18037
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 19334 18028 19340 18080
rect 19392 18068 19398 18080
rect 19705 18071 19763 18077
rect 19705 18068 19717 18071
rect 19392 18040 19717 18068
rect 19392 18028 19398 18040
rect 19705 18037 19717 18040
rect 19751 18037 19763 18071
rect 19705 18031 19763 18037
rect 20254 18028 20260 18080
rect 20312 18068 20318 18080
rect 20625 18071 20683 18077
rect 20625 18068 20637 18071
rect 20312 18040 20637 18068
rect 20312 18028 20318 18040
rect 20625 18037 20637 18040
rect 20671 18037 20683 18071
rect 20625 18031 20683 18037
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 21361 18071 21419 18077
rect 21361 18068 21373 18071
rect 20772 18040 21373 18068
rect 20772 18028 20778 18040
rect 21361 18037 21373 18040
rect 21407 18037 21419 18071
rect 21361 18031 21419 18037
rect 22646 18028 22652 18080
rect 22704 18068 22710 18080
rect 27706 18068 27712 18080
rect 22704 18040 27712 18068
rect 22704 18028 22710 18040
rect 27706 18028 27712 18040
rect 27764 18068 27770 18080
rect 27908 18068 27936 18167
rect 29932 18136 29960 18312
rect 30837 18309 30849 18312
rect 30883 18309 30895 18343
rect 30837 18303 30895 18309
rect 30929 18343 30987 18349
rect 30929 18309 30941 18343
rect 30975 18340 30987 18343
rect 32214 18340 32220 18352
rect 30975 18312 32220 18340
rect 30975 18309 30987 18312
rect 30929 18303 30987 18309
rect 30006 18232 30012 18284
rect 30064 18272 30070 18284
rect 30944 18272 30972 18303
rect 32214 18300 32220 18312
rect 32272 18300 32278 18352
rect 32398 18300 32404 18352
rect 32456 18340 32462 18352
rect 32456 18312 34008 18340
rect 32456 18300 32462 18312
rect 32950 18272 32956 18284
rect 30064 18244 30972 18272
rect 32324 18244 32956 18272
rect 30064 18232 30070 18244
rect 30742 18164 30748 18216
rect 30800 18164 30806 18216
rect 32324 18213 32352 18244
rect 32950 18232 32956 18244
rect 33008 18232 33014 18284
rect 33980 18272 34008 18312
rect 34054 18300 34060 18352
rect 34112 18340 34118 18352
rect 34333 18343 34391 18349
rect 34333 18340 34345 18343
rect 34112 18312 34345 18340
rect 34112 18300 34118 18312
rect 34333 18309 34345 18312
rect 34379 18309 34391 18343
rect 34333 18303 34391 18309
rect 41230 18300 41236 18352
rect 41288 18340 41294 18352
rect 41506 18340 41512 18352
rect 41288 18312 41512 18340
rect 41288 18300 41294 18312
rect 41506 18300 41512 18312
rect 41564 18300 41570 18352
rect 42797 18343 42855 18349
rect 42797 18309 42809 18343
rect 42843 18309 42855 18343
rect 42797 18303 42855 18309
rect 38654 18272 38660 18284
rect 33980 18244 38660 18272
rect 38654 18232 38660 18244
rect 38712 18272 38718 18284
rect 38712 18244 38976 18272
rect 38712 18232 38718 18244
rect 32309 18207 32367 18213
rect 32309 18173 32321 18207
rect 32355 18173 32367 18207
rect 32309 18167 32367 18173
rect 32398 18164 32404 18216
rect 32456 18204 32462 18216
rect 32493 18207 32551 18213
rect 32493 18204 32505 18207
rect 32456 18176 32505 18204
rect 32456 18164 32462 18176
rect 32493 18173 32505 18176
rect 32539 18173 32551 18207
rect 32493 18167 32551 18173
rect 32582 18164 32588 18216
rect 32640 18164 32646 18216
rect 32674 18164 32680 18216
rect 32732 18164 32738 18216
rect 32766 18164 32772 18216
rect 32824 18164 32830 18216
rect 33870 18164 33876 18216
rect 33928 18204 33934 18216
rect 34425 18207 34483 18213
rect 34425 18204 34437 18207
rect 33928 18176 34437 18204
rect 33928 18164 33934 18176
rect 34425 18173 34437 18176
rect 34471 18173 34483 18207
rect 34425 18167 34483 18173
rect 34609 18207 34667 18213
rect 34609 18173 34621 18207
rect 34655 18204 34667 18207
rect 35342 18204 35348 18216
rect 34655 18176 35348 18204
rect 34655 18173 34667 18176
rect 34609 18167 34667 18173
rect 35342 18164 35348 18176
rect 35400 18164 35406 18216
rect 38838 18164 38844 18216
rect 38896 18164 38902 18216
rect 38948 18204 38976 18244
rect 39114 18232 39120 18284
rect 39172 18232 39178 18284
rect 42426 18232 42432 18284
rect 42484 18272 42490 18284
rect 42613 18275 42671 18281
rect 42613 18272 42625 18275
rect 42484 18244 42625 18272
rect 42484 18232 42490 18244
rect 42613 18241 42625 18244
rect 42659 18241 42671 18275
rect 42613 18235 42671 18241
rect 40221 18207 40279 18213
rect 40221 18204 40233 18207
rect 38948 18176 40233 18204
rect 40221 18173 40233 18176
rect 40267 18204 40279 18207
rect 40954 18204 40960 18216
rect 40267 18176 40960 18204
rect 40267 18173 40279 18176
rect 40221 18167 40279 18173
rect 40954 18164 40960 18176
rect 41012 18164 41018 18216
rect 42812 18204 42840 18303
rect 42886 18300 42892 18352
rect 42944 18300 42950 18352
rect 43622 18300 43628 18352
rect 43680 18340 43686 18352
rect 44726 18340 44732 18352
rect 43680 18312 44732 18340
rect 43680 18300 43686 18312
rect 44726 18300 44732 18312
rect 44784 18300 44790 18352
rect 46106 18300 46112 18352
rect 46164 18300 46170 18352
rect 46201 18343 46259 18349
rect 46201 18309 46213 18343
rect 46247 18340 46259 18343
rect 46842 18340 46848 18352
rect 46247 18312 46848 18340
rect 46247 18309 46259 18312
rect 46201 18303 46259 18309
rect 46842 18300 46848 18312
rect 46900 18300 46906 18352
rect 42978 18232 42984 18284
rect 43036 18232 43042 18284
rect 44174 18232 44180 18284
rect 44232 18272 44238 18284
rect 45925 18275 45983 18281
rect 45925 18272 45937 18275
rect 44232 18244 45937 18272
rect 44232 18232 44238 18244
rect 45925 18241 45937 18244
rect 45971 18241 45983 18275
rect 45925 18235 45983 18241
rect 46293 18275 46351 18281
rect 46293 18241 46305 18275
rect 46339 18241 46351 18275
rect 46293 18235 46351 18241
rect 42886 18204 42892 18216
rect 42812 18176 42892 18204
rect 42886 18164 42892 18176
rect 42944 18164 42950 18216
rect 46308 18204 46336 18235
rect 47118 18232 47124 18284
rect 47176 18272 47182 18284
rect 48498 18272 48504 18284
rect 47176 18244 48504 18272
rect 47176 18232 47182 18244
rect 48498 18232 48504 18244
rect 48556 18232 48562 18284
rect 48700 18272 48728 18380
rect 49970 18368 49976 18420
rect 50028 18408 50034 18420
rect 50065 18411 50123 18417
rect 50065 18408 50077 18411
rect 50028 18380 50077 18408
rect 50028 18368 50034 18380
rect 50065 18377 50077 18380
rect 50111 18377 50123 18411
rect 50065 18371 50123 18377
rect 55125 18411 55183 18417
rect 55125 18377 55137 18411
rect 55171 18408 55183 18411
rect 55674 18408 55680 18420
rect 55171 18380 55680 18408
rect 55171 18377 55183 18380
rect 55125 18371 55183 18377
rect 55674 18368 55680 18380
rect 55732 18368 55738 18420
rect 57238 18408 57244 18420
rect 55968 18380 57244 18408
rect 54849 18343 54907 18349
rect 54849 18309 54861 18343
rect 54895 18340 54907 18343
rect 55968 18340 55996 18380
rect 57238 18368 57244 18380
rect 57296 18368 57302 18420
rect 58710 18368 58716 18420
rect 58768 18368 58774 18420
rect 56134 18349 56140 18352
rect 56128 18340 56140 18349
rect 54895 18312 55996 18340
rect 56095 18312 56140 18340
rect 54895 18309 54907 18312
rect 54849 18303 54907 18309
rect 56128 18303 56140 18312
rect 56134 18300 56140 18303
rect 56192 18300 56198 18352
rect 48958 18281 48964 18284
rect 48952 18272 48964 18281
rect 48700 18244 48820 18272
rect 48919 18244 48964 18272
rect 46566 18204 46572 18216
rect 46308 18176 46572 18204
rect 46566 18164 46572 18176
rect 46624 18204 46630 18216
rect 48130 18204 48136 18216
rect 46624 18176 48136 18204
rect 46624 18164 46630 18176
rect 48130 18164 48136 18176
rect 48188 18164 48194 18216
rect 48685 18207 48743 18213
rect 48685 18173 48697 18207
rect 48731 18204 48743 18207
rect 48792 18204 48820 18244
rect 48952 18235 48964 18244
rect 48958 18232 48964 18235
rect 49016 18232 49022 18284
rect 54570 18232 54576 18284
rect 54628 18232 54634 18284
rect 54754 18232 54760 18284
rect 54812 18232 54818 18284
rect 54938 18232 54944 18284
rect 54996 18232 55002 18284
rect 48731 18176 48820 18204
rect 48731 18173 48743 18176
rect 48685 18167 48743 18173
rect 55858 18164 55864 18216
rect 55916 18164 55922 18216
rect 58728 18148 58756 18368
rect 29288 18108 29960 18136
rect 30377 18139 30435 18145
rect 27764 18040 27936 18068
rect 27764 18028 27770 18040
rect 28074 18028 28080 18080
rect 28132 18068 28138 18080
rect 29288 18077 29316 18108
rect 30377 18105 30389 18139
rect 30423 18136 30435 18139
rect 43165 18139 43223 18145
rect 30423 18108 36584 18136
rect 30423 18105 30435 18108
rect 30377 18099 30435 18105
rect 29273 18071 29331 18077
rect 29273 18068 29285 18071
rect 28132 18040 29285 18068
rect 28132 18028 28138 18040
rect 29273 18037 29285 18040
rect 29319 18037 29331 18071
rect 29273 18031 29331 18037
rect 32214 18028 32220 18080
rect 32272 18068 32278 18080
rect 32674 18068 32680 18080
rect 32272 18040 32680 18068
rect 32272 18028 32278 18040
rect 32674 18028 32680 18040
rect 32732 18028 32738 18080
rect 33962 18028 33968 18080
rect 34020 18028 34026 18080
rect 36556 18068 36584 18108
rect 43165 18105 43177 18139
rect 43211 18105 43223 18139
rect 43165 18099 43223 18105
rect 42426 18068 42432 18080
rect 36556 18040 42432 18068
rect 42426 18028 42432 18040
rect 42484 18028 42490 18080
rect 42518 18028 42524 18080
rect 42576 18068 42582 18080
rect 43180 18068 43208 18099
rect 58710 18096 58716 18148
rect 58768 18096 58774 18148
rect 42576 18040 43208 18068
rect 42576 18028 42582 18040
rect 43438 18028 43444 18080
rect 43496 18068 43502 18080
rect 52086 18068 52092 18080
rect 43496 18040 52092 18068
rect 43496 18028 43502 18040
rect 52086 18028 52092 18040
rect 52144 18028 52150 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 5258 17824 5264 17876
rect 5316 17864 5322 17876
rect 9953 17867 10011 17873
rect 5316 17836 8892 17864
rect 5316 17824 5322 17836
rect 8864 17796 8892 17836
rect 9953 17833 9965 17867
rect 9999 17864 10011 17867
rect 10226 17864 10232 17876
rect 9999 17836 10232 17864
rect 9999 17833 10011 17836
rect 9953 17827 10011 17833
rect 10226 17824 10232 17836
rect 10284 17824 10290 17876
rect 10318 17824 10324 17876
rect 10376 17864 10382 17876
rect 13262 17864 13268 17876
rect 10376 17836 13268 17864
rect 10376 17824 10382 17836
rect 13262 17824 13268 17836
rect 13320 17824 13326 17876
rect 14274 17824 14280 17876
rect 14332 17864 14338 17876
rect 14461 17867 14519 17873
rect 14461 17864 14473 17867
rect 14332 17836 14473 17864
rect 14332 17824 14338 17836
rect 14461 17833 14473 17836
rect 14507 17833 14519 17867
rect 14461 17827 14519 17833
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 15289 17867 15347 17873
rect 15289 17864 15301 17867
rect 15252 17836 15301 17864
rect 15252 17824 15258 17836
rect 15289 17833 15301 17836
rect 15335 17833 15347 17867
rect 15289 17827 15347 17833
rect 16758 17824 16764 17876
rect 16816 17824 16822 17876
rect 16942 17824 16948 17876
rect 17000 17864 17006 17876
rect 18601 17867 18659 17873
rect 18601 17864 18613 17867
rect 17000 17836 18613 17864
rect 17000 17824 17006 17836
rect 18601 17833 18613 17836
rect 18647 17833 18659 17867
rect 18601 17827 18659 17833
rect 18690 17824 18696 17876
rect 18748 17864 18754 17876
rect 24486 17864 24492 17876
rect 18748 17836 24492 17864
rect 18748 17824 18754 17836
rect 24486 17824 24492 17836
rect 24544 17824 24550 17876
rect 24946 17824 24952 17876
rect 25004 17864 25010 17876
rect 32033 17867 32091 17873
rect 25004 17836 31754 17864
rect 25004 17824 25010 17836
rect 23658 17796 23664 17808
rect 8864 17768 23664 17796
rect 23658 17756 23664 17768
rect 23716 17756 23722 17808
rect 28534 17796 28540 17808
rect 23860 17768 28540 17796
rect 934 17688 940 17740
rect 992 17728 998 17740
rect 1765 17731 1823 17737
rect 1765 17728 1777 17731
rect 992 17700 1777 17728
rect 992 17688 998 17700
rect 1765 17697 1777 17700
rect 1811 17697 1823 17731
rect 1765 17691 1823 17697
rect 8110 17688 8116 17740
rect 8168 17688 8174 17740
rect 8573 17731 8631 17737
rect 8573 17697 8585 17731
rect 8619 17697 8631 17731
rect 9950 17728 9956 17740
rect 8573 17691 8631 17697
rect 9876 17700 9956 17728
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17660 1639 17663
rect 6454 17660 6460 17672
rect 1627 17632 6460 17660
rect 1627 17629 1639 17632
rect 1581 17623 1639 17629
rect 6454 17620 6460 17632
rect 6512 17620 6518 17672
rect 6546 17620 6552 17672
rect 6604 17620 6610 17672
rect 8205 17663 8263 17669
rect 8205 17629 8217 17663
rect 8251 17629 8263 17663
rect 8588 17660 8616 17691
rect 9876 17669 9904 17700
rect 9950 17688 9956 17700
rect 10008 17728 10014 17740
rect 10318 17728 10324 17740
rect 10008 17700 10324 17728
rect 10008 17688 10014 17700
rect 10318 17688 10324 17700
rect 10376 17688 10382 17740
rect 18690 17728 18696 17740
rect 12406 17700 18696 17728
rect 9125 17663 9183 17669
rect 9125 17660 9137 17663
rect 8588 17632 9137 17660
rect 8205 17623 8263 17629
rect 9125 17629 9137 17632
rect 9171 17629 9183 17663
rect 9125 17623 9183 17629
rect 9861 17663 9919 17669
rect 9861 17629 9873 17663
rect 9907 17629 9919 17663
rect 9861 17623 9919 17629
rect 8220 17592 8248 17623
rect 10042 17620 10048 17672
rect 10100 17660 10106 17672
rect 12406 17660 12434 17700
rect 10100 17632 12434 17660
rect 14277 17663 14335 17669
rect 10100 17620 10106 17632
rect 14277 17629 14289 17663
rect 14323 17660 14335 17663
rect 14826 17660 14832 17672
rect 14323 17632 14832 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 15102 17620 15108 17672
rect 15160 17620 15166 17672
rect 15856 17669 15884 17700
rect 18690 17688 18696 17700
rect 18748 17688 18754 17740
rect 18782 17688 18788 17740
rect 18840 17728 18846 17740
rect 19521 17731 19579 17737
rect 19521 17728 19533 17731
rect 18840 17700 19533 17728
rect 18840 17688 18846 17700
rect 19521 17697 19533 17700
rect 19567 17697 19579 17731
rect 23290 17728 23296 17740
rect 19521 17691 19579 17697
rect 20088 17700 23296 17728
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 16206 17620 16212 17672
rect 16264 17660 16270 17672
rect 16577 17663 16635 17669
rect 16577 17660 16589 17663
rect 16264 17632 16589 17660
rect 16264 17620 16270 17632
rect 16577 17629 16589 17632
rect 16623 17629 16635 17663
rect 16577 17623 16635 17629
rect 17681 17663 17739 17669
rect 17681 17629 17693 17663
rect 17727 17660 17739 17663
rect 17727 17632 18000 17660
rect 17727 17629 17739 17632
rect 17681 17623 17739 17629
rect 8220 17564 16068 17592
rect 6730 17484 6736 17536
rect 6788 17484 6794 17536
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 16040 17533 16068 17564
rect 9309 17527 9367 17533
rect 9309 17524 9321 17527
rect 8628 17496 9321 17524
rect 8628 17484 8634 17496
rect 9309 17493 9321 17496
rect 9355 17493 9367 17527
rect 9309 17487 9367 17493
rect 16025 17527 16083 17533
rect 16025 17493 16037 17527
rect 16071 17493 16083 17527
rect 16025 17487 16083 17493
rect 17770 17484 17776 17536
rect 17828 17524 17834 17536
rect 17865 17527 17923 17533
rect 17865 17524 17877 17527
rect 17828 17496 17877 17524
rect 17828 17484 17834 17496
rect 17865 17493 17877 17496
rect 17911 17493 17923 17527
rect 17972 17524 18000 17632
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 18417 17663 18475 17669
rect 18417 17660 18429 17663
rect 18104 17632 18429 17660
rect 18104 17620 18110 17632
rect 18417 17629 18429 17632
rect 18463 17629 18475 17663
rect 18417 17623 18475 17629
rect 19426 17620 19432 17672
rect 19484 17620 19490 17672
rect 19610 17620 19616 17672
rect 19668 17620 19674 17672
rect 20088 17669 20116 17700
rect 23290 17688 23296 17700
rect 23348 17688 23354 17740
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17629 20131 17663
rect 20073 17623 20131 17629
rect 20898 17620 20904 17672
rect 20956 17620 20962 17672
rect 20990 17620 20996 17672
rect 21048 17620 21054 17672
rect 23860 17660 23888 17768
rect 28534 17756 28540 17768
rect 28592 17796 28598 17808
rect 28592 17768 28672 17796
rect 28592 17756 28598 17768
rect 24210 17688 24216 17740
rect 24268 17728 24274 17740
rect 24268 17700 25268 17728
rect 24268 17688 24274 17700
rect 21091 17632 23888 17660
rect 18138 17552 18144 17604
rect 18196 17592 18202 17604
rect 18196 17564 20300 17592
rect 18196 17552 18202 17564
rect 18690 17524 18696 17536
rect 17972 17496 18696 17524
rect 17865 17487 17923 17493
rect 18690 17484 18696 17496
rect 18748 17484 18754 17536
rect 20272 17533 20300 17564
rect 20438 17552 20444 17604
rect 20496 17592 20502 17604
rect 21091 17592 21119 17632
rect 23934 17620 23940 17672
rect 23992 17660 23998 17672
rect 24765 17663 24823 17669
rect 24765 17660 24777 17663
rect 23992 17632 24777 17660
rect 23992 17620 23998 17632
rect 24765 17629 24777 17632
rect 24811 17629 24823 17663
rect 25133 17663 25191 17669
rect 25133 17660 25145 17663
rect 24765 17623 24823 17629
rect 24863 17632 25145 17660
rect 20496 17564 21119 17592
rect 20496 17552 20502 17564
rect 21542 17552 21548 17604
rect 21600 17592 21606 17604
rect 23952 17592 23980 17620
rect 21600 17564 23980 17592
rect 21600 17552 21606 17564
rect 24302 17552 24308 17604
rect 24360 17592 24366 17604
rect 24863 17592 24891 17632
rect 25133 17629 25145 17632
rect 25179 17629 25191 17663
rect 25240 17660 25268 17700
rect 25590 17688 25596 17740
rect 25648 17688 25654 17740
rect 25792 17700 27568 17728
rect 25792 17669 25820 17700
rect 25777 17663 25835 17669
rect 25777 17660 25789 17663
rect 25240 17632 25789 17660
rect 25133 17623 25191 17629
rect 25777 17629 25789 17632
rect 25823 17629 25835 17663
rect 25777 17623 25835 17629
rect 27062 17620 27068 17672
rect 27120 17620 27126 17672
rect 27338 17620 27344 17672
rect 27396 17620 27402 17672
rect 27433 17663 27491 17669
rect 27433 17629 27445 17663
rect 27479 17629 27491 17663
rect 27540 17660 27568 17700
rect 27890 17688 27896 17740
rect 27948 17728 27954 17740
rect 27948 17700 28580 17728
rect 27948 17688 27954 17700
rect 27982 17660 27988 17672
rect 27540 17632 27988 17660
rect 27433 17623 27491 17629
rect 24360 17564 24891 17592
rect 24360 17552 24366 17564
rect 25038 17552 25044 17604
rect 25096 17592 25102 17604
rect 27249 17595 27307 17601
rect 27249 17592 27261 17595
rect 25096 17564 27261 17592
rect 25096 17552 25102 17564
rect 27249 17561 27261 17564
rect 27295 17561 27307 17595
rect 27249 17555 27307 17561
rect 20257 17527 20315 17533
rect 20257 17493 20269 17527
rect 20303 17493 20315 17527
rect 20257 17487 20315 17493
rect 21082 17484 21088 17536
rect 21140 17524 21146 17536
rect 21177 17527 21235 17533
rect 21177 17524 21189 17527
rect 21140 17496 21189 17524
rect 21140 17484 21146 17496
rect 21177 17493 21189 17496
rect 21223 17493 21235 17527
rect 21177 17487 21235 17493
rect 24670 17484 24676 17536
rect 24728 17484 24734 17536
rect 24854 17484 24860 17536
rect 24912 17484 24918 17536
rect 24949 17527 25007 17533
rect 24949 17493 24961 17527
rect 24995 17524 25007 17527
rect 25222 17524 25228 17536
rect 24995 17496 25228 17524
rect 24995 17493 25007 17496
rect 24949 17487 25007 17493
rect 25222 17484 25228 17496
rect 25280 17484 25286 17536
rect 25406 17484 25412 17536
rect 25464 17524 25470 17536
rect 25961 17527 26019 17533
rect 25961 17524 25973 17527
rect 25464 17496 25973 17524
rect 25464 17484 25470 17496
rect 25961 17493 25973 17496
rect 26007 17493 26019 17527
rect 25961 17487 26019 17493
rect 27154 17484 27160 17536
rect 27212 17524 27218 17536
rect 27338 17524 27344 17536
rect 27212 17496 27344 17524
rect 27212 17484 27218 17496
rect 27338 17484 27344 17496
rect 27396 17524 27402 17536
rect 27448 17524 27476 17623
rect 27982 17620 27988 17632
rect 28040 17620 28046 17672
rect 28350 17669 28356 17672
rect 28169 17663 28227 17669
rect 28169 17629 28181 17663
rect 28215 17629 28227 17663
rect 28169 17623 28227 17629
rect 28317 17663 28356 17669
rect 28317 17629 28329 17663
rect 28317 17623 28356 17629
rect 27396 17496 27476 17524
rect 27617 17527 27675 17533
rect 27396 17484 27402 17496
rect 27617 17493 27629 17527
rect 27663 17524 27675 17527
rect 28184 17524 28212 17623
rect 28350 17620 28356 17623
rect 28408 17620 28414 17672
rect 28552 17669 28580 17700
rect 28644 17669 28672 17768
rect 29822 17756 29828 17808
rect 29880 17756 29886 17808
rect 31726 17796 31754 17836
rect 32033 17833 32045 17867
rect 32079 17864 32091 17867
rect 32766 17864 32772 17876
rect 32079 17836 32772 17864
rect 32079 17833 32091 17836
rect 32033 17827 32091 17833
rect 32766 17824 32772 17836
rect 32824 17824 32830 17876
rect 37182 17824 37188 17876
rect 37240 17864 37246 17876
rect 38838 17864 38844 17876
rect 37240 17836 38844 17864
rect 37240 17824 37246 17836
rect 38838 17824 38844 17836
rect 38896 17824 38902 17876
rect 38930 17824 38936 17876
rect 38988 17864 38994 17876
rect 38988 17836 52960 17864
rect 38988 17824 38994 17836
rect 31726 17768 36584 17796
rect 31018 17688 31024 17740
rect 31076 17728 31082 17740
rect 31665 17731 31723 17737
rect 31665 17728 31677 17731
rect 31076 17700 31677 17728
rect 31076 17688 31082 17700
rect 31665 17697 31677 17700
rect 31711 17697 31723 17731
rect 31665 17691 31723 17697
rect 31772 17700 32444 17728
rect 28537 17663 28595 17669
rect 28537 17629 28549 17663
rect 28583 17629 28595 17663
rect 28537 17623 28595 17629
rect 28634 17663 28692 17669
rect 28634 17629 28646 17663
rect 28680 17629 28692 17663
rect 29733 17663 29791 17669
rect 29733 17660 29745 17663
rect 28634 17623 28692 17629
rect 28828 17632 29745 17660
rect 28445 17595 28503 17601
rect 28445 17561 28457 17595
rect 28491 17561 28503 17595
rect 28445 17555 28503 17561
rect 27663 17496 28212 17524
rect 28460 17524 28488 17555
rect 28718 17524 28724 17536
rect 28460 17496 28724 17524
rect 27663 17493 27675 17496
rect 27617 17487 27675 17493
rect 28718 17484 28724 17496
rect 28776 17484 28782 17536
rect 28828 17533 28856 17632
rect 29733 17629 29745 17632
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 30006 17620 30012 17672
rect 30064 17620 30070 17672
rect 31772 17660 31800 17700
rect 31726 17632 31800 17660
rect 31849 17663 31907 17669
rect 28902 17552 28908 17604
rect 28960 17592 28966 17604
rect 31726 17592 31754 17632
rect 31849 17629 31861 17663
rect 31895 17660 31907 17663
rect 31938 17660 31944 17672
rect 31895 17632 31944 17660
rect 31895 17629 31907 17632
rect 31849 17623 31907 17629
rect 31938 17620 31944 17632
rect 31996 17620 32002 17672
rect 32416 17660 32444 17700
rect 32490 17688 32496 17740
rect 32548 17688 32554 17740
rect 33870 17728 33876 17740
rect 32600 17700 33876 17728
rect 32600 17660 32628 17700
rect 33870 17688 33876 17700
rect 33928 17688 33934 17740
rect 34054 17688 34060 17740
rect 34112 17728 34118 17740
rect 35069 17731 35127 17737
rect 35069 17728 35081 17731
rect 34112 17700 35081 17728
rect 34112 17688 34118 17700
rect 35069 17697 35081 17700
rect 35115 17697 35127 17731
rect 35069 17691 35127 17697
rect 32416 17632 32628 17660
rect 32677 17663 32735 17669
rect 32677 17629 32689 17663
rect 32723 17629 32735 17663
rect 32677 17623 32735 17629
rect 32692 17592 32720 17623
rect 33778 17620 33784 17672
rect 33836 17620 33842 17672
rect 33888 17660 33916 17688
rect 34790 17660 34796 17672
rect 33888 17632 34796 17660
rect 34790 17620 34796 17632
rect 34848 17620 34854 17672
rect 34885 17663 34943 17669
rect 34885 17629 34897 17663
rect 34931 17660 34943 17663
rect 36556 17660 36584 17768
rect 38746 17756 38752 17808
rect 38804 17756 38810 17808
rect 38856 17796 38884 17824
rect 38856 17768 40264 17796
rect 40236 17740 40264 17768
rect 41230 17756 41236 17808
rect 41288 17796 41294 17808
rect 41601 17799 41659 17805
rect 41601 17796 41613 17799
rect 41288 17768 41613 17796
rect 41288 17756 41294 17768
rect 41601 17765 41613 17768
rect 41647 17765 41659 17799
rect 41601 17759 41659 17765
rect 48501 17799 48559 17805
rect 48501 17765 48513 17799
rect 48547 17796 48559 17799
rect 48682 17796 48688 17808
rect 48547 17768 48688 17796
rect 48547 17765 48559 17768
rect 48501 17759 48559 17765
rect 48682 17756 48688 17768
rect 48740 17756 48746 17808
rect 52932 17796 52960 17836
rect 53006 17824 53012 17876
rect 53064 17864 53070 17876
rect 54478 17864 54484 17876
rect 53064 17836 54484 17864
rect 53064 17824 53070 17836
rect 54478 17824 54484 17836
rect 54536 17824 54542 17876
rect 57146 17824 57152 17876
rect 57204 17864 57210 17876
rect 58253 17867 58311 17873
rect 58253 17864 58265 17867
rect 57204 17836 58265 17864
rect 57204 17824 57210 17836
rect 58253 17833 58265 17836
rect 58299 17833 58311 17867
rect 58253 17827 58311 17833
rect 52932 17768 55812 17796
rect 39206 17688 39212 17740
rect 39264 17728 39270 17740
rect 39393 17731 39451 17737
rect 39393 17728 39405 17731
rect 39264 17700 39405 17728
rect 39264 17688 39270 17700
rect 39393 17697 39405 17700
rect 39439 17728 39451 17731
rect 39850 17728 39856 17740
rect 39439 17700 39856 17728
rect 39439 17697 39451 17700
rect 39393 17691 39451 17697
rect 39850 17688 39856 17700
rect 39908 17688 39914 17740
rect 40218 17688 40224 17740
rect 40276 17688 40282 17740
rect 48130 17688 48136 17740
rect 48188 17728 48194 17740
rect 48188 17700 51028 17728
rect 48188 17688 48194 17700
rect 40494 17669 40500 17672
rect 40488 17660 40500 17669
rect 34931 17632 36492 17660
rect 36556 17632 39344 17660
rect 40455 17632 40500 17660
rect 34931 17629 34943 17632
rect 34885 17623 34943 17629
rect 28960 17564 31754 17592
rect 31956 17564 32720 17592
rect 28960 17552 28966 17564
rect 28813 17527 28871 17533
rect 28813 17493 28825 17527
rect 28859 17493 28871 17527
rect 28813 17487 28871 17493
rect 30193 17527 30251 17533
rect 30193 17493 30205 17527
rect 30239 17524 30251 17527
rect 30282 17524 30288 17536
rect 30239 17496 30288 17524
rect 30239 17493 30251 17496
rect 30193 17487 30251 17493
rect 30282 17484 30288 17496
rect 30340 17484 30346 17536
rect 31386 17484 31392 17536
rect 31444 17524 31450 17536
rect 31956 17524 31984 17564
rect 33686 17552 33692 17604
rect 33744 17592 33750 17604
rect 36464 17592 36492 17632
rect 36906 17592 36912 17604
rect 33744 17564 34008 17592
rect 36464 17564 36912 17592
rect 33744 17552 33750 17564
rect 31444 17496 31984 17524
rect 31444 17484 31450 17496
rect 32766 17484 32772 17536
rect 32824 17524 32830 17536
rect 32861 17527 32919 17533
rect 32861 17524 32873 17527
rect 32824 17496 32873 17524
rect 32824 17484 32830 17496
rect 32861 17493 32873 17496
rect 32907 17493 32919 17527
rect 32861 17487 32919 17493
rect 33226 17484 33232 17536
rect 33284 17524 33290 17536
rect 33413 17527 33471 17533
rect 33413 17524 33425 17527
rect 33284 17496 33425 17524
rect 33284 17484 33290 17496
rect 33413 17493 33425 17496
rect 33459 17493 33471 17527
rect 33413 17487 33471 17493
rect 33870 17484 33876 17536
rect 33928 17484 33934 17536
rect 33980 17524 34008 17564
rect 36906 17552 36912 17564
rect 36964 17552 36970 17604
rect 38654 17552 38660 17604
rect 38712 17592 38718 17604
rect 39117 17595 39175 17601
rect 39117 17592 39129 17595
rect 38712 17564 39129 17592
rect 38712 17552 38718 17564
rect 39117 17561 39129 17564
rect 39163 17561 39175 17595
rect 39117 17555 39175 17561
rect 39206 17552 39212 17604
rect 39264 17552 39270 17604
rect 39316 17592 39344 17632
rect 40488 17623 40500 17632
rect 40494 17620 40500 17623
rect 40552 17620 40558 17672
rect 47946 17620 47952 17672
rect 48004 17620 48010 17672
rect 48332 17669 48360 17700
rect 51000 17672 51028 17700
rect 51552 17700 51764 17728
rect 48317 17663 48375 17669
rect 48317 17629 48329 17663
rect 48363 17660 48375 17663
rect 50617 17663 50675 17669
rect 48363 17632 48397 17660
rect 48363 17629 48375 17632
rect 48317 17623 48375 17629
rect 50617 17629 50629 17663
rect 50663 17629 50675 17663
rect 50617 17623 50675 17629
rect 39316 17564 41414 17592
rect 38930 17524 38936 17536
rect 33980 17496 38936 17524
rect 38930 17484 38936 17496
rect 38988 17484 38994 17536
rect 41386 17524 41414 17564
rect 46934 17552 46940 17604
rect 46992 17592 46998 17604
rect 48133 17595 48191 17601
rect 48133 17592 48145 17595
rect 46992 17564 48145 17592
rect 46992 17552 46998 17564
rect 48133 17561 48145 17564
rect 48179 17561 48191 17595
rect 48133 17555 48191 17561
rect 48225 17595 48283 17601
rect 48225 17561 48237 17595
rect 48271 17592 48283 17595
rect 49970 17592 49976 17604
rect 48271 17564 49976 17592
rect 48271 17561 48283 17564
rect 48225 17555 48283 17561
rect 49970 17552 49976 17564
rect 50028 17552 50034 17604
rect 50632 17524 50660 17623
rect 50982 17620 50988 17672
rect 51040 17620 51046 17672
rect 50801 17595 50859 17601
rect 50801 17561 50813 17595
rect 50847 17561 50859 17595
rect 50801 17555 50859 17561
rect 50893 17595 50951 17601
rect 50893 17561 50905 17595
rect 50939 17592 50951 17595
rect 51552 17592 51580 17700
rect 51626 17620 51632 17672
rect 51684 17620 51690 17672
rect 51736 17660 51764 17700
rect 54754 17688 54760 17740
rect 54812 17728 54818 17740
rect 55677 17731 55735 17737
rect 55677 17728 55689 17731
rect 54812 17700 55689 17728
rect 54812 17688 54818 17700
rect 55677 17697 55689 17700
rect 55723 17697 55735 17731
rect 55677 17691 55735 17697
rect 53006 17660 53012 17672
rect 51736 17632 53012 17660
rect 53006 17620 53012 17632
rect 53064 17620 53070 17672
rect 53834 17620 53840 17672
rect 53892 17660 53898 17672
rect 55493 17663 55551 17669
rect 55493 17660 55505 17663
rect 53892 17632 55505 17660
rect 53892 17620 53898 17632
rect 55493 17629 55505 17632
rect 55539 17629 55551 17663
rect 55784 17660 55812 17768
rect 55858 17688 55864 17740
rect 55916 17728 55922 17740
rect 56873 17731 56931 17737
rect 56873 17728 56885 17731
rect 55916 17700 56885 17728
rect 55916 17688 55922 17700
rect 56873 17697 56885 17700
rect 56919 17697 56931 17731
rect 56873 17691 56931 17697
rect 58250 17660 58256 17672
rect 55784 17632 58256 17660
rect 55493 17623 55551 17629
rect 58250 17620 58256 17632
rect 58308 17620 58314 17672
rect 51902 17601 51908 17604
rect 50939 17564 51580 17592
rect 50939 17561 50951 17564
rect 50893 17555 50951 17561
rect 51896 17555 51908 17601
rect 41386 17496 50660 17524
rect 50816 17524 50844 17555
rect 51902 17552 51908 17555
rect 51960 17552 51966 17604
rect 56318 17552 56324 17604
rect 56376 17592 56382 17604
rect 57118 17595 57176 17601
rect 57118 17592 57130 17595
rect 56376 17564 57130 17592
rect 56376 17552 56382 17564
rect 57118 17561 57130 17564
rect 57164 17561 57176 17595
rect 57118 17555 57176 17561
rect 51074 17524 51080 17536
rect 50816 17496 51080 17524
rect 51074 17484 51080 17496
rect 51132 17484 51138 17536
rect 51169 17527 51227 17533
rect 51169 17493 51181 17527
rect 51215 17524 51227 17527
rect 51626 17524 51632 17536
rect 51215 17496 51632 17524
rect 51215 17493 51227 17496
rect 51169 17487 51227 17493
rect 51626 17484 51632 17496
rect 51684 17484 51690 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 8478 17280 8484 17332
rect 8536 17320 8542 17332
rect 8757 17323 8815 17329
rect 8757 17320 8769 17323
rect 8536 17292 8769 17320
rect 8536 17280 8542 17292
rect 8757 17289 8769 17292
rect 8803 17289 8815 17323
rect 8757 17283 8815 17289
rect 15378 17280 15384 17332
rect 15436 17280 15442 17332
rect 17221 17323 17279 17329
rect 17221 17289 17233 17323
rect 17267 17289 17279 17323
rect 17221 17283 17279 17289
rect 6454 17212 6460 17264
rect 6512 17252 6518 17264
rect 11146 17252 11152 17264
rect 6512 17224 11152 17252
rect 6512 17212 6518 17224
rect 11146 17212 11152 17224
rect 11204 17212 11210 17264
rect 17236 17252 17264 17283
rect 17954 17280 17960 17332
rect 18012 17280 18018 17332
rect 18785 17323 18843 17329
rect 18785 17289 18797 17323
rect 18831 17320 18843 17323
rect 18874 17320 18880 17332
rect 18831 17292 18880 17320
rect 18831 17289 18843 17292
rect 18785 17283 18843 17289
rect 18874 17280 18880 17292
rect 18932 17280 18938 17332
rect 19150 17280 19156 17332
rect 19208 17320 19214 17332
rect 20717 17323 20775 17329
rect 19208 17292 20024 17320
rect 19208 17280 19214 17292
rect 19996 17252 20024 17292
rect 20717 17289 20729 17323
rect 20763 17320 20775 17323
rect 20990 17320 20996 17332
rect 20763 17292 20996 17320
rect 20763 17289 20775 17292
rect 20717 17283 20775 17289
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 24946 17280 24952 17332
rect 25004 17280 25010 17332
rect 25222 17280 25228 17332
rect 25280 17280 25286 17332
rect 25332 17292 36584 17320
rect 22646 17252 22652 17264
rect 16040 17224 17172 17252
rect 17236 17224 19932 17252
rect 19996 17224 22652 17252
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17184 1639 17187
rect 2406 17184 2412 17196
rect 1627 17156 2412 17184
rect 1627 17153 1639 17156
rect 1581 17147 1639 17153
rect 2406 17144 2412 17156
rect 2464 17144 2470 17196
rect 8570 17144 8576 17196
rect 8628 17144 8634 17196
rect 15286 17144 15292 17196
rect 15344 17144 15350 17196
rect 15473 17187 15531 17193
rect 15473 17153 15485 17187
rect 15519 17184 15531 17187
rect 15562 17184 15568 17196
rect 15519 17156 15568 17184
rect 15519 17153 15531 17156
rect 15473 17147 15531 17153
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 16040 17193 16068 17224
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17153 16083 17187
rect 16025 17147 16083 17153
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17153 17095 17187
rect 17144 17184 17172 17224
rect 17144 17156 17724 17184
rect 17037 17147 17095 17153
rect 934 17076 940 17128
rect 992 17116 998 17128
rect 1765 17119 1823 17125
rect 1765 17116 1777 17119
rect 992 17088 1777 17116
rect 992 17076 998 17088
rect 1765 17085 1777 17088
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 17052 17048 17080 17147
rect 17696 17116 17724 17156
rect 17770 17144 17776 17196
rect 17828 17144 17834 17196
rect 18601 17187 18659 17193
rect 18601 17153 18613 17187
rect 18647 17184 18659 17187
rect 18782 17184 18788 17196
rect 18647 17156 18788 17184
rect 18647 17153 18659 17156
rect 18601 17147 18659 17153
rect 18782 17144 18788 17156
rect 18840 17144 18846 17196
rect 19334 17144 19340 17196
rect 19392 17144 19398 17196
rect 19904 17193 19932 17224
rect 22646 17212 22652 17224
rect 22704 17212 22710 17264
rect 24670 17212 24676 17264
rect 24728 17252 24734 17264
rect 25332 17252 25360 17292
rect 24728 17224 25360 17252
rect 24728 17212 24734 17224
rect 25406 17212 25412 17264
rect 25464 17212 25470 17264
rect 26050 17212 26056 17264
rect 26108 17252 26114 17264
rect 28077 17255 28135 17261
rect 28077 17252 28089 17255
rect 26108 17224 28089 17252
rect 26108 17212 26114 17224
rect 28077 17221 28089 17224
rect 28123 17221 28135 17255
rect 28077 17215 28135 17221
rect 28166 17212 28172 17264
rect 28224 17212 28230 17264
rect 28442 17212 28448 17264
rect 28500 17252 28506 17264
rect 33686 17252 33692 17264
rect 28500 17224 33692 17252
rect 28500 17212 28506 17224
rect 33686 17212 33692 17224
rect 33744 17212 33750 17264
rect 33864 17255 33922 17261
rect 33864 17221 33876 17255
rect 33910 17252 33922 17255
rect 33962 17252 33968 17264
rect 33910 17224 33968 17252
rect 33910 17221 33922 17224
rect 33864 17215 33922 17221
rect 33962 17212 33968 17224
rect 34020 17212 34026 17264
rect 36556 17252 36584 17292
rect 38286 17280 38292 17332
rect 38344 17280 38350 17332
rect 51813 17323 51871 17329
rect 38396 17292 51764 17320
rect 38396 17252 38424 17292
rect 36556 17224 38424 17252
rect 38657 17255 38715 17261
rect 38657 17221 38669 17255
rect 38703 17252 38715 17255
rect 39206 17252 39212 17264
rect 38703 17224 39212 17252
rect 38703 17221 38715 17224
rect 38657 17215 38715 17221
rect 39206 17212 39212 17224
rect 39264 17212 39270 17264
rect 40880 17224 41092 17252
rect 19889 17187 19947 17193
rect 19889 17153 19901 17187
rect 19935 17153 19947 17187
rect 19889 17147 19947 17153
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17184 20131 17187
rect 20530 17184 20536 17196
rect 20119 17156 20536 17184
rect 20119 17153 20131 17156
rect 20073 17147 20131 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 21085 17187 21143 17193
rect 21085 17153 21097 17187
rect 21131 17184 21143 17187
rect 21910 17184 21916 17196
rect 21131 17156 21916 17184
rect 21131 17153 21143 17156
rect 21085 17147 21143 17153
rect 21910 17144 21916 17156
rect 21968 17144 21974 17196
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17184 22063 17187
rect 24118 17184 24124 17196
rect 22051 17156 24124 17184
rect 22051 17153 22063 17156
rect 22005 17147 22063 17153
rect 24118 17144 24124 17156
rect 24176 17144 24182 17196
rect 24854 17144 24860 17196
rect 24912 17184 24918 17196
rect 25041 17187 25099 17193
rect 25041 17184 25053 17187
rect 24912 17156 25053 17184
rect 24912 17144 24918 17156
rect 25041 17153 25053 17156
rect 25087 17153 25099 17187
rect 25153 17187 25211 17193
rect 25153 17184 25165 17187
rect 25041 17147 25099 17153
rect 25148 17153 25165 17184
rect 25199 17153 25211 17187
rect 25148 17147 25211 17153
rect 19981 17119 20039 17125
rect 19981 17116 19993 17119
rect 17696 17088 19993 17116
rect 19981 17085 19993 17088
rect 20027 17085 20039 17119
rect 19981 17079 20039 17085
rect 20346 17076 20352 17128
rect 20404 17076 20410 17128
rect 20441 17119 20499 17125
rect 20441 17085 20453 17119
rect 20487 17116 20499 17119
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 20487 17088 21189 17116
rect 20487 17085 20499 17088
rect 20441 17079 20499 17085
rect 21177 17085 21189 17088
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 21361 17119 21419 17125
rect 21361 17085 21373 17119
rect 21407 17116 21419 17119
rect 21450 17116 21456 17128
rect 21407 17088 21456 17116
rect 21407 17085 21419 17088
rect 21361 17079 21419 17085
rect 19242 17048 19248 17060
rect 17052 17020 19248 17048
rect 19242 17008 19248 17020
rect 19300 17008 19306 17060
rect 20364 17048 20392 17076
rect 19444 17020 20392 17048
rect 21192 17048 21220 17079
rect 21450 17076 21456 17088
rect 21508 17076 21514 17128
rect 24762 17076 24768 17128
rect 24820 17116 24826 17128
rect 25148 17116 25176 17147
rect 27614 17144 27620 17196
rect 27672 17184 27678 17196
rect 27893 17187 27951 17193
rect 27893 17184 27905 17187
rect 27672 17156 27905 17184
rect 27672 17144 27678 17156
rect 27893 17153 27905 17156
rect 27939 17153 27951 17187
rect 27893 17147 27951 17153
rect 27982 17144 27988 17196
rect 28040 17184 28046 17196
rect 28313 17187 28371 17193
rect 28313 17184 28325 17187
rect 28040 17156 28325 17184
rect 28040 17144 28046 17156
rect 28313 17153 28325 17156
rect 28359 17184 28371 17187
rect 28810 17184 28816 17196
rect 28359 17156 28816 17184
rect 28359 17153 28371 17156
rect 28313 17147 28371 17153
rect 28810 17144 28816 17156
rect 28868 17184 28874 17196
rect 31386 17184 31392 17196
rect 28868 17156 31392 17184
rect 28868 17144 28874 17156
rect 31386 17144 31392 17156
rect 31444 17144 31450 17196
rect 32766 17144 32772 17196
rect 32824 17144 32830 17196
rect 32858 17144 32864 17196
rect 32916 17184 32922 17196
rect 33597 17187 33655 17193
rect 33597 17184 33609 17187
rect 32916 17156 33609 17184
rect 32916 17144 32922 17156
rect 33597 17153 33609 17156
rect 33643 17153 33655 17187
rect 40880 17184 40908 17224
rect 33597 17147 33655 17153
rect 33704 17156 40908 17184
rect 28994 17116 29000 17128
rect 24820 17088 25176 17116
rect 25332 17088 29000 17116
rect 24820 17076 24826 17088
rect 22278 17048 22284 17060
rect 21192 17020 22284 17048
rect 2406 16940 2412 16992
rect 2464 16940 2470 16992
rect 16209 16983 16267 16989
rect 16209 16949 16221 16983
rect 16255 16980 16267 16983
rect 17126 16980 17132 16992
rect 16255 16952 17132 16980
rect 16255 16949 16267 16952
rect 16209 16943 16267 16949
rect 17126 16940 17132 16952
rect 17184 16940 17190 16992
rect 17218 16940 17224 16992
rect 17276 16980 17282 16992
rect 19444 16980 19472 17020
rect 22278 17008 22284 17020
rect 22336 17048 22342 17060
rect 25332 17048 25360 17088
rect 28994 17076 29000 17088
rect 29052 17076 29058 17128
rect 32214 17076 32220 17128
rect 32272 17116 32278 17128
rect 32493 17119 32551 17125
rect 32493 17116 32505 17119
rect 32272 17088 32505 17116
rect 32272 17076 32278 17088
rect 32493 17085 32505 17088
rect 32539 17085 32551 17119
rect 32493 17079 32551 17085
rect 32582 17076 32588 17128
rect 32640 17076 32646 17128
rect 32674 17076 32680 17128
rect 32732 17116 32738 17128
rect 33410 17116 33416 17128
rect 32732 17088 33416 17116
rect 32732 17076 32738 17088
rect 33410 17076 33416 17088
rect 33468 17076 33474 17128
rect 33502 17076 33508 17128
rect 33560 17116 33566 17128
rect 33704 17116 33732 17156
rect 40954 17144 40960 17196
rect 41012 17144 41018 17196
rect 41064 17184 41092 17224
rect 41138 17212 41144 17264
rect 41196 17252 41202 17264
rect 51736 17252 51764 17292
rect 51813 17289 51825 17323
rect 51859 17320 51871 17323
rect 51902 17320 51908 17332
rect 51859 17292 51908 17320
rect 51859 17289 51871 17292
rect 51813 17283 51871 17289
rect 51902 17280 51908 17292
rect 51960 17280 51966 17332
rect 53926 17280 53932 17332
rect 53984 17320 53990 17332
rect 55950 17320 55956 17332
rect 53984 17292 55956 17320
rect 53984 17280 53990 17292
rect 55950 17280 55956 17292
rect 56008 17280 56014 17332
rect 56318 17280 56324 17332
rect 56376 17280 56382 17332
rect 54570 17252 54576 17264
rect 41196 17224 51580 17252
rect 51736 17224 54576 17252
rect 41196 17212 41202 17224
rect 47946 17184 47952 17196
rect 41064 17156 47952 17184
rect 47946 17144 47952 17156
rect 48004 17144 48010 17196
rect 51442 17144 51448 17196
rect 51500 17144 51506 17196
rect 38749 17119 38807 17125
rect 33560 17088 33732 17116
rect 34624 17088 38654 17116
rect 33560 17076 33566 17088
rect 22336 17020 25360 17048
rect 22336 17008 22342 17020
rect 27706 17008 27712 17060
rect 27764 17048 27770 17060
rect 27890 17048 27896 17060
rect 27764 17020 27896 17048
rect 27764 17008 27770 17020
rect 27890 17008 27896 17020
rect 27948 17008 27954 17060
rect 28445 17051 28503 17057
rect 28445 17017 28457 17051
rect 28491 17048 28503 17051
rect 28491 17020 33640 17048
rect 28491 17017 28503 17020
rect 28445 17011 28503 17017
rect 17276 16952 19472 16980
rect 17276 16940 17282 16952
rect 19518 16940 19524 16992
rect 19576 16940 19582 16992
rect 20346 16940 20352 16992
rect 20404 16980 20410 16992
rect 22189 16983 22247 16989
rect 22189 16980 22201 16983
rect 20404 16952 22201 16980
rect 20404 16940 20410 16952
rect 22189 16949 22201 16952
rect 22235 16949 22247 16983
rect 22189 16943 22247 16949
rect 23658 16940 23664 16992
rect 23716 16980 23722 16992
rect 29178 16980 29184 16992
rect 23716 16952 29184 16980
rect 23716 16940 23722 16952
rect 29178 16940 29184 16952
rect 29236 16940 29242 16992
rect 32309 16983 32367 16989
rect 32309 16949 32321 16983
rect 32355 16980 32367 16983
rect 33502 16980 33508 16992
rect 32355 16952 33508 16980
rect 32355 16949 32367 16952
rect 32309 16943 32367 16949
rect 33502 16940 33508 16952
rect 33560 16940 33566 16992
rect 33612 16980 33640 17020
rect 34624 16980 34652 17088
rect 38626 17048 38654 17088
rect 38749 17085 38761 17119
rect 38795 17116 38807 17119
rect 38838 17116 38844 17128
rect 38795 17088 38844 17116
rect 38795 17085 38807 17088
rect 38749 17079 38807 17085
rect 38838 17076 38844 17088
rect 38896 17076 38902 17128
rect 38933 17119 38991 17125
rect 38933 17085 38945 17119
rect 38979 17116 38991 17119
rect 39942 17116 39948 17128
rect 38979 17088 39948 17116
rect 38979 17085 38991 17088
rect 38933 17079 38991 17085
rect 39942 17076 39948 17088
rect 40000 17076 40006 17128
rect 40862 17076 40868 17128
rect 40920 17116 40926 17128
rect 41049 17119 41107 17125
rect 41049 17116 41061 17119
rect 40920 17088 41061 17116
rect 40920 17076 40926 17088
rect 41049 17085 41061 17088
rect 41095 17085 41107 17119
rect 41049 17079 41107 17085
rect 41233 17119 41291 17125
rect 41233 17085 41245 17119
rect 41279 17116 41291 17119
rect 41322 17116 41328 17128
rect 41279 17088 41328 17116
rect 41279 17085 41291 17088
rect 41233 17079 41291 17085
rect 41322 17076 41328 17088
rect 41380 17076 41386 17128
rect 51552 17116 51580 17224
rect 54570 17212 54576 17224
rect 54628 17212 54634 17264
rect 58066 17252 58072 17264
rect 54680 17224 58072 17252
rect 51626 17144 51632 17196
rect 51684 17144 51690 17196
rect 51736 17156 54064 17184
rect 51736 17116 51764 17156
rect 51552 17088 51764 17116
rect 51810 17076 51816 17128
rect 51868 17116 51874 17128
rect 53926 17116 53932 17128
rect 51868 17088 53932 17116
rect 51868 17076 51874 17088
rect 53926 17076 53932 17088
rect 53984 17076 53990 17128
rect 54036 17116 54064 17156
rect 54110 17144 54116 17196
rect 54168 17144 54174 17196
rect 54680 17116 54708 17224
rect 58066 17212 58072 17224
rect 58124 17212 58130 17264
rect 54941 17187 54999 17193
rect 54941 17153 54953 17187
rect 54987 17153 54999 17187
rect 54941 17147 54999 17153
rect 54036 17088 54708 17116
rect 54956 17048 54984 17147
rect 55122 17144 55128 17196
rect 55180 17144 55186 17196
rect 55217 17187 55275 17193
rect 55217 17153 55229 17187
rect 55263 17153 55275 17187
rect 55217 17147 55275 17153
rect 38626 17020 54984 17048
rect 33612 16952 34652 16980
rect 34790 16940 34796 16992
rect 34848 16980 34854 16992
rect 34977 16983 35035 16989
rect 34977 16980 34989 16983
rect 34848 16952 34989 16980
rect 34848 16940 34854 16952
rect 34977 16949 34989 16952
rect 35023 16949 35035 16983
rect 34977 16943 35035 16949
rect 36906 16940 36912 16992
rect 36964 16980 36970 16992
rect 40218 16980 40224 16992
rect 36964 16952 40224 16980
rect 36964 16940 36970 16952
rect 40218 16940 40224 16952
rect 40276 16940 40282 16992
rect 40589 16983 40647 16989
rect 40589 16949 40601 16983
rect 40635 16980 40647 16983
rect 44174 16980 44180 16992
rect 40635 16952 44180 16980
rect 40635 16949 40647 16952
rect 40589 16943 40647 16949
rect 44174 16940 44180 16952
rect 44232 16940 44238 16992
rect 54294 16940 54300 16992
rect 54352 16940 54358 16992
rect 55232 16980 55260 17147
rect 55306 17144 55312 17196
rect 55364 17144 55370 17196
rect 56137 17187 56195 17193
rect 56137 17184 56149 17187
rect 55508 17156 56149 17184
rect 55508 17057 55536 17156
rect 56137 17153 56149 17156
rect 56183 17153 56195 17187
rect 56137 17147 56195 17153
rect 56226 17144 56232 17196
rect 56284 17184 56290 17196
rect 57057 17187 57115 17193
rect 57057 17184 57069 17187
rect 56284 17156 57069 17184
rect 56284 17144 56290 17156
rect 57057 17153 57069 17156
rect 57103 17153 57115 17187
rect 57057 17147 57115 17153
rect 55950 17076 55956 17128
rect 56008 17076 56014 17128
rect 57333 17119 57391 17125
rect 57333 17085 57345 17119
rect 57379 17116 57391 17119
rect 58986 17116 58992 17128
rect 57379 17088 58992 17116
rect 57379 17085 57391 17088
rect 57333 17079 57391 17085
rect 58986 17076 58992 17088
rect 59044 17076 59050 17128
rect 55493 17051 55551 17057
rect 55493 17017 55505 17051
rect 55539 17017 55551 17051
rect 55493 17011 55551 17017
rect 57146 16980 57152 16992
rect 55232 16952 57152 16980
rect 57146 16940 57152 16952
rect 57204 16940 57210 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 16206 16736 16212 16788
rect 16264 16736 16270 16788
rect 18782 16736 18788 16788
rect 18840 16776 18846 16788
rect 18840 16748 22094 16776
rect 18840 16736 18846 16748
rect 12802 16668 12808 16720
rect 12860 16708 12866 16720
rect 12860 16680 13676 16708
rect 12860 16668 12866 16680
rect 13446 16600 13452 16652
rect 13504 16600 13510 16652
rect 13648 16649 13676 16680
rect 18690 16668 18696 16720
rect 18748 16668 18754 16720
rect 19518 16708 19524 16720
rect 18892 16680 19524 16708
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16609 13691 16643
rect 18892 16640 18920 16680
rect 19518 16668 19524 16680
rect 19576 16668 19582 16720
rect 19613 16711 19671 16717
rect 19613 16677 19625 16711
rect 19659 16677 19671 16711
rect 22066 16708 22094 16748
rect 22646 16736 22652 16788
rect 22704 16736 22710 16788
rect 28902 16776 28908 16788
rect 22756 16748 28908 16776
rect 22756 16708 22784 16748
rect 28902 16736 28908 16748
rect 28960 16736 28966 16788
rect 28994 16736 29000 16788
rect 29052 16776 29058 16788
rect 41138 16776 41144 16788
rect 29052 16748 41144 16776
rect 29052 16736 29058 16748
rect 41138 16736 41144 16748
rect 41196 16736 41202 16788
rect 52914 16736 52920 16788
rect 52972 16776 52978 16788
rect 55306 16776 55312 16788
rect 52972 16748 55312 16776
rect 52972 16736 52978 16748
rect 55306 16736 55312 16748
rect 55364 16736 55370 16788
rect 56594 16736 56600 16788
rect 56652 16776 56658 16788
rect 57149 16779 57207 16785
rect 57149 16776 57161 16779
rect 56652 16748 57161 16776
rect 56652 16736 56658 16748
rect 57149 16745 57161 16748
rect 57195 16745 57207 16779
rect 57149 16739 57207 16745
rect 22066 16680 22784 16708
rect 19613 16671 19671 16677
rect 13633 16603 13691 16609
rect 16224 16612 16804 16640
rect 1581 16575 1639 16581
rect 1581 16541 1593 16575
rect 1627 16572 1639 16575
rect 10410 16572 10416 16584
rect 1627 16544 10416 16572
rect 1627 16541 1639 16544
rect 1581 16535 1639 16541
rect 10410 16532 10416 16544
rect 10468 16532 10474 16584
rect 12250 16532 12256 16584
rect 12308 16532 12314 16584
rect 13354 16532 13360 16584
rect 13412 16532 13418 16584
rect 16224 16581 16252 16612
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16541 13599 16575
rect 13541 16535 13599 16541
rect 16209 16575 16267 16581
rect 16209 16541 16221 16575
rect 16255 16541 16267 16575
rect 16209 16535 16267 16541
rect 934 16464 940 16516
rect 992 16504 998 16516
rect 1857 16507 1915 16513
rect 1857 16504 1869 16507
rect 992 16476 1869 16504
rect 992 16464 998 16476
rect 1857 16473 1869 16476
rect 1903 16473 1915 16507
rect 1857 16467 1915 16473
rect 11146 16464 11152 16516
rect 11204 16504 11210 16516
rect 13556 16504 13584 16535
rect 16390 16532 16396 16584
rect 16448 16532 16454 16584
rect 13906 16504 13912 16516
rect 11204 16476 13216 16504
rect 13556 16476 13912 16504
rect 11204 16464 11210 16476
rect 11698 16396 11704 16448
rect 11756 16436 11762 16448
rect 13188 16445 13216 16476
rect 13906 16464 13912 16476
rect 13964 16464 13970 16516
rect 16776 16504 16804 16612
rect 18708 16612 18920 16640
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 16942 16572 16948 16584
rect 16899 16544 16948 16572
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 17126 16581 17132 16584
rect 17120 16572 17132 16581
rect 17087 16544 17132 16572
rect 17120 16535 17132 16544
rect 17126 16532 17132 16535
rect 17184 16532 17190 16584
rect 18708 16581 18736 16612
rect 19242 16600 19248 16652
rect 19300 16640 19306 16652
rect 19628 16640 19656 16671
rect 31754 16668 31760 16720
rect 31812 16708 31818 16720
rect 32766 16708 32772 16720
rect 31812 16680 32772 16708
rect 31812 16668 31818 16680
rect 32766 16668 32772 16680
rect 32824 16668 32830 16720
rect 40678 16668 40684 16720
rect 40736 16708 40742 16720
rect 41322 16708 41328 16720
rect 40736 16680 41328 16708
rect 40736 16668 40742 16680
rect 41322 16668 41328 16680
rect 41380 16708 41386 16720
rect 41380 16680 41736 16708
rect 41380 16668 41386 16680
rect 19300 16612 19656 16640
rect 19300 16600 19306 16612
rect 20806 16600 20812 16652
rect 20864 16600 20870 16652
rect 25961 16643 26019 16649
rect 25961 16609 25973 16643
rect 26007 16609 26019 16643
rect 25961 16603 26019 16609
rect 18693 16575 18751 16581
rect 18693 16541 18705 16575
rect 18739 16541 18751 16575
rect 18693 16535 18751 16541
rect 18874 16532 18880 16584
rect 18932 16532 18938 16584
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 17218 16504 17224 16516
rect 16776 16476 17224 16504
rect 17218 16464 17224 16476
rect 17276 16464 17282 16516
rect 19444 16504 19472 16535
rect 19518 16532 19524 16584
rect 19576 16572 19582 16584
rect 20165 16575 20223 16581
rect 20165 16572 20177 16575
rect 19576 16544 20177 16572
rect 19576 16532 19582 16544
rect 20165 16541 20177 16544
rect 20211 16541 20223 16575
rect 20165 16535 20223 16541
rect 20346 16532 20352 16584
rect 20404 16532 20410 16584
rect 21082 16581 21088 16584
rect 21076 16572 21088 16581
rect 21043 16544 21088 16572
rect 21076 16535 21088 16544
rect 21082 16532 21088 16535
rect 21140 16532 21146 16584
rect 22646 16532 22652 16584
rect 22704 16532 22710 16584
rect 22830 16532 22836 16584
rect 22888 16532 22894 16584
rect 24578 16532 24584 16584
rect 24636 16572 24642 16584
rect 25976 16572 26004 16603
rect 27522 16600 27528 16652
rect 27580 16640 27586 16652
rect 27709 16643 27767 16649
rect 27709 16640 27721 16643
rect 27580 16612 27721 16640
rect 27580 16600 27586 16612
rect 27709 16609 27721 16612
rect 27755 16640 27767 16643
rect 28442 16640 28448 16652
rect 27755 16612 28448 16640
rect 27755 16609 27767 16612
rect 27709 16603 27767 16609
rect 28442 16600 28448 16612
rect 28500 16600 28506 16652
rect 28626 16600 28632 16652
rect 28684 16640 28690 16652
rect 28994 16640 29000 16652
rect 28684 16612 29000 16640
rect 28684 16600 28690 16612
rect 28994 16600 29000 16612
rect 29052 16600 29058 16652
rect 30006 16600 30012 16652
rect 30064 16640 30070 16652
rect 32493 16643 32551 16649
rect 32493 16640 32505 16643
rect 30064 16612 32505 16640
rect 30064 16600 30070 16612
rect 32493 16609 32505 16612
rect 32539 16640 32551 16643
rect 32539 16612 32812 16640
rect 32539 16609 32551 16612
rect 32493 16603 32551 16609
rect 26510 16572 26516 16584
rect 24636 16544 26516 16572
rect 24636 16532 24642 16544
rect 26510 16532 26516 16544
rect 26568 16532 26574 16584
rect 26602 16532 26608 16584
rect 26660 16572 26666 16584
rect 26660 16544 31754 16572
rect 26660 16532 26666 16544
rect 20257 16507 20315 16513
rect 20257 16504 20269 16507
rect 18248 16476 19380 16504
rect 19444 16476 20269 16504
rect 18248 16445 18276 16476
rect 12437 16439 12495 16445
rect 12437 16436 12449 16439
rect 11756 16408 12449 16436
rect 11756 16396 11762 16408
rect 12437 16405 12449 16408
rect 12483 16405 12495 16439
rect 12437 16399 12495 16405
rect 13173 16439 13231 16445
rect 13173 16405 13185 16439
rect 13219 16405 13231 16439
rect 13173 16399 13231 16405
rect 18233 16439 18291 16445
rect 18233 16405 18245 16439
rect 18279 16405 18291 16439
rect 18233 16399 18291 16405
rect 18414 16396 18420 16448
rect 18472 16436 18478 16448
rect 18782 16436 18788 16448
rect 18472 16408 18788 16436
rect 18472 16396 18478 16408
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 19352 16436 19380 16476
rect 20257 16473 20269 16476
rect 20303 16473 20315 16507
rect 26050 16504 26056 16516
rect 20257 16467 20315 16473
rect 20364 16476 26056 16504
rect 20364 16436 20392 16476
rect 26050 16464 26056 16476
rect 26108 16464 26114 16516
rect 26228 16507 26286 16513
rect 26228 16473 26240 16507
rect 26274 16504 26286 16507
rect 27154 16504 27160 16516
rect 26274 16476 27160 16504
rect 26274 16473 26286 16476
rect 26228 16467 26286 16473
rect 27154 16464 27160 16476
rect 27212 16464 27218 16516
rect 31726 16504 31754 16544
rect 32125 16507 32183 16513
rect 32125 16504 32137 16507
rect 31726 16476 32137 16504
rect 32125 16473 32137 16476
rect 32171 16473 32183 16507
rect 32125 16467 32183 16473
rect 32309 16507 32367 16513
rect 32309 16473 32321 16507
rect 32355 16504 32367 16507
rect 32398 16504 32404 16516
rect 32355 16476 32404 16504
rect 32355 16473 32367 16476
rect 32309 16467 32367 16473
rect 19352 16408 20392 16436
rect 21910 16396 21916 16448
rect 21968 16436 21974 16448
rect 22189 16439 22247 16445
rect 22189 16436 22201 16439
rect 21968 16408 22201 16436
rect 21968 16396 21974 16408
rect 22189 16405 22201 16408
rect 22235 16405 22247 16439
rect 22189 16399 22247 16405
rect 24486 16396 24492 16448
rect 24544 16436 24550 16448
rect 26142 16436 26148 16448
rect 24544 16408 26148 16436
rect 24544 16396 24550 16408
rect 26142 16396 26148 16408
rect 26200 16396 26206 16448
rect 27246 16396 27252 16448
rect 27304 16436 27310 16448
rect 27341 16439 27399 16445
rect 27341 16436 27353 16439
rect 27304 16408 27353 16436
rect 27304 16396 27310 16408
rect 27341 16405 27353 16408
rect 27387 16405 27399 16439
rect 27341 16399 27399 16405
rect 27706 16396 27712 16448
rect 27764 16436 27770 16448
rect 27985 16439 28043 16445
rect 27985 16436 27997 16439
rect 27764 16408 27997 16436
rect 27764 16396 27770 16408
rect 27985 16405 27997 16408
rect 28031 16405 28043 16439
rect 27985 16399 28043 16405
rect 28350 16396 28356 16448
rect 28408 16396 28414 16448
rect 32140 16436 32168 16467
rect 32398 16464 32404 16476
rect 32456 16464 32462 16516
rect 32784 16504 32812 16612
rect 32858 16600 32864 16652
rect 32916 16640 32922 16652
rect 32953 16643 33011 16649
rect 32953 16640 32965 16643
rect 32916 16612 32965 16640
rect 32916 16600 32922 16612
rect 32953 16609 32965 16612
rect 32999 16609 33011 16643
rect 32953 16603 33011 16609
rect 36722 16600 36728 16652
rect 36780 16600 36786 16652
rect 36906 16600 36912 16652
rect 36964 16600 36970 16652
rect 37182 16600 37188 16652
rect 37240 16640 37246 16652
rect 37461 16643 37519 16649
rect 37461 16640 37473 16643
rect 37240 16612 37473 16640
rect 37240 16600 37246 16612
rect 37461 16609 37473 16612
rect 37507 16609 37519 16643
rect 37461 16603 37519 16609
rect 40034 16600 40040 16652
rect 40092 16640 40098 16652
rect 41509 16643 41567 16649
rect 41509 16640 41521 16643
rect 40092 16612 41521 16640
rect 40092 16600 40098 16612
rect 41509 16609 41521 16612
rect 41555 16609 41567 16643
rect 41509 16603 41567 16609
rect 41708 16640 41736 16680
rect 51534 16668 51540 16720
rect 51592 16708 51598 16720
rect 51592 16680 53604 16708
rect 51592 16668 51598 16680
rect 42794 16640 42800 16652
rect 41708 16612 42800 16640
rect 33226 16581 33232 16584
rect 33220 16572 33232 16581
rect 33187 16544 33232 16572
rect 33220 16535 33232 16544
rect 33226 16532 33232 16535
rect 33284 16532 33290 16584
rect 36538 16532 36544 16584
rect 36596 16572 36602 16584
rect 37200 16572 37228 16600
rect 36596 16544 37228 16572
rect 37728 16575 37786 16581
rect 36596 16532 36602 16544
rect 37728 16541 37740 16575
rect 37774 16572 37786 16575
rect 38286 16572 38292 16584
rect 37774 16544 38292 16572
rect 37774 16541 37786 16544
rect 37728 16535 37786 16541
rect 38286 16532 38292 16544
rect 38344 16532 38350 16584
rect 40678 16532 40684 16584
rect 40736 16532 40742 16584
rect 40846 16575 40904 16581
rect 40846 16541 40858 16575
rect 40892 16572 40904 16575
rect 40892 16541 40908 16572
rect 40846 16535 40908 16541
rect 35802 16504 35808 16516
rect 32784 16476 35808 16504
rect 35802 16464 35808 16476
rect 35860 16464 35866 16516
rect 36170 16464 36176 16516
rect 36228 16504 36234 16516
rect 36633 16507 36691 16513
rect 36633 16504 36645 16507
rect 36228 16476 36645 16504
rect 36228 16464 36234 16476
rect 36633 16473 36645 16476
rect 36679 16473 36691 16507
rect 36633 16467 36691 16473
rect 32490 16436 32496 16448
rect 32140 16408 32496 16436
rect 32490 16396 32496 16408
rect 32548 16396 32554 16448
rect 33962 16396 33968 16448
rect 34020 16436 34026 16448
rect 34333 16439 34391 16445
rect 34333 16436 34345 16439
rect 34020 16408 34345 16436
rect 34020 16396 34026 16408
rect 34333 16405 34345 16408
rect 34379 16405 34391 16439
rect 34333 16399 34391 16405
rect 36262 16396 36268 16448
rect 36320 16396 36326 16448
rect 38838 16396 38844 16448
rect 38896 16396 38902 16448
rect 40494 16396 40500 16448
rect 40552 16396 40558 16448
rect 40880 16436 40908 16535
rect 40954 16532 40960 16584
rect 41012 16532 41018 16584
rect 41046 16532 41052 16584
rect 41104 16532 41110 16584
rect 41708 16581 41736 16612
rect 42794 16600 42800 16612
rect 42852 16600 42858 16652
rect 44266 16600 44272 16652
rect 44324 16640 44330 16652
rect 45189 16643 45247 16649
rect 45189 16640 45201 16643
rect 44324 16612 45201 16640
rect 44324 16600 44330 16612
rect 45189 16609 45201 16612
rect 45235 16609 45247 16643
rect 45189 16603 45247 16609
rect 46750 16600 46756 16652
rect 46808 16640 46814 16652
rect 51445 16643 51503 16649
rect 51445 16640 51457 16643
rect 46808 16612 51457 16640
rect 46808 16600 46814 16612
rect 51445 16609 51457 16612
rect 51491 16640 51503 16643
rect 51810 16640 51816 16652
rect 51491 16612 51816 16640
rect 51491 16609 51503 16612
rect 51445 16603 51503 16609
rect 51810 16600 51816 16612
rect 51868 16600 51874 16652
rect 53576 16649 53604 16680
rect 53561 16643 53619 16649
rect 53561 16609 53573 16643
rect 53607 16609 53619 16643
rect 53561 16603 53619 16609
rect 41693 16575 41751 16581
rect 41693 16541 41705 16575
rect 41739 16541 41751 16575
rect 41693 16535 41751 16541
rect 41785 16575 41843 16581
rect 41785 16541 41797 16575
rect 41831 16541 41843 16575
rect 41785 16535 41843 16541
rect 41800 16504 41828 16535
rect 41966 16532 41972 16584
rect 42024 16532 42030 16584
rect 42058 16532 42064 16584
rect 42116 16532 42122 16584
rect 51626 16532 51632 16584
rect 51684 16532 51690 16584
rect 53828 16575 53886 16581
rect 53828 16541 53840 16575
rect 53874 16572 53886 16575
rect 54294 16572 54300 16584
rect 53874 16544 54300 16572
rect 53874 16541 53886 16544
rect 53828 16535 53886 16541
rect 54294 16532 54300 16544
rect 54352 16532 54358 16584
rect 57977 16575 58035 16581
rect 57977 16541 57989 16575
rect 58023 16572 58035 16575
rect 58802 16572 58808 16584
rect 58023 16544 58808 16572
rect 58023 16541 58035 16544
rect 57977 16535 58035 16541
rect 58802 16532 58808 16544
rect 58860 16532 58866 16584
rect 43438 16504 43444 16516
rect 41800 16476 43444 16504
rect 43438 16464 43444 16476
rect 43496 16464 43502 16516
rect 45456 16507 45514 16513
rect 45456 16473 45468 16507
rect 45502 16504 45514 16507
rect 46382 16504 46388 16516
rect 45502 16476 46388 16504
rect 45502 16473 45514 16476
rect 45456 16467 45514 16473
rect 46382 16464 46388 16476
rect 46440 16464 46446 16516
rect 47670 16464 47676 16516
rect 47728 16504 47734 16516
rect 52365 16507 52423 16513
rect 52365 16504 52377 16507
rect 47728 16476 52377 16504
rect 47728 16464 47734 16476
rect 52365 16473 52377 16476
rect 52411 16504 52423 16507
rect 56778 16504 56784 16516
rect 52411 16476 56784 16504
rect 52411 16473 52423 16476
rect 52365 16467 52423 16473
rect 56778 16464 56784 16476
rect 56836 16464 56842 16516
rect 57057 16507 57115 16513
rect 57057 16473 57069 16507
rect 57103 16504 57115 16507
rect 58986 16504 58992 16516
rect 57103 16476 58992 16504
rect 57103 16473 57115 16476
rect 57057 16467 57115 16473
rect 58986 16464 58992 16476
rect 59044 16464 59050 16516
rect 41690 16436 41696 16448
rect 40880 16408 41696 16436
rect 41690 16396 41696 16408
rect 41748 16396 41754 16448
rect 42702 16396 42708 16448
rect 42760 16436 42766 16448
rect 45554 16436 45560 16448
rect 42760 16408 45560 16436
rect 42760 16396 42766 16408
rect 45554 16396 45560 16408
rect 45612 16396 45618 16448
rect 46566 16396 46572 16448
rect 46624 16396 46630 16448
rect 51810 16396 51816 16448
rect 51868 16396 51874 16448
rect 52457 16439 52515 16445
rect 52457 16405 52469 16439
rect 52503 16436 52515 16439
rect 52914 16436 52920 16448
rect 52503 16408 52920 16436
rect 52503 16405 52515 16408
rect 52457 16399 52515 16405
rect 52914 16396 52920 16408
rect 52972 16396 52978 16448
rect 54941 16439 54999 16445
rect 54941 16405 54953 16439
rect 54987 16436 54999 16439
rect 55306 16436 55312 16448
rect 54987 16408 55312 16436
rect 54987 16405 54999 16408
rect 54941 16399 54999 16405
rect 55306 16396 55312 16408
rect 55364 16436 55370 16448
rect 56226 16436 56232 16448
rect 55364 16408 56232 16436
rect 55364 16396 55370 16408
rect 56226 16396 56232 16408
rect 56284 16396 56290 16448
rect 58066 16396 58072 16448
rect 58124 16396 58130 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 13538 16192 13544 16244
rect 13596 16192 13602 16244
rect 20346 16232 20352 16244
rect 18892 16204 20352 16232
rect 18892 16173 18920 16204
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 22189 16235 22247 16241
rect 22189 16232 22201 16235
rect 22066 16204 22201 16232
rect 18877 16167 18935 16173
rect 18877 16133 18889 16167
rect 18923 16133 18935 16167
rect 18877 16127 18935 16133
rect 18966 16124 18972 16176
rect 19024 16164 19030 16176
rect 19242 16164 19248 16176
rect 19024 16136 19248 16164
rect 19024 16124 19030 16136
rect 19242 16124 19248 16136
rect 19300 16124 19306 16176
rect 19429 16167 19487 16173
rect 19429 16133 19441 16167
rect 19475 16164 19487 16167
rect 20530 16164 20536 16176
rect 19475 16136 20536 16164
rect 19475 16133 19487 16136
rect 19429 16127 19487 16133
rect 20530 16124 20536 16136
rect 20588 16124 20594 16176
rect 22066 16164 22094 16204
rect 22189 16201 22201 16204
rect 22235 16201 22247 16235
rect 22189 16195 22247 16201
rect 22922 16192 22928 16244
rect 22980 16232 22986 16244
rect 23290 16232 23296 16244
rect 22980 16204 23296 16232
rect 22980 16192 22986 16204
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 24118 16192 24124 16244
rect 24176 16192 24182 16244
rect 24670 16192 24676 16244
rect 24728 16232 24734 16244
rect 26602 16232 26608 16244
rect 24728 16204 26608 16232
rect 24728 16192 24734 16204
rect 26602 16192 26608 16204
rect 26660 16192 26666 16244
rect 27154 16192 27160 16244
rect 27212 16192 27218 16244
rect 27522 16192 27528 16244
rect 27580 16192 27586 16244
rect 29457 16235 29515 16241
rect 29457 16201 29469 16235
rect 29503 16232 29515 16235
rect 31110 16232 31116 16244
rect 29503 16204 31116 16232
rect 29503 16201 29515 16204
rect 29457 16195 29515 16201
rect 31110 16192 31116 16204
rect 31168 16192 31174 16244
rect 31294 16192 31300 16244
rect 31352 16232 31358 16244
rect 36722 16232 36728 16244
rect 31352 16204 36728 16232
rect 31352 16192 31358 16204
rect 36722 16192 36728 16204
rect 36780 16192 36786 16244
rect 40034 16232 40040 16244
rect 37476 16204 40040 16232
rect 21100 16136 22094 16164
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 1854 16096 1860 16108
rect 1627 16068 1860 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 1854 16056 1860 16068
rect 1912 16096 1918 16108
rect 2317 16099 2375 16105
rect 2317 16096 2329 16099
rect 1912 16068 2329 16096
rect 1912 16056 1918 16068
rect 2317 16065 2329 16068
rect 2363 16065 2375 16099
rect 2317 16059 2375 16065
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 10318 16096 10324 16108
rect 9907 16068 10324 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 11698 16056 11704 16108
rect 11756 16056 11762 16108
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 11900 16068 12449 16096
rect 934 15988 940 16040
rect 992 16028 998 16040
rect 1765 16031 1823 16037
rect 1765 16028 1777 16031
rect 992 16000 1777 16028
rect 992 15988 998 16000
rect 1765 15997 1777 16000
rect 1811 15997 1823 16031
rect 1765 15991 1823 15997
rect 11900 15969 11928 16068
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 13354 16056 13360 16108
rect 13412 16096 13418 16108
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 13412 16068 13737 16096
rect 13412 16056 13418 16068
rect 13725 16065 13737 16068
rect 13771 16065 13783 16099
rect 13725 16059 13783 16065
rect 13814 16056 13820 16108
rect 13872 16056 13878 16108
rect 13906 16056 13912 16108
rect 13964 16056 13970 16108
rect 15746 16056 15752 16108
rect 15804 16056 15810 16108
rect 17034 16056 17040 16108
rect 17092 16056 17098 16108
rect 17304 16099 17362 16105
rect 17304 16065 17316 16099
rect 17350 16096 17362 16099
rect 17770 16096 17776 16108
rect 17350 16068 17776 16096
rect 17350 16065 17362 16068
rect 17304 16059 17362 16065
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 18690 16056 18696 16108
rect 18748 16096 18754 16108
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 18748 16068 19073 16096
rect 18748 16056 18754 16068
rect 19061 16065 19073 16068
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 19150 16056 19156 16108
rect 19208 16056 19214 16108
rect 21100 16105 21128 16136
rect 23566 16124 23572 16176
rect 23624 16164 23630 16176
rect 23624 16136 25360 16164
rect 23624 16124 23630 16136
rect 20349 16099 20407 16105
rect 20349 16065 20361 16099
rect 20395 16065 20407 16099
rect 20349 16059 20407 16065
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 16028 14059 16031
rect 14090 16028 14096 16040
rect 14047 16000 14096 16028
rect 14047 15997 14059 16000
rect 14001 15991 14059 15997
rect 14090 15988 14096 16000
rect 14148 15988 14154 16040
rect 20364 16028 20392 16059
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21968 16068 22017 16096
rect 21968 16056 21974 16068
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16096 23167 16099
rect 23198 16096 23204 16108
rect 23155 16068 23204 16096
rect 23155 16065 23167 16068
rect 23109 16059 23167 16065
rect 23198 16056 23204 16068
rect 23256 16056 23262 16108
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16096 23351 16099
rect 23842 16096 23848 16108
rect 23339 16068 23848 16096
rect 23339 16065 23351 16068
rect 23293 16059 23351 16065
rect 23842 16056 23848 16068
rect 23900 16056 23906 16108
rect 23937 16099 23995 16105
rect 23937 16065 23949 16099
rect 23983 16065 23995 16099
rect 23937 16059 23995 16065
rect 20364 16000 21312 16028
rect 21284 15969 21312 16000
rect 11885 15963 11943 15969
rect 11885 15929 11897 15963
rect 11931 15929 11943 15963
rect 11885 15923 11943 15929
rect 18417 15963 18475 15969
rect 18417 15929 18429 15963
rect 18463 15960 18475 15963
rect 21269 15963 21327 15969
rect 18463 15932 20944 15960
rect 18463 15929 18475 15932
rect 18417 15923 18475 15929
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 10045 15895 10103 15901
rect 10045 15892 10057 15895
rect 9732 15864 10057 15892
rect 9732 15852 9738 15864
rect 10045 15861 10057 15864
rect 10091 15861 10103 15895
rect 10045 15855 10103 15861
rect 12618 15852 12624 15904
rect 12676 15852 12682 15904
rect 15194 15852 15200 15904
rect 15252 15892 15258 15904
rect 15933 15895 15991 15901
rect 15933 15892 15945 15895
rect 15252 15864 15945 15892
rect 15252 15852 15258 15864
rect 15933 15861 15945 15864
rect 15979 15861 15991 15895
rect 15933 15855 15991 15861
rect 19886 15852 19892 15904
rect 19944 15892 19950 15904
rect 20533 15895 20591 15901
rect 20533 15892 20545 15895
rect 19944 15864 20545 15892
rect 19944 15852 19950 15864
rect 20533 15861 20545 15864
rect 20579 15861 20591 15895
rect 20916 15892 20944 15932
rect 21269 15929 21281 15963
rect 21315 15960 21327 15963
rect 23842 15960 23848 15972
rect 21315 15932 23848 15960
rect 21315 15929 21327 15932
rect 21269 15923 21327 15929
rect 23842 15920 23848 15932
rect 23900 15920 23906 15972
rect 23952 15960 23980 16059
rect 24302 16056 24308 16108
rect 24360 16096 24366 16108
rect 25041 16099 25099 16105
rect 25041 16096 25053 16099
rect 24360 16068 25053 16096
rect 24360 16056 24366 16068
rect 25041 16065 25053 16068
rect 25087 16096 25099 16099
rect 25130 16096 25136 16108
rect 25087 16068 25136 16096
rect 25087 16065 25099 16068
rect 25041 16059 25099 16065
rect 25130 16056 25136 16068
rect 25188 16056 25194 16108
rect 25332 16037 25360 16136
rect 25590 16124 25596 16176
rect 25648 16164 25654 16176
rect 25648 16136 28488 16164
rect 25648 16124 25654 16136
rect 26050 16056 26056 16108
rect 26108 16096 26114 16108
rect 26329 16099 26387 16105
rect 26329 16096 26341 16099
rect 26108 16068 26341 16096
rect 26108 16056 26114 16068
rect 26329 16065 26341 16068
rect 26375 16096 26387 16099
rect 28350 16096 28356 16108
rect 26375 16068 28356 16096
rect 26375 16065 26387 16068
rect 26329 16059 26387 16065
rect 28350 16056 28356 16068
rect 28408 16056 28414 16108
rect 28460 16096 28488 16136
rect 29546 16124 29552 16176
rect 29604 16124 29610 16176
rect 31202 16124 31208 16176
rect 31260 16124 31266 16176
rect 32306 16124 32312 16176
rect 32364 16164 32370 16176
rect 37476 16173 37504 16204
rect 40034 16192 40040 16204
rect 40092 16192 40098 16244
rect 40126 16192 40132 16244
rect 40184 16232 40190 16244
rect 40954 16232 40960 16244
rect 40184 16204 40960 16232
rect 40184 16192 40190 16204
rect 40954 16192 40960 16204
rect 41012 16192 41018 16244
rect 41046 16192 41052 16244
rect 41104 16232 41110 16244
rect 43165 16235 43223 16241
rect 43165 16232 43177 16235
rect 41104 16204 43177 16232
rect 41104 16192 41110 16204
rect 43165 16201 43177 16204
rect 43211 16201 43223 16235
rect 43165 16195 43223 16201
rect 45462 16192 45468 16244
rect 45520 16192 45526 16244
rect 46382 16192 46388 16244
rect 46440 16192 46446 16244
rect 46566 16192 46572 16244
rect 46624 16232 46630 16244
rect 46845 16235 46903 16241
rect 46845 16232 46857 16235
rect 46624 16204 46857 16232
rect 46624 16192 46630 16204
rect 46845 16201 46857 16204
rect 46891 16201 46903 16235
rect 46845 16195 46903 16201
rect 51074 16192 51080 16244
rect 51132 16232 51138 16244
rect 51132 16204 51304 16232
rect 51132 16192 51138 16204
rect 37461 16167 37519 16173
rect 32364 16136 32720 16164
rect 32364 16124 32370 16136
rect 31665 16099 31723 16105
rect 28460 16068 31616 16096
rect 25317 16031 25375 16037
rect 25317 15997 25329 16031
rect 25363 16028 25375 16031
rect 25682 16028 25688 16040
rect 25363 16000 25688 16028
rect 25363 15997 25375 16000
rect 25317 15991 25375 15997
rect 25682 15988 25688 16000
rect 25740 15988 25746 16040
rect 27246 15988 27252 16040
rect 27304 16028 27310 16040
rect 27617 16031 27675 16037
rect 27617 16028 27629 16031
rect 27304 16000 27629 16028
rect 27304 15988 27310 16000
rect 27617 15997 27629 16000
rect 27663 15997 27675 16031
rect 27617 15991 27675 15997
rect 27801 16031 27859 16037
rect 27801 15997 27813 16031
rect 27847 16028 27859 16031
rect 27890 16028 27896 16040
rect 27847 16000 27896 16028
rect 27847 15997 27859 16000
rect 27801 15991 27859 15997
rect 27890 15988 27896 16000
rect 27948 16028 27954 16040
rect 28166 16028 28172 16040
rect 27948 16000 28172 16028
rect 27948 15988 27954 16000
rect 28166 15988 28172 16000
rect 28224 16028 28230 16040
rect 29730 16028 29736 16040
rect 28224 16000 29736 16028
rect 28224 15988 28230 16000
rect 29730 15988 29736 16000
rect 29788 15988 29794 16040
rect 26513 15963 26571 15969
rect 26513 15960 26525 15963
rect 23952 15932 26525 15960
rect 26513 15929 26525 15932
rect 26559 15929 26571 15963
rect 26513 15923 26571 15929
rect 26602 15920 26608 15972
rect 26660 15960 26666 15972
rect 31294 15960 31300 15972
rect 26660 15932 31300 15960
rect 26660 15920 26666 15932
rect 31294 15920 31300 15932
rect 31352 15920 31358 15972
rect 31588 15960 31616 16068
rect 31665 16065 31677 16099
rect 31711 16096 31723 16099
rect 31754 16096 31760 16108
rect 31711 16068 31760 16096
rect 31711 16065 31723 16068
rect 31665 16059 31723 16065
rect 31754 16056 31760 16068
rect 31812 16056 31818 16108
rect 31846 16056 31852 16108
rect 31904 16096 31910 16108
rect 32692 16105 32720 16136
rect 37461 16133 37473 16167
rect 37507 16133 37519 16167
rect 37461 16127 37519 16133
rect 38473 16167 38531 16173
rect 38473 16133 38485 16167
rect 38519 16164 38531 16167
rect 40494 16164 40500 16176
rect 38519 16136 40500 16164
rect 38519 16133 38531 16136
rect 38473 16127 38531 16133
rect 40494 16124 40500 16136
rect 40552 16124 40558 16176
rect 41782 16124 41788 16176
rect 41840 16164 41846 16176
rect 42702 16164 42708 16176
rect 41840 16136 42708 16164
rect 41840 16124 41846 16136
rect 42702 16124 42708 16136
rect 42760 16124 42766 16176
rect 42889 16167 42947 16173
rect 42889 16133 42901 16167
rect 42935 16164 42947 16167
rect 43070 16164 43076 16176
rect 42935 16136 43076 16164
rect 42935 16133 42947 16136
rect 42889 16127 42947 16133
rect 43070 16124 43076 16136
rect 43128 16124 43134 16176
rect 46753 16167 46811 16173
rect 46753 16133 46765 16167
rect 46799 16164 46811 16167
rect 51166 16164 51172 16176
rect 46799 16136 51172 16164
rect 46799 16133 46811 16136
rect 46753 16127 46811 16133
rect 51166 16124 51172 16136
rect 51224 16124 51230 16176
rect 51276 16173 51304 16204
rect 51626 16192 51632 16244
rect 51684 16192 51690 16244
rect 53009 16235 53067 16241
rect 53009 16201 53021 16235
rect 53055 16232 53067 16235
rect 53834 16232 53840 16244
rect 53055 16204 53840 16232
rect 53055 16201 53067 16204
rect 53009 16195 53067 16201
rect 51261 16167 51319 16173
rect 51261 16133 51273 16167
rect 51307 16164 51319 16167
rect 51534 16164 51540 16176
rect 51307 16136 51540 16164
rect 51307 16133 51319 16136
rect 51261 16127 51319 16133
rect 51534 16124 51540 16136
rect 51592 16124 51598 16176
rect 53024 16164 53052 16195
rect 53834 16192 53840 16204
rect 53892 16192 53898 16244
rect 54110 16192 54116 16244
rect 54168 16232 54174 16244
rect 54205 16235 54263 16241
rect 54205 16232 54217 16235
rect 54168 16204 54217 16232
rect 54168 16192 54174 16204
rect 54205 16201 54217 16204
rect 54251 16201 54263 16235
rect 54205 16195 54263 16201
rect 52104 16136 53052 16164
rect 53929 16167 53987 16173
rect 32585 16099 32643 16105
rect 32585 16096 32597 16099
rect 31904 16068 32597 16096
rect 31904 16056 31910 16068
rect 32585 16065 32597 16068
rect 32631 16065 32643 16099
rect 32585 16059 32643 16065
rect 32677 16099 32735 16105
rect 32677 16065 32689 16099
rect 32723 16065 32735 16099
rect 32677 16059 32735 16065
rect 32861 16099 32919 16105
rect 32861 16065 32873 16099
rect 32907 16065 32919 16099
rect 32861 16059 32919 16065
rect 32953 16102 33011 16105
rect 32953 16099 33088 16102
rect 32953 16065 32965 16099
rect 32999 16074 33088 16099
rect 32999 16065 33011 16074
rect 32953 16059 33011 16065
rect 32876 15960 32904 16059
rect 33060 16028 33088 16074
rect 35802 16056 35808 16108
rect 35860 16096 35866 16108
rect 37645 16099 37703 16105
rect 37645 16096 37657 16099
rect 35860 16068 37657 16096
rect 35860 16056 35866 16068
rect 37645 16065 37657 16068
rect 37691 16096 37703 16099
rect 38657 16099 38715 16105
rect 38657 16096 38669 16099
rect 37691 16068 38669 16096
rect 37691 16065 37703 16068
rect 37645 16059 37703 16065
rect 38657 16065 38669 16068
rect 38703 16065 38715 16099
rect 38657 16059 38715 16065
rect 41509 16099 41567 16105
rect 41509 16065 41521 16099
rect 41555 16096 41567 16099
rect 41690 16096 41696 16108
rect 41555 16068 41696 16096
rect 41555 16065 41567 16068
rect 41509 16059 41567 16065
rect 41690 16056 41696 16068
rect 41748 16056 41754 16108
rect 41877 16099 41935 16105
rect 41877 16065 41889 16099
rect 41923 16096 41935 16099
rect 42058 16096 42064 16108
rect 41923 16068 42064 16096
rect 41923 16065 41935 16068
rect 41877 16059 41935 16065
rect 42058 16056 42064 16068
rect 42116 16056 42122 16108
rect 42426 16056 42432 16108
rect 42484 16096 42490 16108
rect 42613 16099 42671 16105
rect 42613 16096 42625 16099
rect 42484 16068 42625 16096
rect 42484 16056 42490 16068
rect 42613 16065 42625 16068
rect 42659 16065 42671 16099
rect 42613 16059 42671 16065
rect 42797 16099 42855 16105
rect 42797 16065 42809 16099
rect 42843 16065 42855 16099
rect 42797 16059 42855 16065
rect 37550 16028 37556 16040
rect 33060 16000 37556 16028
rect 37550 15988 37556 16000
rect 37608 15988 37614 16040
rect 41598 15988 41604 16040
rect 41656 15988 41662 16040
rect 41969 16031 42027 16037
rect 41969 15997 41981 16031
rect 42015 16028 42027 16031
rect 42812 16028 42840 16059
rect 42978 16056 42984 16108
rect 43036 16056 43042 16108
rect 44174 16056 44180 16108
rect 44232 16056 44238 16108
rect 47854 16056 47860 16108
rect 47912 16096 47918 16108
rect 48021 16099 48079 16105
rect 48021 16096 48033 16099
rect 47912 16068 48033 16096
rect 47912 16056 47918 16068
rect 48021 16065 48033 16068
rect 48067 16065 48079 16099
rect 48021 16059 48079 16065
rect 50706 16056 50712 16108
rect 50764 16096 50770 16108
rect 51077 16099 51135 16105
rect 51077 16096 51089 16099
rect 50764 16068 51089 16096
rect 50764 16056 50770 16068
rect 51077 16065 51089 16068
rect 51123 16065 51135 16099
rect 51077 16059 51135 16065
rect 51350 16056 51356 16108
rect 51408 16056 51414 16108
rect 52104 16105 52132 16136
rect 53929 16133 53941 16167
rect 53975 16164 53987 16167
rect 55306 16164 55312 16176
rect 53975 16136 55312 16164
rect 53975 16133 53987 16136
rect 53929 16127 53987 16133
rect 55306 16124 55312 16136
rect 55364 16124 55370 16176
rect 51445 16099 51503 16105
rect 51445 16065 51457 16099
rect 51491 16065 51503 16099
rect 51445 16059 51503 16065
rect 52089 16099 52147 16105
rect 52089 16065 52101 16099
rect 52135 16065 52147 16099
rect 52089 16059 52147 16065
rect 42886 16028 42892 16040
rect 42015 16000 42892 16028
rect 42015 15997 42027 16000
rect 41969 15991 42027 15997
rect 32950 15960 32956 15972
rect 31588 15932 32536 15960
rect 32876 15932 32956 15960
rect 21910 15892 21916 15904
rect 20916 15864 21916 15892
rect 20533 15855 20591 15861
rect 21910 15852 21916 15864
rect 21968 15852 21974 15904
rect 23106 15852 23112 15904
rect 23164 15892 23170 15904
rect 23477 15895 23535 15901
rect 23477 15892 23489 15895
rect 23164 15864 23489 15892
rect 23164 15852 23170 15864
rect 23477 15861 23489 15864
rect 23523 15861 23535 15895
rect 23477 15855 23535 15861
rect 23658 15852 23664 15904
rect 23716 15892 23722 15904
rect 23934 15892 23940 15904
rect 23716 15864 23940 15892
rect 23716 15852 23722 15864
rect 23934 15852 23940 15864
rect 23992 15892 23998 15904
rect 24670 15892 24676 15904
rect 23992 15864 24676 15892
rect 23992 15852 23998 15864
rect 24670 15852 24676 15864
rect 24728 15852 24734 15904
rect 28718 15852 28724 15904
rect 28776 15892 28782 15904
rect 29089 15895 29147 15901
rect 29089 15892 29101 15895
rect 28776 15864 29101 15892
rect 28776 15852 28782 15864
rect 29089 15861 29101 15864
rect 29135 15861 29147 15895
rect 29089 15855 29147 15861
rect 32214 15852 32220 15904
rect 32272 15892 32278 15904
rect 32401 15895 32459 15901
rect 32401 15892 32413 15895
rect 32272 15864 32413 15892
rect 32272 15852 32278 15864
rect 32401 15861 32413 15864
rect 32447 15861 32459 15895
rect 32508 15892 32536 15932
rect 32950 15920 32956 15932
rect 33008 15920 33014 15972
rect 40862 15960 40868 15972
rect 33060 15932 40868 15960
rect 33060 15892 33088 15932
rect 40862 15920 40868 15932
rect 40920 15960 40926 15972
rect 40957 15963 41015 15969
rect 40957 15960 40969 15963
rect 40920 15932 40969 15960
rect 40920 15920 40926 15932
rect 40957 15929 40969 15932
rect 41003 15929 41015 15963
rect 40957 15923 41015 15929
rect 41506 15920 41512 15972
rect 41564 15960 41570 15972
rect 41984 15960 42012 15991
rect 42886 15988 42892 16000
rect 42944 15988 42950 16040
rect 46937 16031 46995 16037
rect 46937 15997 46949 16031
rect 46983 15997 46995 16031
rect 46937 15991 46995 15997
rect 46952 15960 46980 15991
rect 47762 15988 47768 16040
rect 47820 15988 47826 16040
rect 50982 15988 50988 16040
rect 51040 16028 51046 16040
rect 51460 16028 51488 16059
rect 52914 16056 52920 16108
rect 52972 16056 52978 16108
rect 53098 16056 53104 16108
rect 53156 16056 53162 16108
rect 53190 16056 53196 16108
rect 53248 16096 53254 16108
rect 53653 16099 53711 16105
rect 53653 16096 53665 16099
rect 53248 16068 53665 16096
rect 53248 16056 53254 16068
rect 53653 16065 53665 16068
rect 53699 16065 53711 16099
rect 53653 16059 53711 16065
rect 53834 16056 53840 16108
rect 53892 16056 53898 16108
rect 54021 16099 54079 16105
rect 54021 16065 54033 16099
rect 54067 16096 54079 16099
rect 54938 16096 54944 16108
rect 54067 16068 54944 16096
rect 54067 16065 54079 16068
rect 54021 16059 54079 16065
rect 54036 16028 54064 16059
rect 54938 16056 54944 16068
rect 54996 16056 55002 16108
rect 51040 16000 54064 16028
rect 51040 15988 51046 16000
rect 41564 15932 42012 15960
rect 46860 15932 46980 15960
rect 41564 15920 41570 15932
rect 46860 15904 46888 15932
rect 32508 15864 33088 15892
rect 32401 15855 32459 15861
rect 36446 15852 36452 15904
rect 36504 15892 36510 15904
rect 37090 15892 37096 15904
rect 36504 15864 37096 15892
rect 36504 15852 36510 15864
rect 37090 15852 37096 15864
rect 37148 15892 37154 15904
rect 37737 15895 37795 15901
rect 37737 15892 37749 15895
rect 37148 15864 37749 15892
rect 37148 15852 37154 15864
rect 37737 15861 37749 15864
rect 37783 15861 37795 15895
rect 37737 15855 37795 15861
rect 38194 15852 38200 15904
rect 38252 15892 38258 15904
rect 38749 15895 38807 15901
rect 38749 15892 38761 15895
rect 38252 15864 38761 15892
rect 38252 15852 38258 15864
rect 38749 15861 38761 15864
rect 38795 15861 38807 15895
rect 38749 15855 38807 15861
rect 46842 15852 46848 15904
rect 46900 15852 46906 15904
rect 48130 15852 48136 15904
rect 48188 15892 48194 15904
rect 49145 15895 49203 15901
rect 49145 15892 49157 15895
rect 48188 15864 49157 15892
rect 48188 15852 48194 15864
rect 49145 15861 49157 15864
rect 49191 15861 49203 15895
rect 49145 15855 49203 15861
rect 50706 15852 50712 15904
rect 50764 15852 50770 15904
rect 51534 15852 51540 15904
rect 51592 15892 51598 15904
rect 52273 15895 52331 15901
rect 52273 15892 52285 15895
rect 51592 15864 52285 15892
rect 51592 15852 51598 15864
rect 52273 15861 52285 15864
rect 52319 15892 52331 15895
rect 53834 15892 53840 15904
rect 52319 15864 53840 15892
rect 52319 15861 52331 15864
rect 52273 15855 52331 15861
rect 53834 15852 53840 15864
rect 53892 15892 53898 15904
rect 55122 15892 55128 15904
rect 53892 15864 55128 15892
rect 53892 15852 53898 15864
rect 55122 15852 55128 15864
rect 55180 15852 55186 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 10318 15648 10324 15700
rect 10376 15648 10382 15700
rect 10410 15648 10416 15700
rect 10468 15688 10474 15700
rect 13081 15691 13139 15697
rect 13081 15688 13093 15691
rect 10468 15660 13093 15688
rect 10468 15648 10474 15660
rect 13081 15657 13093 15660
rect 13127 15657 13139 15691
rect 13081 15651 13139 15657
rect 17770 15648 17776 15700
rect 17828 15648 17834 15700
rect 21729 15691 21787 15697
rect 21729 15688 21741 15691
rect 18064 15660 21741 15688
rect 12437 15623 12495 15629
rect 12437 15589 12449 15623
rect 12483 15620 12495 15623
rect 17126 15620 17132 15632
rect 12483 15592 17132 15620
rect 12483 15589 12495 15592
rect 12437 15583 12495 15589
rect 17126 15580 17132 15592
rect 17184 15580 17190 15632
rect 11054 15512 11060 15564
rect 11112 15512 11118 15564
rect 12066 15512 12072 15564
rect 12124 15552 12130 15564
rect 13449 15555 13507 15561
rect 13449 15552 13461 15555
rect 12124 15524 13461 15552
rect 12124 15512 12130 15524
rect 13449 15521 13461 15524
rect 13495 15552 13507 15555
rect 13814 15552 13820 15564
rect 13495 15524 13820 15552
rect 13495 15521 13507 15524
rect 13449 15515 13507 15521
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 18064 15552 18092 15660
rect 21729 15657 21741 15660
rect 21775 15657 21787 15691
rect 21729 15651 21787 15657
rect 23293 15691 23351 15697
rect 23293 15657 23305 15691
rect 23339 15688 23351 15691
rect 23339 15660 41414 15688
rect 23339 15657 23351 15660
rect 23293 15651 23351 15657
rect 18693 15623 18751 15629
rect 18693 15589 18705 15623
rect 18739 15620 18751 15623
rect 20625 15623 20683 15629
rect 20625 15620 20637 15623
rect 18739 15592 20637 15620
rect 18739 15589 18751 15592
rect 18693 15583 18751 15589
rect 20625 15589 20637 15592
rect 20671 15589 20683 15623
rect 20625 15583 20683 15589
rect 22830 15580 22836 15632
rect 22888 15620 22894 15632
rect 23382 15620 23388 15632
rect 22888 15592 23388 15620
rect 22888 15580 22894 15592
rect 23382 15580 23388 15592
rect 23440 15620 23446 15632
rect 23937 15623 23995 15629
rect 23937 15620 23949 15623
rect 23440 15592 23949 15620
rect 23440 15580 23446 15592
rect 23937 15589 23949 15592
rect 23983 15589 23995 15623
rect 23937 15583 23995 15589
rect 24026 15580 24032 15632
rect 24084 15620 24090 15632
rect 24302 15620 24308 15632
rect 24084 15592 24308 15620
rect 24084 15580 24090 15592
rect 24302 15580 24308 15592
rect 24360 15580 24366 15632
rect 28534 15580 28540 15632
rect 28592 15620 28598 15632
rect 36446 15620 36452 15632
rect 28592 15592 36452 15620
rect 28592 15580 28598 15592
rect 36446 15580 36452 15592
rect 36504 15580 36510 15632
rect 41386 15620 41414 15660
rect 41690 15648 41696 15700
rect 41748 15648 41754 15700
rect 42058 15648 42064 15700
rect 42116 15688 42122 15700
rect 45278 15688 45284 15700
rect 42116 15660 45284 15688
rect 42116 15648 42122 15660
rect 45278 15648 45284 15660
rect 45336 15648 45342 15700
rect 48133 15691 48191 15697
rect 48133 15657 48145 15691
rect 48179 15688 48191 15691
rect 48222 15688 48228 15700
rect 48179 15660 48228 15688
rect 48179 15657 48191 15660
rect 48133 15651 48191 15657
rect 48222 15648 48228 15660
rect 48280 15648 48286 15700
rect 51350 15648 51356 15700
rect 51408 15688 51414 15700
rect 51408 15660 52960 15688
rect 51408 15648 51414 15660
rect 52932 15629 52960 15660
rect 53098 15648 53104 15700
rect 53156 15688 53162 15700
rect 58526 15688 58532 15700
rect 53156 15660 58532 15688
rect 53156 15648 53162 15660
rect 58526 15648 58532 15660
rect 58584 15648 58590 15700
rect 52917 15623 52975 15629
rect 41386 15592 48314 15620
rect 15304 15524 16712 15552
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 9953 15487 10011 15493
rect 9953 15484 9965 15487
rect 9824 15456 9965 15484
rect 9824 15444 9830 15456
rect 9953 15453 9965 15456
rect 9999 15453 10011 15487
rect 9953 15447 10011 15453
rect 10134 15444 10140 15496
rect 10192 15444 10198 15496
rect 13262 15444 13268 15496
rect 13320 15444 13326 15496
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15484 13599 15487
rect 13906 15484 13912 15496
rect 13587 15456 13912 15484
rect 13587 15453 13599 15456
rect 13541 15447 13599 15453
rect 11324 15419 11382 15425
rect 11324 15385 11336 15419
rect 11370 15416 11382 15419
rect 12618 15416 12624 15428
rect 11370 15388 12624 15416
rect 11370 15385 11382 15388
rect 11324 15379 11382 15385
rect 12618 15376 12624 15388
rect 12676 15376 12682 15428
rect 13372 15416 13400 15447
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 14274 15444 14280 15496
rect 14332 15444 14338 15496
rect 15304 15493 15332 15524
rect 15289 15487 15347 15493
rect 15289 15453 15301 15487
rect 15335 15453 15347 15487
rect 15289 15447 15347 15453
rect 16114 15444 16120 15496
rect 16172 15444 16178 15496
rect 16482 15416 16488 15428
rect 13372 15388 16488 15416
rect 16482 15376 16488 15388
rect 16540 15376 16546 15428
rect 16684 15416 16712 15524
rect 16868 15524 18092 15552
rect 18785 15555 18843 15561
rect 16868 15493 16896 15524
rect 18785 15521 18797 15555
rect 18831 15521 18843 15555
rect 18785 15515 18843 15521
rect 16853 15487 16911 15493
rect 16853 15453 16865 15487
rect 16899 15453 16911 15487
rect 16853 15447 16911 15453
rect 17589 15487 17647 15493
rect 17589 15453 17601 15487
rect 17635 15484 17647 15487
rect 18800 15484 18828 15515
rect 19150 15512 19156 15564
rect 19208 15552 19214 15564
rect 19613 15555 19671 15561
rect 19613 15552 19625 15555
rect 19208 15524 19625 15552
rect 19208 15512 19214 15524
rect 19613 15521 19625 15524
rect 19659 15521 19671 15555
rect 19613 15515 19671 15521
rect 19886 15512 19892 15564
rect 19944 15512 19950 15564
rect 24118 15552 24124 15564
rect 22756 15524 24124 15552
rect 17635 15456 18828 15484
rect 17635 15453 17647 15456
rect 17589 15447 17647 15453
rect 18874 15444 18880 15496
rect 18932 15484 18938 15496
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 18932 15456 19717 15484
rect 18932 15444 18938 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15484 19855 15487
rect 20254 15484 20260 15496
rect 19843 15456 20260 15484
rect 19843 15453 19855 15456
rect 19797 15447 19855 15453
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 20438 15444 20444 15496
rect 20496 15444 20502 15496
rect 22756 15493 22784 15524
rect 24118 15512 24124 15524
rect 24176 15512 24182 15564
rect 25608 15524 27660 15552
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 22741 15487 22799 15493
rect 22741 15453 22753 15487
rect 22787 15453 22799 15487
rect 22741 15447 22799 15453
rect 23161 15487 23219 15493
rect 23161 15453 23173 15487
rect 23207 15484 23219 15487
rect 23207 15456 23796 15484
rect 23207 15453 23219 15456
rect 23161 15447 23219 15453
rect 16684 15388 16896 15416
rect 14458 15308 14464 15360
rect 14516 15308 14522 15360
rect 15470 15308 15476 15360
rect 15528 15308 15534 15360
rect 16301 15351 16359 15357
rect 16301 15317 16313 15351
rect 16347 15348 16359 15351
rect 16758 15348 16764 15360
rect 16347 15320 16764 15348
rect 16347 15317 16359 15320
rect 16301 15311 16359 15317
rect 16758 15308 16764 15320
rect 16816 15308 16822 15360
rect 16868 15348 16896 15388
rect 17126 15376 17132 15428
rect 17184 15416 17190 15428
rect 18325 15419 18383 15425
rect 17184 15388 18092 15416
rect 17184 15376 17190 15388
rect 17037 15351 17095 15357
rect 17037 15348 17049 15351
rect 16868 15320 17049 15348
rect 17037 15317 17049 15320
rect 17083 15348 17095 15351
rect 17954 15348 17960 15360
rect 17083 15320 17960 15348
rect 17083 15317 17095 15320
rect 17037 15311 17095 15317
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 18064 15348 18092 15388
rect 18325 15385 18337 15419
rect 18371 15416 18383 15419
rect 19242 15416 19248 15428
rect 18371 15388 19248 15416
rect 18371 15385 18383 15388
rect 18325 15379 18383 15385
rect 19242 15376 19248 15388
rect 19300 15376 19306 15428
rect 21560 15416 21588 15447
rect 19352 15388 21588 15416
rect 19352 15348 19380 15388
rect 18064 15320 19380 15348
rect 19426 15308 19432 15360
rect 19484 15308 19490 15360
rect 21560 15348 21588 15388
rect 21726 15376 21732 15428
rect 21784 15416 21790 15428
rect 22925 15419 22983 15425
rect 22925 15416 22937 15419
rect 21784 15388 22937 15416
rect 21784 15376 21790 15388
rect 22925 15385 22937 15388
rect 22971 15385 22983 15419
rect 22925 15379 22983 15385
rect 23014 15376 23020 15428
rect 23072 15376 23078 15428
rect 23768 15416 23796 15456
rect 23842 15444 23848 15496
rect 23900 15444 23906 15496
rect 24578 15444 24584 15496
rect 24636 15444 24642 15496
rect 24670 15444 24676 15496
rect 24728 15484 24734 15496
rect 25608 15484 25636 15524
rect 24728 15456 25636 15484
rect 24728 15444 24734 15456
rect 25682 15444 25688 15496
rect 25740 15484 25746 15496
rect 26513 15487 26571 15493
rect 26513 15484 26525 15487
rect 25740 15456 26525 15484
rect 25740 15444 25746 15456
rect 26513 15453 26525 15456
rect 26559 15453 26571 15487
rect 26513 15447 26571 15453
rect 26694 15444 26700 15496
rect 26752 15444 26758 15496
rect 27522 15444 27528 15496
rect 27580 15444 27586 15496
rect 27632 15484 27660 15524
rect 31202 15512 31208 15564
rect 31260 15552 31266 15564
rect 34054 15552 34060 15564
rect 31260 15524 34060 15552
rect 31260 15512 31266 15524
rect 34054 15512 34060 15524
rect 34112 15512 34118 15564
rect 35342 15512 35348 15564
rect 35400 15552 35406 15564
rect 35437 15555 35495 15561
rect 35437 15552 35449 15555
rect 35400 15524 35449 15552
rect 35400 15512 35406 15524
rect 35437 15521 35449 15524
rect 35483 15521 35495 15555
rect 35437 15515 35495 15521
rect 36262 15512 36268 15564
rect 36320 15552 36326 15564
rect 36320 15524 36676 15552
rect 36320 15512 36326 15524
rect 27632 15456 28028 15484
rect 24210 15416 24216 15428
rect 23768 15388 24216 15416
rect 24210 15376 24216 15388
rect 24268 15376 24274 15428
rect 24848 15419 24906 15425
rect 24848 15385 24860 15419
rect 24894 15416 24906 15419
rect 26881 15419 26939 15425
rect 26881 15416 26893 15419
rect 24894 15388 26893 15416
rect 24894 15385 24906 15388
rect 24848 15379 24906 15385
rect 26881 15385 26893 15388
rect 26927 15385 26939 15419
rect 26881 15379 26939 15385
rect 27792 15419 27850 15425
rect 27792 15385 27804 15419
rect 27838 15416 27850 15419
rect 27890 15416 27896 15428
rect 27838 15388 27896 15416
rect 27838 15385 27850 15388
rect 27792 15379 27850 15385
rect 27890 15376 27896 15388
rect 27948 15376 27954 15428
rect 28000 15416 28028 15456
rect 31754 15444 31760 15496
rect 31812 15484 31818 15496
rect 32674 15484 32680 15496
rect 31812 15456 32680 15484
rect 31812 15444 31818 15456
rect 32674 15444 32680 15456
rect 32732 15444 32738 15496
rect 35253 15487 35311 15493
rect 35253 15453 35265 15487
rect 35299 15484 35311 15487
rect 35618 15484 35624 15496
rect 35299 15456 35624 15484
rect 35299 15453 35311 15456
rect 35253 15447 35311 15453
rect 35618 15444 35624 15456
rect 35676 15444 35682 15496
rect 36538 15444 36544 15496
rect 36596 15444 36602 15496
rect 36648 15484 36676 15524
rect 37550 15512 37556 15564
rect 37608 15552 37614 15564
rect 42058 15552 42064 15564
rect 37608 15524 42064 15552
rect 37608 15512 37614 15524
rect 42058 15512 42064 15524
rect 42116 15512 42122 15564
rect 48286 15552 48314 15592
rect 52917 15589 52929 15623
rect 52963 15620 52975 15623
rect 52963 15592 57928 15620
rect 52963 15589 52975 15592
rect 52917 15583 52975 15589
rect 48286 15524 51672 15552
rect 36797 15487 36855 15493
rect 36797 15484 36809 15487
rect 36648 15456 36809 15484
rect 36797 15453 36809 15456
rect 36843 15453 36855 15487
rect 36797 15447 36855 15453
rect 41046 15444 41052 15496
rect 41104 15444 41110 15496
rect 41230 15493 41236 15496
rect 41197 15487 41236 15493
rect 41197 15453 41209 15487
rect 41197 15447 41236 15453
rect 41230 15444 41236 15447
rect 41288 15444 41294 15496
rect 41322 15444 41328 15496
rect 41380 15444 41386 15496
rect 41414 15444 41420 15496
rect 41472 15444 41478 15496
rect 41598 15493 41604 15496
rect 41555 15487 41604 15493
rect 41555 15453 41567 15487
rect 41601 15453 41604 15487
rect 41555 15447 41604 15453
rect 41598 15444 41604 15447
rect 41656 15484 41662 15496
rect 42978 15484 42984 15496
rect 41656 15456 42984 15484
rect 41656 15444 41662 15456
rect 42978 15444 42984 15456
rect 43036 15444 43042 15496
rect 48222 15444 48228 15496
rect 48280 15484 48286 15496
rect 51442 15484 51448 15496
rect 48280 15456 51448 15484
rect 48280 15444 48286 15456
rect 51442 15444 51448 15456
rect 51500 15484 51506 15496
rect 51537 15487 51595 15493
rect 51537 15484 51549 15487
rect 51500 15456 51549 15484
rect 51500 15444 51506 15456
rect 51537 15453 51549 15456
rect 51583 15453 51595 15487
rect 51644 15484 51672 15524
rect 53190 15484 53196 15496
rect 51644 15456 53196 15484
rect 51537 15447 51595 15453
rect 53190 15444 53196 15456
rect 53248 15444 53254 15496
rect 57900 15493 57928 15592
rect 57885 15487 57943 15493
rect 57885 15453 57897 15487
rect 57931 15453 57943 15487
rect 57885 15447 57943 15453
rect 28000 15388 38056 15416
rect 24946 15348 24952 15360
rect 21560 15320 24952 15348
rect 24946 15308 24952 15320
rect 25004 15348 25010 15360
rect 25961 15351 26019 15357
rect 25961 15348 25973 15351
rect 25004 15320 25973 15348
rect 25004 15308 25010 15320
rect 25961 15317 25973 15320
rect 26007 15317 26019 15351
rect 25961 15311 26019 15317
rect 28350 15308 28356 15360
rect 28408 15348 28414 15360
rect 28905 15351 28963 15357
rect 28905 15348 28917 15351
rect 28408 15320 28917 15348
rect 28408 15308 28414 15320
rect 28905 15317 28917 15320
rect 28951 15317 28963 15351
rect 28905 15311 28963 15317
rect 34698 15308 34704 15360
rect 34756 15348 34762 15360
rect 34885 15351 34943 15357
rect 34885 15348 34897 15351
rect 34756 15320 34897 15348
rect 34756 15308 34762 15320
rect 34885 15317 34897 15320
rect 34931 15317 34943 15351
rect 34885 15311 34943 15317
rect 35345 15351 35403 15357
rect 35345 15317 35357 15351
rect 35391 15348 35403 15351
rect 35618 15348 35624 15360
rect 35391 15320 35624 15348
rect 35391 15317 35403 15320
rect 35345 15311 35403 15317
rect 35618 15308 35624 15320
rect 35676 15308 35682 15360
rect 36722 15308 36728 15360
rect 36780 15348 36786 15360
rect 37921 15351 37979 15357
rect 37921 15348 37933 15351
rect 36780 15320 37933 15348
rect 36780 15308 36786 15320
rect 37921 15317 37933 15320
rect 37967 15317 37979 15351
rect 38028 15348 38056 15388
rect 44174 15376 44180 15428
rect 44232 15416 44238 15428
rect 51810 15425 51816 15428
rect 46845 15419 46903 15425
rect 46845 15416 46857 15419
rect 44232 15388 46857 15416
rect 44232 15376 44238 15388
rect 46845 15385 46857 15388
rect 46891 15385 46903 15419
rect 51804 15416 51816 15425
rect 51771 15388 51816 15416
rect 46845 15379 46903 15385
rect 51804 15379 51816 15388
rect 51810 15376 51816 15379
rect 51868 15376 51874 15428
rect 58158 15376 58164 15428
rect 58216 15376 58222 15428
rect 50706 15348 50712 15360
rect 38028 15320 50712 15348
rect 37921 15311 37979 15317
rect 50706 15308 50712 15320
rect 50764 15308 50770 15360
rect 51166 15308 51172 15360
rect 51224 15348 51230 15360
rect 58618 15348 58624 15360
rect 51224 15320 58624 15348
rect 51224 15308 51230 15320
rect 58618 15308 58624 15320
rect 58676 15308 58682 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 15470 15144 15476 15156
rect 11900 15116 15476 15144
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 15008 1639 15011
rect 1627 14980 2774 15008
rect 1627 14977 1639 14980
rect 1581 14971 1639 14977
rect 934 14900 940 14952
rect 992 14940 998 14952
rect 1765 14943 1823 14949
rect 1765 14940 1777 14943
rect 992 14912 1777 14940
rect 992 14900 998 14912
rect 1765 14909 1777 14912
rect 1811 14909 1823 14943
rect 1765 14903 1823 14909
rect 2746 14804 2774 14980
rect 9306 14968 9312 15020
rect 9364 15008 9370 15020
rect 9401 15011 9459 15017
rect 9401 15008 9413 15011
rect 9364 14980 9413 15008
rect 9364 14968 9370 14980
rect 9401 14977 9413 14980
rect 9447 15008 9459 15011
rect 11054 15008 11060 15020
rect 9447 14980 11060 15008
rect 9447 14977 9459 14980
rect 9401 14971 9459 14977
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 11900 15017 11928 15116
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 16482 15104 16488 15156
rect 16540 15144 16546 15156
rect 16540 15116 18092 15144
rect 16540 15104 16546 15116
rect 17957 15079 18015 15085
rect 17957 15076 17969 15079
rect 14384 15048 17969 15076
rect 14384 15020 14412 15048
rect 17957 15045 17969 15048
rect 18003 15045 18015 15079
rect 17957 15039 18015 15045
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 14977 11943 15011
rect 12618 15008 12624 15020
rect 11885 14971 11943 14977
rect 11992 14980 12624 15008
rect 9674 14900 9680 14952
rect 9732 14900 9738 14952
rect 11072 14872 11100 14968
rect 11992 14949 12020 14980
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 12710 14968 12716 15020
rect 12768 14968 12774 15020
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 15008 13507 15011
rect 14182 15008 14188 15020
rect 13495 14980 14188 15008
rect 13495 14977 13507 14980
rect 13449 14971 13507 14977
rect 11977 14943 12035 14949
rect 11977 14909 11989 14943
rect 12023 14909 12035 14943
rect 13464 14940 13492 14971
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 14366 14968 14372 15020
rect 14424 14968 14430 15020
rect 16025 15011 16083 15017
rect 16025 15008 16037 15011
rect 14568 14980 16037 15008
rect 11977 14903 12035 14909
rect 12084 14912 13492 14940
rect 13725 14943 13783 14949
rect 11422 14872 11428 14884
rect 11072 14844 11428 14872
rect 11422 14832 11428 14844
rect 11480 14872 11486 14884
rect 12084 14872 12112 14912
rect 13725 14909 13737 14943
rect 13771 14940 13783 14943
rect 14458 14940 14464 14952
rect 13771 14912 14464 14940
rect 13771 14909 13783 14912
rect 13725 14903 13783 14909
rect 14458 14900 14464 14912
rect 14516 14900 14522 14952
rect 11480 14844 12112 14872
rect 11480 14832 11486 14844
rect 12250 14832 12256 14884
rect 12308 14832 12314 14884
rect 12986 14872 12992 14884
rect 12406 14844 12992 14872
rect 10870 14804 10876 14816
rect 2746 14776 10876 14804
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 10965 14807 11023 14813
rect 10965 14773 10977 14807
rect 11011 14804 11023 14807
rect 12406 14804 12434 14844
rect 12986 14832 12992 14844
rect 13044 14832 13050 14884
rect 11011 14776 12434 14804
rect 12897 14807 12955 14813
rect 11011 14773 11023 14776
rect 10965 14767 11023 14773
rect 12897 14773 12909 14807
rect 12943 14804 12955 14807
rect 13446 14804 13452 14816
rect 12943 14776 13452 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 13722 14764 13728 14816
rect 13780 14804 13786 14816
rect 14568 14804 14596 14980
rect 16025 14977 16037 14980
rect 16071 15008 16083 15011
rect 16071 14980 16804 15008
rect 16071 14977 16083 14980
rect 16025 14971 16083 14977
rect 16776 14940 16804 14980
rect 16850 14968 16856 15020
rect 16908 14968 16914 15020
rect 18064 15008 18092 15116
rect 18966 15104 18972 15156
rect 19024 15144 19030 15156
rect 19077 15147 19135 15153
rect 19077 15144 19089 15147
rect 19024 15116 19089 15144
rect 19024 15104 19030 15116
rect 19077 15113 19089 15116
rect 19123 15113 19135 15147
rect 19077 15107 19135 15113
rect 19242 15104 19248 15156
rect 19300 15104 19306 15156
rect 19889 15147 19947 15153
rect 19889 15113 19901 15147
rect 19935 15144 19947 15147
rect 20438 15144 20444 15156
rect 19935 15116 20444 15144
rect 19935 15113 19947 15116
rect 19889 15107 19947 15113
rect 20438 15104 20444 15116
rect 20496 15104 20502 15156
rect 22554 15144 22560 15156
rect 22066 15116 22560 15144
rect 18138 15036 18144 15088
rect 18196 15036 18202 15088
rect 18690 15036 18696 15088
rect 18748 15076 18754 15088
rect 18874 15076 18880 15088
rect 18748 15048 18880 15076
rect 18748 15036 18754 15048
rect 18874 15036 18880 15048
rect 18932 15036 18938 15088
rect 22066 15076 22094 15116
rect 22554 15104 22560 15116
rect 22612 15144 22618 15156
rect 22738 15144 22744 15156
rect 22612 15116 22744 15144
rect 22612 15104 22618 15116
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 22833 15147 22891 15153
rect 22833 15113 22845 15147
rect 22879 15144 22891 15147
rect 23658 15144 23664 15156
rect 22879 15116 23664 15144
rect 22879 15113 22891 15116
rect 22833 15107 22891 15113
rect 23658 15104 23664 15116
rect 23716 15104 23722 15156
rect 25130 15144 25136 15156
rect 24044 15116 25136 15144
rect 18984 15048 22094 15076
rect 18984 15008 19012 15048
rect 16960 14980 17816 15008
rect 18064 14980 19012 15008
rect 16960 14940 16988 14980
rect 16776 14912 16988 14940
rect 17034 14900 17040 14952
rect 17092 14900 17098 14952
rect 17052 14872 17080 14900
rect 17681 14875 17739 14881
rect 17681 14872 17693 14875
rect 17052 14844 17693 14872
rect 17681 14841 17693 14844
rect 17727 14841 17739 14875
rect 17788 14872 17816 14980
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19705 15011 19763 15017
rect 19705 15008 19717 15011
rect 19484 14980 19717 15008
rect 19484 14968 19490 14980
rect 19705 14977 19717 14980
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 20254 14968 20260 15020
rect 20312 15008 20318 15020
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 20312 14980 22017 15008
rect 20312 14968 20318 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 15008 22155 15011
rect 22646 15008 22652 15020
rect 22143 14980 22652 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 22646 14968 22652 14980
rect 22704 14968 22710 15020
rect 22738 14968 22744 15020
rect 22796 15017 22802 15020
rect 22796 15011 22832 15017
rect 22820 14977 22832 15011
rect 22796 14971 22832 14977
rect 23201 15011 23259 15017
rect 23201 14977 23213 15011
rect 23247 15008 23259 15011
rect 23474 15008 23480 15020
rect 23247 14980 23480 15008
rect 23247 14977 23259 14980
rect 23201 14971 23259 14977
rect 22796 14968 22802 14971
rect 23474 14968 23480 14980
rect 23532 15008 23538 15020
rect 24044 15008 24072 15116
rect 25130 15104 25136 15116
rect 25188 15104 25194 15156
rect 25317 15147 25375 15153
rect 25317 15113 25329 15147
rect 25363 15144 25375 15147
rect 26694 15144 26700 15156
rect 25363 15116 26700 15144
rect 25363 15113 25375 15116
rect 25317 15107 25375 15113
rect 26694 15104 26700 15116
rect 26752 15104 26758 15156
rect 27890 15104 27896 15156
rect 27948 15104 27954 15156
rect 29454 15144 29460 15156
rect 28000 15116 29460 15144
rect 24302 15036 24308 15088
rect 24360 15036 24366 15088
rect 24397 15079 24455 15085
rect 24397 15045 24409 15079
rect 24443 15076 24455 15079
rect 24946 15076 24952 15088
rect 24443 15048 24952 15076
rect 24443 15045 24455 15048
rect 24397 15039 24455 15045
rect 24946 15036 24952 15048
rect 25004 15076 25010 15088
rect 25685 15079 25743 15085
rect 25685 15076 25697 15079
rect 25004 15048 25697 15076
rect 25004 15036 25010 15048
rect 25685 15045 25697 15048
rect 25731 15045 25743 15079
rect 25685 15039 25743 15045
rect 26326 15036 26332 15088
rect 26384 15076 26390 15088
rect 27430 15076 27436 15088
rect 26384 15048 27436 15076
rect 26384 15036 26390 15048
rect 27430 15036 27436 15048
rect 27488 15076 27494 15088
rect 28000 15076 28028 15116
rect 29454 15104 29460 15116
rect 29512 15104 29518 15156
rect 29546 15104 29552 15156
rect 29604 15144 29610 15156
rect 29825 15147 29883 15153
rect 29825 15144 29837 15147
rect 29604 15116 29837 15144
rect 29604 15104 29610 15116
rect 29825 15113 29837 15116
rect 29871 15113 29883 15147
rect 29825 15107 29883 15113
rect 30834 15104 30840 15156
rect 30892 15144 30898 15156
rect 32950 15144 32956 15156
rect 30892 15116 32956 15144
rect 30892 15104 30898 15116
rect 32950 15104 32956 15116
rect 33008 15104 33014 15156
rect 34422 15104 34428 15156
rect 34480 15144 34486 15156
rect 34480 15116 36676 15144
rect 34480 15104 34486 15116
rect 28718 15085 28724 15088
rect 28712 15076 28724 15085
rect 27488 15048 28028 15076
rect 28679 15048 28724 15076
rect 27488 15036 27494 15048
rect 28712 15039 28724 15048
rect 28718 15036 28724 15039
rect 28776 15036 28782 15088
rect 29086 15076 29092 15088
rect 28920 15048 29092 15076
rect 23532 14980 24072 15008
rect 23532 14968 23538 14980
rect 24118 14968 24124 15020
rect 24176 14968 24182 15020
rect 24210 14968 24216 15020
rect 24268 15008 24274 15020
rect 24494 15011 24552 15017
rect 24494 15008 24506 15011
rect 24268 14980 24506 15008
rect 24268 14968 24274 14980
rect 24494 14977 24506 14980
rect 24540 14977 24552 15011
rect 24494 14971 24552 14977
rect 25130 14968 25136 15020
rect 25188 15008 25194 15020
rect 25498 15008 25504 15020
rect 25188 14980 25504 15008
rect 25188 14968 25194 14980
rect 25498 14968 25504 14980
rect 25556 15008 25562 15020
rect 25556 14980 25728 15008
rect 25556 14968 25562 14980
rect 18233 14943 18291 14949
rect 18233 14909 18245 14943
rect 18279 14940 18291 14943
rect 19978 14940 19984 14952
rect 18279 14912 19984 14940
rect 18279 14909 18291 14912
rect 18233 14903 18291 14909
rect 19978 14900 19984 14912
rect 20036 14900 20042 14952
rect 22670 14940 22698 14968
rect 23293 14943 23351 14949
rect 23293 14940 23305 14943
rect 22670 14912 23305 14940
rect 23293 14909 23305 14912
rect 23339 14909 23351 14943
rect 25700 14940 25728 14980
rect 25774 14968 25780 15020
rect 25832 14968 25838 15020
rect 27706 14968 27712 15020
rect 27764 14968 27770 15020
rect 28920 15008 28948 15048
rect 29086 15036 29092 15048
rect 29144 15076 29150 15088
rect 30190 15076 30196 15088
rect 29144 15048 30196 15076
rect 29144 15036 29150 15048
rect 30190 15036 30196 15048
rect 30248 15036 30254 15088
rect 30926 15036 30932 15088
rect 30984 15076 30990 15088
rect 31478 15076 31484 15088
rect 30984 15048 31484 15076
rect 30984 15036 30990 15048
rect 31478 15036 31484 15048
rect 31536 15036 31542 15088
rect 36538 15076 36544 15088
rect 34440 15048 36544 15076
rect 28368 14980 28948 15008
rect 25869 14943 25927 14949
rect 25869 14940 25881 14943
rect 25700 14912 25881 14940
rect 23293 14903 23351 14909
rect 25869 14909 25881 14912
rect 25915 14940 25927 14943
rect 27430 14940 27436 14952
rect 25915 14912 27436 14940
rect 25915 14909 25927 14912
rect 25869 14903 25927 14909
rect 27430 14900 27436 14912
rect 27488 14900 27494 14952
rect 27525 14943 27583 14949
rect 27525 14909 27537 14943
rect 27571 14940 27583 14943
rect 28368 14940 28396 14980
rect 28994 14968 29000 15020
rect 29052 15008 29058 15020
rect 30377 15011 30435 15017
rect 30377 15008 30389 15011
rect 29052 14980 30389 15008
rect 29052 14968 29058 14980
rect 30377 14977 30389 14980
rect 30423 14977 30435 15011
rect 30377 14971 30435 14977
rect 30558 14968 30564 15020
rect 30616 15008 30622 15020
rect 32122 15008 32128 15020
rect 30616 14980 32128 15008
rect 30616 14968 30622 14980
rect 32122 14968 32128 14980
rect 32180 14968 32186 15020
rect 32306 14968 32312 15020
rect 32364 15008 32370 15020
rect 32858 15008 32864 15020
rect 32364 14980 32864 15008
rect 32364 14968 32370 14980
rect 32858 14968 32864 14980
rect 32916 14968 32922 15020
rect 34440 15017 34468 15048
rect 36538 15036 36544 15048
rect 36596 15036 36602 15088
rect 36648 15076 36676 15116
rect 37918 15104 37924 15156
rect 37976 15144 37982 15156
rect 38657 15147 38715 15153
rect 38657 15144 38669 15147
rect 37976 15116 38669 15144
rect 37976 15104 37982 15116
rect 38657 15113 38669 15116
rect 38703 15113 38715 15147
rect 38657 15107 38715 15113
rect 39298 15104 39304 15156
rect 39356 15144 39362 15156
rect 41506 15144 41512 15156
rect 39356 15116 41512 15144
rect 39356 15104 39362 15116
rect 40862 15076 40868 15088
rect 36648 15048 40868 15076
rect 40862 15036 40868 15048
rect 40920 15036 40926 15088
rect 41432 15085 41460 15116
rect 41506 15104 41512 15116
rect 41564 15104 41570 15156
rect 41785 15147 41843 15153
rect 41785 15113 41797 15147
rect 41831 15144 41843 15147
rect 41966 15144 41972 15156
rect 41831 15116 41972 15144
rect 41831 15113 41843 15116
rect 41785 15107 41843 15113
rect 41966 15104 41972 15116
rect 42024 15104 42030 15156
rect 42242 15104 42248 15156
rect 42300 15144 42306 15156
rect 43073 15147 43131 15153
rect 43073 15144 43085 15147
rect 42300 15116 43085 15144
rect 42300 15104 42306 15116
rect 43073 15113 43085 15116
rect 43119 15113 43131 15147
rect 43073 15107 43131 15113
rect 47765 15147 47823 15153
rect 47765 15113 47777 15147
rect 47811 15144 47823 15147
rect 47854 15144 47860 15156
rect 47811 15116 47860 15144
rect 47811 15113 47823 15116
rect 47765 15107 47823 15113
rect 47854 15104 47860 15116
rect 47912 15104 47918 15156
rect 41417 15079 41475 15085
rect 41417 15045 41429 15079
rect 41463 15045 41475 15079
rect 41417 15039 41475 15045
rect 42702 15036 42708 15088
rect 42760 15076 42766 15088
rect 48406 15076 48412 15088
rect 42760 15048 48412 15076
rect 42760 15036 42766 15048
rect 48406 15036 48412 15048
rect 48464 15036 48470 15088
rect 34698 15017 34704 15020
rect 34425 15011 34483 15017
rect 34425 14977 34437 15011
rect 34471 14977 34483 15011
rect 34692 15008 34704 15017
rect 34659 14980 34704 15008
rect 34425 14971 34483 14977
rect 34692 14971 34704 14980
rect 34698 14968 34704 14971
rect 34756 14968 34762 15020
rect 38654 15011 38712 15017
rect 38654 14977 38666 15011
rect 38700 15008 38712 15011
rect 40034 15008 40040 15020
rect 38700 14980 40040 15008
rect 38700 14977 38712 14980
rect 38654 14971 38712 14977
rect 40034 14968 40040 14980
rect 40092 14968 40098 15020
rect 41233 15011 41291 15017
rect 41233 14977 41245 15011
rect 41279 14977 41291 15011
rect 41233 14971 41291 14977
rect 27571 14912 28396 14940
rect 28445 14943 28503 14949
rect 27571 14909 27583 14912
rect 27525 14903 27583 14909
rect 28445 14909 28457 14943
rect 28491 14909 28503 14943
rect 28445 14903 28503 14909
rect 21818 14872 21824 14884
rect 17788 14844 21824 14872
rect 17681 14835 17739 14841
rect 21818 14832 21824 14844
rect 21876 14832 21882 14884
rect 22664 14844 24624 14872
rect 13780 14776 14596 14804
rect 13780 14764 13786 14776
rect 15010 14764 15016 14816
rect 15068 14764 15074 14816
rect 16206 14764 16212 14816
rect 16264 14764 16270 14816
rect 16850 14764 16856 14816
rect 16908 14804 16914 14816
rect 17037 14807 17095 14813
rect 17037 14804 17049 14807
rect 16908 14776 17049 14804
rect 16908 14764 16914 14776
rect 17037 14773 17049 14776
rect 17083 14773 17095 14807
rect 17037 14767 17095 14773
rect 19061 14807 19119 14813
rect 19061 14773 19073 14807
rect 19107 14804 19119 14807
rect 19150 14804 19156 14816
rect 19107 14776 19156 14804
rect 19107 14773 19119 14776
rect 19061 14767 19119 14773
rect 19150 14764 19156 14776
rect 19208 14764 19214 14816
rect 22664 14813 22692 14844
rect 22649 14807 22707 14813
rect 22649 14773 22661 14807
rect 22695 14773 22707 14807
rect 22649 14767 22707 14773
rect 23290 14764 23296 14816
rect 23348 14804 23354 14816
rect 24302 14804 24308 14816
rect 23348 14776 24308 14804
rect 23348 14764 23354 14776
rect 24302 14764 24308 14776
rect 24360 14764 24366 14816
rect 24596 14804 24624 14844
rect 24670 14832 24676 14884
rect 24728 14832 24734 14884
rect 25498 14832 25504 14884
rect 25556 14872 25562 14884
rect 25774 14872 25780 14884
rect 25556 14844 25780 14872
rect 25556 14832 25562 14844
rect 25774 14832 25780 14844
rect 25832 14832 25838 14884
rect 26050 14804 26056 14816
rect 24596 14776 26056 14804
rect 26050 14764 26056 14776
rect 26108 14764 26114 14816
rect 28460 14804 28488 14903
rect 31754 14900 31760 14952
rect 31812 14940 31818 14952
rect 32585 14943 32643 14949
rect 32585 14940 32597 14943
rect 31812 14912 32597 14940
rect 31812 14900 31818 14912
rect 32585 14909 32597 14912
rect 32631 14909 32643 14943
rect 32585 14903 32643 14909
rect 38746 14900 38752 14952
rect 38804 14940 38810 14952
rect 39117 14943 39175 14949
rect 39117 14940 39129 14943
rect 38804 14912 39129 14940
rect 38804 14900 38810 14912
rect 39117 14909 39129 14912
rect 39163 14909 39175 14943
rect 41248 14940 41276 14971
rect 41506 14968 41512 15020
rect 41564 14968 41570 15020
rect 41598 14968 41604 15020
rect 41656 14968 41662 15020
rect 42794 14968 42800 15020
rect 42852 15008 42858 15020
rect 42981 15011 43039 15017
rect 42981 15008 42993 15011
rect 42852 14980 42993 15008
rect 42852 14968 42858 14980
rect 42981 14977 42993 14980
rect 43027 14977 43039 15011
rect 42981 14971 43039 14977
rect 48133 15011 48191 15017
rect 48133 14977 48145 15011
rect 48179 15008 48191 15011
rect 58434 15008 58440 15020
rect 48179 14980 58440 15008
rect 48179 14977 48191 14980
rect 48133 14971 48191 14977
rect 58434 14968 58440 14980
rect 58492 14968 58498 15020
rect 41248 14912 46336 14940
rect 39117 14903 39175 14909
rect 29454 14832 29460 14884
rect 29512 14872 29518 14884
rect 46198 14872 46204 14884
rect 29512 14844 31754 14872
rect 29512 14832 29518 14844
rect 29730 14804 29736 14816
rect 28460 14776 29736 14804
rect 29730 14764 29736 14776
rect 29788 14764 29794 14816
rect 31726 14804 31754 14844
rect 35544 14844 46204 14872
rect 31938 14804 31944 14816
rect 31726 14776 31944 14804
rect 31938 14764 31944 14776
rect 31996 14764 32002 14816
rect 32674 14764 32680 14816
rect 32732 14804 32738 14816
rect 33873 14807 33931 14813
rect 33873 14804 33885 14807
rect 32732 14776 33885 14804
rect 32732 14764 32738 14776
rect 33873 14773 33885 14776
rect 33919 14804 33931 14807
rect 35544 14804 35572 14844
rect 46198 14832 46204 14844
rect 46256 14832 46262 14884
rect 33919 14776 35572 14804
rect 33919 14773 33931 14776
rect 33873 14767 33931 14773
rect 35618 14764 35624 14816
rect 35676 14804 35682 14816
rect 35805 14807 35863 14813
rect 35805 14804 35817 14807
rect 35676 14776 35817 14804
rect 35676 14764 35682 14776
rect 35805 14773 35817 14776
rect 35851 14773 35863 14807
rect 35805 14767 35863 14773
rect 38473 14807 38531 14813
rect 38473 14773 38485 14807
rect 38519 14804 38531 14807
rect 38930 14804 38936 14816
rect 38519 14776 38936 14804
rect 38519 14773 38531 14776
rect 38473 14767 38531 14773
rect 38930 14764 38936 14776
rect 38988 14764 38994 14816
rect 39025 14807 39083 14813
rect 39025 14773 39037 14807
rect 39071 14804 39083 14807
rect 39114 14804 39120 14816
rect 39071 14776 39120 14804
rect 39071 14773 39083 14776
rect 39025 14767 39083 14773
rect 39114 14764 39120 14776
rect 39172 14764 39178 14816
rect 40862 14764 40868 14816
rect 40920 14804 40926 14816
rect 42702 14804 42708 14816
rect 40920 14776 42708 14804
rect 40920 14764 40926 14776
rect 42702 14764 42708 14776
rect 42760 14764 42766 14816
rect 42978 14764 42984 14816
rect 43036 14804 43042 14816
rect 44266 14804 44272 14816
rect 43036 14776 44272 14804
rect 43036 14764 43042 14776
rect 44266 14764 44272 14776
rect 44324 14764 44330 14816
rect 46308 14804 46336 14912
rect 48222 14900 48228 14952
rect 48280 14900 48286 14952
rect 48317 14943 48375 14949
rect 48317 14909 48329 14943
rect 48363 14909 48375 14943
rect 48317 14903 48375 14909
rect 46842 14832 46848 14884
rect 46900 14872 46906 14884
rect 48332 14872 48360 14903
rect 46900 14844 48360 14872
rect 46900 14832 46906 14844
rect 50154 14804 50160 14816
rect 46308 14776 50160 14804
rect 50154 14764 50160 14776
rect 50212 14764 50218 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 12805 14603 12863 14609
rect 12805 14569 12817 14603
rect 12851 14600 12863 14603
rect 17034 14600 17040 14612
rect 12851 14572 16712 14600
rect 12851 14569 12863 14572
rect 12805 14563 12863 14569
rect 9306 14424 9312 14476
rect 9364 14424 9370 14476
rect 11422 14424 11428 14476
rect 11480 14424 11486 14476
rect 13998 14464 14004 14476
rect 13464 14436 14004 14464
rect 1578 14356 1584 14408
rect 1636 14356 1642 14408
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 8846 14396 8852 14408
rect 8343 14368 8852 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 9585 14399 9643 14405
rect 9585 14365 9597 14399
rect 9631 14396 9643 14399
rect 9858 14396 9864 14408
rect 9631 14368 9864 14396
rect 9631 14365 9643 14368
rect 9585 14359 9643 14365
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 13464 14405 13492 14436
rect 13998 14424 14004 14436
rect 14056 14424 14062 14476
rect 14182 14424 14188 14476
rect 14240 14464 14246 14476
rect 14369 14467 14427 14473
rect 14369 14464 14381 14467
rect 14240 14436 14381 14464
rect 14240 14424 14246 14436
rect 14369 14433 14381 14436
rect 14415 14464 14427 14467
rect 14415 14436 16620 14464
rect 14415 14433 14427 14436
rect 14369 14427 14427 14433
rect 13449 14399 13507 14405
rect 13449 14365 13461 14399
rect 13495 14365 13507 14399
rect 14645 14399 14703 14405
rect 14645 14396 14657 14399
rect 13449 14359 13507 14365
rect 13648 14368 14657 14396
rect 934 14288 940 14340
rect 992 14328 998 14340
rect 1857 14331 1915 14337
rect 1857 14328 1869 14331
rect 992 14300 1869 14328
rect 992 14288 998 14300
rect 1857 14297 1869 14300
rect 1903 14297 1915 14331
rect 1857 14291 1915 14297
rect 11692 14331 11750 14337
rect 11692 14297 11704 14331
rect 11738 14328 11750 14331
rect 11882 14328 11888 14340
rect 11738 14300 11888 14328
rect 11738 14297 11750 14300
rect 11692 14291 11750 14297
rect 11882 14288 11888 14300
rect 11940 14288 11946 14340
rect 8481 14263 8539 14269
rect 8481 14229 8493 14263
rect 8527 14260 8539 14263
rect 9674 14260 9680 14272
rect 8527 14232 9680 14260
rect 8527 14229 8539 14232
rect 8481 14223 8539 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 10226 14220 10232 14272
rect 10284 14260 10290 14272
rect 13648 14269 13676 14368
rect 14645 14365 14657 14368
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 10689 14263 10747 14269
rect 10689 14260 10701 14263
rect 10284 14232 10701 14260
rect 10284 14220 10290 14232
rect 10689 14229 10701 14232
rect 10735 14229 10747 14263
rect 10689 14223 10747 14229
rect 13633 14263 13691 14269
rect 13633 14229 13645 14263
rect 13679 14229 13691 14263
rect 13633 14223 13691 14229
rect 15562 14220 15568 14272
rect 15620 14260 15626 14272
rect 15749 14263 15807 14269
rect 15749 14260 15761 14263
rect 15620 14232 15761 14260
rect 15620 14220 15626 14232
rect 15749 14229 15761 14232
rect 15795 14229 15807 14263
rect 16592 14260 16620 14436
rect 16684 14328 16712 14572
rect 16776 14572 17040 14600
rect 16776 14476 16804 14572
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 18690 14560 18696 14612
rect 18748 14600 18754 14612
rect 19150 14600 19156 14612
rect 18748 14572 19156 14600
rect 18748 14560 18754 14572
rect 19150 14560 19156 14572
rect 19208 14600 19214 14612
rect 19797 14603 19855 14609
rect 19797 14600 19809 14603
rect 19208 14572 19809 14600
rect 19208 14560 19214 14572
rect 19797 14569 19809 14572
rect 19843 14569 19855 14603
rect 19797 14563 19855 14569
rect 21818 14560 21824 14612
rect 21876 14560 21882 14612
rect 26605 14603 26663 14609
rect 26605 14600 26617 14603
rect 22066 14572 26617 14600
rect 17954 14492 17960 14544
rect 18012 14532 18018 14544
rect 22066 14532 22094 14572
rect 26605 14569 26617 14572
rect 26651 14569 26663 14603
rect 26605 14563 26663 14569
rect 26694 14560 26700 14612
rect 26752 14600 26758 14612
rect 31662 14600 31668 14612
rect 26752 14572 31668 14600
rect 26752 14560 26758 14572
rect 31662 14560 31668 14572
rect 31720 14560 31726 14612
rect 31754 14560 31760 14612
rect 31812 14560 31818 14612
rect 32122 14560 32128 14612
rect 32180 14600 32186 14612
rect 33594 14600 33600 14612
rect 32180 14572 33600 14600
rect 32180 14560 32186 14572
rect 33594 14560 33600 14572
rect 33652 14560 33658 14612
rect 38010 14560 38016 14612
rect 38068 14600 38074 14612
rect 39393 14603 39451 14609
rect 39393 14600 39405 14603
rect 38068 14572 39405 14600
rect 38068 14560 38074 14572
rect 39393 14569 39405 14572
rect 39439 14600 39451 14603
rect 52362 14600 52368 14612
rect 39439 14572 52368 14600
rect 39439 14569 39451 14572
rect 39393 14563 39451 14569
rect 52362 14560 52368 14572
rect 52420 14560 52426 14612
rect 58066 14560 58072 14612
rect 58124 14560 58130 14612
rect 18012 14504 19656 14532
rect 18012 14492 18018 14504
rect 16758 14424 16764 14476
rect 16816 14424 16822 14476
rect 17770 14424 17776 14476
rect 17828 14464 17834 14476
rect 18785 14467 18843 14473
rect 18785 14464 18797 14467
rect 17828 14436 18797 14464
rect 17828 14424 17834 14436
rect 18785 14433 18797 14436
rect 18831 14433 18843 14467
rect 18785 14427 18843 14433
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 17017 14399 17075 14405
rect 17017 14396 17029 14399
rect 16908 14368 17029 14396
rect 16908 14356 16914 14368
rect 17017 14365 17029 14368
rect 17063 14365 17075 14399
rect 17017 14359 17075 14365
rect 18690 14356 18696 14408
rect 18748 14356 18754 14408
rect 18874 14356 18880 14408
rect 18932 14356 18938 14408
rect 19334 14356 19340 14408
rect 19392 14396 19398 14408
rect 19628 14405 19656 14504
rect 21652 14504 22094 14532
rect 22833 14535 22891 14541
rect 19429 14399 19487 14405
rect 19429 14396 19441 14399
rect 19392 14368 19441 14396
rect 19392 14356 19398 14368
rect 19429 14365 19441 14368
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 20254 14356 20260 14408
rect 20312 14356 20318 14408
rect 21652 14405 21680 14504
rect 22833 14501 22845 14535
rect 22879 14532 22891 14535
rect 25314 14532 25320 14544
rect 22879 14504 25320 14532
rect 22879 14501 22891 14504
rect 22833 14495 22891 14501
rect 25314 14492 25320 14504
rect 25372 14492 25378 14544
rect 25958 14492 25964 14544
rect 26016 14532 26022 14544
rect 32493 14535 32551 14541
rect 26016 14504 29684 14532
rect 26016 14492 26022 14504
rect 23293 14467 23351 14473
rect 23293 14433 23305 14467
rect 23339 14464 23351 14467
rect 23474 14464 23480 14476
rect 23339 14436 23480 14464
rect 23339 14433 23351 14436
rect 23293 14427 23351 14433
rect 23474 14424 23480 14436
rect 23532 14424 23538 14476
rect 23658 14424 23664 14476
rect 23716 14464 23722 14476
rect 23937 14467 23995 14473
rect 23937 14464 23949 14467
rect 23716 14436 23949 14464
rect 23716 14424 23722 14436
rect 23937 14433 23949 14436
rect 23983 14433 23995 14467
rect 23937 14427 23995 14433
rect 28813 14467 28871 14473
rect 28813 14433 28825 14467
rect 28859 14464 28871 14467
rect 29086 14464 29092 14476
rect 28859 14436 29092 14464
rect 28859 14433 28871 14436
rect 28813 14427 28871 14433
rect 29086 14424 29092 14436
rect 29144 14424 29150 14476
rect 21637 14399 21695 14405
rect 21637 14365 21649 14399
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 22922 14396 22928 14408
rect 22152 14368 22928 14396
rect 22152 14356 22158 14368
rect 22922 14356 22928 14368
rect 22980 14396 22986 14408
rect 23017 14399 23075 14405
rect 23017 14396 23029 14399
rect 22980 14368 23029 14396
rect 22980 14356 22986 14368
rect 23017 14365 23029 14368
rect 23063 14365 23075 14399
rect 23017 14359 23075 14365
rect 23106 14356 23112 14408
rect 23164 14356 23170 14408
rect 23382 14356 23388 14408
rect 23440 14356 23446 14408
rect 23845 14399 23903 14405
rect 23845 14365 23857 14399
rect 23891 14365 23903 14399
rect 23845 14359 23903 14365
rect 24029 14399 24087 14405
rect 24029 14365 24041 14399
rect 24075 14396 24087 14399
rect 24210 14396 24216 14408
rect 24075 14368 24216 14396
rect 24075 14365 24087 14368
rect 24029 14359 24087 14365
rect 22554 14328 22560 14340
rect 16684 14300 22560 14328
rect 22554 14288 22560 14300
rect 22612 14288 22618 14340
rect 22646 14288 22652 14340
rect 22704 14328 22710 14340
rect 23198 14328 23204 14340
rect 22704 14300 23204 14328
rect 22704 14288 22710 14300
rect 23198 14288 23204 14300
rect 23256 14328 23262 14340
rect 23860 14328 23888 14359
rect 24210 14356 24216 14368
rect 24268 14356 24274 14408
rect 24946 14356 24952 14408
rect 25004 14356 25010 14408
rect 25317 14399 25375 14405
rect 25317 14365 25329 14399
rect 25363 14396 25375 14399
rect 25498 14398 25504 14408
rect 25424 14396 25504 14398
rect 25363 14370 25504 14396
rect 25363 14368 25452 14370
rect 25363 14365 25375 14368
rect 25317 14359 25375 14365
rect 25498 14356 25504 14370
rect 25556 14396 25562 14408
rect 25682 14396 25688 14408
rect 25556 14368 25688 14396
rect 25556 14356 25562 14368
rect 25682 14356 25688 14368
rect 25740 14356 25746 14408
rect 25958 14356 25964 14408
rect 26016 14396 26022 14408
rect 26421 14399 26479 14405
rect 26421 14396 26433 14399
rect 26016 14368 26433 14396
rect 26016 14356 26022 14368
rect 26421 14365 26433 14368
rect 26467 14365 26479 14399
rect 26421 14359 26479 14365
rect 28997 14399 29055 14405
rect 28997 14365 29009 14399
rect 29043 14396 29055 14399
rect 29362 14396 29368 14408
rect 29043 14368 29368 14396
rect 29043 14365 29055 14368
rect 28997 14359 29055 14365
rect 29362 14356 29368 14368
rect 29420 14356 29426 14408
rect 29656 14396 29684 14504
rect 32493 14501 32505 14535
rect 32539 14501 32551 14535
rect 32493 14495 32551 14501
rect 29730 14424 29736 14476
rect 29788 14424 29794 14476
rect 32508 14464 32536 14495
rect 32950 14492 32956 14544
rect 33008 14532 33014 14544
rect 37918 14532 37924 14544
rect 33008 14504 37924 14532
rect 33008 14492 33014 14504
rect 37918 14492 37924 14504
rect 37976 14492 37982 14544
rect 42978 14464 42984 14476
rect 31772 14436 32536 14464
rect 32600 14436 37596 14464
rect 31772 14405 31800 14436
rect 31757 14399 31815 14405
rect 29656 14368 31248 14396
rect 23256 14300 23888 14328
rect 23256 14288 23262 14300
rect 24670 14288 24676 14340
rect 24728 14328 24734 14340
rect 25133 14331 25191 14337
rect 25133 14328 25145 14331
rect 24728 14300 25145 14328
rect 24728 14288 24734 14300
rect 25133 14297 25145 14300
rect 25179 14297 25191 14331
rect 25133 14291 25191 14297
rect 25225 14331 25283 14337
rect 25225 14297 25237 14331
rect 25271 14297 25283 14331
rect 25225 14291 25283 14297
rect 29181 14331 29239 14337
rect 29181 14297 29193 14331
rect 29227 14328 29239 14331
rect 29978 14331 30036 14337
rect 29978 14328 29990 14331
rect 29227 14300 29990 14328
rect 29227 14297 29239 14300
rect 29181 14291 29239 14297
rect 29978 14297 29990 14300
rect 30024 14297 30036 14331
rect 29978 14291 30036 14297
rect 16758 14260 16764 14272
rect 16592 14232 16764 14260
rect 15749 14223 15807 14229
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 18141 14263 18199 14269
rect 18141 14229 18153 14263
rect 18187 14260 18199 14263
rect 20162 14260 20168 14272
rect 18187 14232 20168 14260
rect 18187 14229 18199 14232
rect 18141 14223 18199 14229
rect 20162 14220 20168 14232
rect 20220 14220 20226 14272
rect 20441 14263 20499 14269
rect 20441 14229 20453 14263
rect 20487 14260 20499 14263
rect 20622 14260 20628 14272
rect 20487 14232 20628 14260
rect 20487 14229 20499 14232
rect 20441 14223 20499 14229
rect 20622 14220 20628 14232
rect 20680 14220 20686 14272
rect 25240 14260 25268 14291
rect 25314 14260 25320 14272
rect 25240 14232 25320 14260
rect 25314 14220 25320 14232
rect 25372 14220 25378 14272
rect 25498 14220 25504 14272
rect 25556 14220 25562 14272
rect 27430 14220 27436 14272
rect 27488 14260 27494 14272
rect 29454 14260 29460 14272
rect 27488 14232 29460 14260
rect 27488 14220 27494 14232
rect 29454 14220 29460 14232
rect 29512 14220 29518 14272
rect 31018 14220 31024 14272
rect 31076 14260 31082 14272
rect 31113 14263 31171 14269
rect 31113 14260 31125 14263
rect 31076 14232 31125 14260
rect 31076 14220 31082 14232
rect 31113 14229 31125 14232
rect 31159 14229 31171 14263
rect 31220 14260 31248 14368
rect 31757 14365 31769 14399
rect 31803 14365 31815 14399
rect 31757 14359 31815 14365
rect 31941 14399 31999 14405
rect 31941 14365 31953 14399
rect 31987 14396 31999 14399
rect 32600 14396 32628 14436
rect 37568 14408 37596 14436
rect 41386 14436 42984 14464
rect 31987 14368 32628 14396
rect 31987 14365 31999 14368
rect 31941 14359 31999 14365
rect 31294 14288 31300 14340
rect 31352 14328 31358 14340
rect 31956 14328 31984 14359
rect 32674 14356 32680 14408
rect 32732 14356 32738 14408
rect 32950 14356 32956 14408
rect 33008 14356 33014 14408
rect 33137 14399 33195 14405
rect 33137 14365 33149 14399
rect 33183 14365 33195 14399
rect 33137 14359 33195 14365
rect 31352 14300 31984 14328
rect 31352 14288 31358 14300
rect 32582 14288 32588 14340
rect 32640 14328 32646 14340
rect 32858 14328 32864 14340
rect 32640 14300 32864 14328
rect 32640 14288 32646 14300
rect 32858 14288 32864 14300
rect 32916 14328 32922 14340
rect 33152 14328 33180 14359
rect 33594 14356 33600 14408
rect 33652 14356 33658 14408
rect 37366 14356 37372 14408
rect 37424 14356 37430 14408
rect 37550 14356 37556 14408
rect 37608 14356 37614 14408
rect 38013 14399 38071 14405
rect 38013 14365 38025 14399
rect 38059 14396 38071 14399
rect 40037 14399 40095 14405
rect 40037 14396 40049 14399
rect 38059 14368 40049 14396
rect 38059 14365 38071 14368
rect 38013 14359 38071 14365
rect 40037 14365 40049 14368
rect 40083 14396 40095 14399
rect 40678 14396 40684 14408
rect 40083 14368 40684 14396
rect 40083 14365 40095 14368
rect 40037 14359 40095 14365
rect 40678 14356 40684 14368
rect 40736 14396 40742 14408
rect 41386 14396 41414 14436
rect 42978 14424 42984 14436
rect 43036 14424 43042 14476
rect 43254 14424 43260 14476
rect 43312 14424 43318 14476
rect 40736 14368 41414 14396
rect 40736 14356 40742 14368
rect 41966 14356 41972 14408
rect 42024 14396 42030 14408
rect 42061 14399 42119 14405
rect 42061 14396 42073 14399
rect 42024 14368 42073 14396
rect 42024 14356 42030 14368
rect 42061 14365 42073 14368
rect 42107 14396 42119 14399
rect 42242 14396 42248 14408
rect 42107 14368 42248 14396
rect 42107 14365 42119 14368
rect 42061 14359 42119 14365
rect 42242 14356 42248 14368
rect 42300 14356 42306 14408
rect 42334 14356 42340 14408
rect 42392 14396 42398 14408
rect 42702 14396 42708 14408
rect 42392 14368 42708 14396
rect 42392 14356 42398 14368
rect 42702 14356 42708 14368
rect 42760 14356 42766 14408
rect 49050 14396 49056 14408
rect 43088 14368 49056 14396
rect 32916 14300 33180 14328
rect 34333 14331 34391 14337
rect 32916 14288 32922 14300
rect 34333 14297 34345 14331
rect 34379 14328 34391 14331
rect 36078 14328 36084 14340
rect 34379 14300 36084 14328
rect 34379 14297 34391 14300
rect 34333 14291 34391 14297
rect 36078 14288 36084 14300
rect 36136 14288 36142 14340
rect 37461 14331 37519 14337
rect 37461 14297 37473 14331
rect 37507 14328 37519 14331
rect 38258 14331 38316 14337
rect 38258 14328 38270 14331
rect 37507 14300 38270 14328
rect 37507 14297 37519 14300
rect 37461 14291 37519 14297
rect 38258 14297 38270 14300
rect 38304 14297 38316 14331
rect 38258 14291 38316 14297
rect 39022 14288 39028 14340
rect 39080 14328 39086 14340
rect 40282 14331 40340 14337
rect 40282 14328 40294 14331
rect 39080 14300 40294 14328
rect 39080 14288 39086 14300
rect 40282 14297 40294 14300
rect 40328 14297 40340 14331
rect 43088 14328 43116 14368
rect 49050 14356 49056 14368
rect 49108 14356 49114 14408
rect 57974 14356 57980 14408
rect 58032 14356 58038 14408
rect 40282 14291 40340 14297
rect 41432 14300 43116 14328
rect 39114 14260 39120 14272
rect 31220 14232 39120 14260
rect 31113 14223 31171 14229
rect 39114 14220 39120 14232
rect 39172 14220 39178 14272
rect 40034 14220 40040 14272
rect 40092 14260 40098 14272
rect 41432 14269 41460 14300
rect 41417 14263 41475 14269
rect 41417 14260 41429 14263
rect 40092 14232 41429 14260
rect 40092 14220 40098 14232
rect 41417 14229 41429 14232
rect 41463 14229 41475 14263
rect 41417 14223 41475 14229
rect 41506 14220 41512 14272
rect 41564 14260 41570 14272
rect 43990 14260 43996 14272
rect 41564 14232 43996 14260
rect 41564 14220 41570 14232
rect 43990 14220 43996 14232
rect 44048 14220 44054 14272
rect 44542 14220 44548 14272
rect 44600 14260 44606 14272
rect 56870 14260 56876 14272
rect 44600 14232 56876 14260
rect 44600 14220 44606 14232
rect 56870 14220 56876 14232
rect 56928 14220 56934 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 8846 14016 8852 14068
rect 8904 14016 8910 14068
rect 9953 14059 10011 14065
rect 9953 14025 9965 14059
rect 9999 14025 10011 14059
rect 9953 14019 10011 14025
rect 11701 14059 11759 14065
rect 11701 14025 11713 14059
rect 11747 14056 11759 14059
rect 12434 14056 12440 14068
rect 11747 14028 12440 14056
rect 11747 14025 11759 14028
rect 11701 14019 11759 14025
rect 9968 13988 9996 14019
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 12710 14016 12716 14068
rect 12768 14056 12774 14068
rect 13725 14059 13783 14065
rect 13725 14056 13737 14059
rect 12768 14028 13737 14056
rect 12768 14016 12774 14028
rect 13725 14025 13737 14028
rect 13771 14025 13783 14059
rect 16206 14056 16212 14068
rect 13725 14019 13783 14025
rect 14292 14028 16212 14056
rect 11790 13988 11796 14000
rect 8680 13960 9996 13988
rect 11440 13960 11796 13988
rect 8680 13929 8708 13960
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13920 1639 13923
rect 8665 13923 8723 13929
rect 1627 13892 2452 13920
rect 1627 13889 1639 13892
rect 1581 13883 1639 13889
rect 934 13812 940 13864
rect 992 13852 998 13864
rect 2424 13861 2452 13892
rect 8665 13889 8677 13923
rect 8711 13889 8723 13923
rect 8665 13883 8723 13889
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13920 9643 13923
rect 11440 13920 11468 13960
rect 11790 13948 11796 13960
rect 11848 13948 11854 14000
rect 11974 13948 11980 14000
rect 12032 13948 12038 14000
rect 14292 13988 14320 14028
rect 16206 14016 16212 14028
rect 16264 14016 16270 14068
rect 16850 14016 16856 14068
rect 16908 14056 16914 14068
rect 17586 14056 17592 14068
rect 16908 14028 17592 14056
rect 16908 14016 16914 14028
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 18138 14016 18144 14068
rect 18196 14056 18202 14068
rect 18767 14059 18825 14065
rect 18767 14056 18779 14059
rect 18196 14028 18779 14056
rect 18196 14016 18202 14028
rect 18767 14025 18779 14028
rect 18813 14025 18825 14059
rect 20806 14056 20812 14068
rect 18767 14019 18825 14025
rect 19076 14028 20812 14056
rect 19076 13997 19104 14028
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 22005 14059 22063 14065
rect 22005 14056 22017 14059
rect 21468 14028 22017 14056
rect 19061 13991 19119 13997
rect 12406 13960 14320 13988
rect 15120 13960 17540 13988
rect 9631 13892 11468 13920
rect 11992 13920 12020 13948
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11992 13892 12081 13920
rect 9631 13889 9643 13892
rect 9585 13883 9643 13889
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13920 12219 13923
rect 12406 13920 12434 13960
rect 12207 13892 12434 13920
rect 12207 13889 12219 13892
rect 12161 13883 12219 13889
rect 13354 13880 13360 13932
rect 13412 13880 13418 13932
rect 14182 13880 14188 13932
rect 14240 13880 14246 13932
rect 14550 13920 14556 13932
rect 14384 13892 14556 13920
rect 1765 13855 1823 13861
rect 1765 13852 1777 13855
rect 992 13824 1777 13852
rect 992 13812 998 13824
rect 1765 13821 1777 13824
rect 1811 13821 1823 13855
rect 1765 13815 1823 13821
rect 2409 13855 2467 13861
rect 2409 13821 2421 13855
rect 2455 13852 2467 13855
rect 2498 13852 2504 13864
rect 2455 13824 2504 13852
rect 2455 13821 2467 13824
rect 2409 13815 2467 13821
rect 2498 13812 2504 13824
rect 2556 13812 2562 13864
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13852 9551 13855
rect 9766 13852 9772 13864
rect 9539 13824 9772 13852
rect 9539 13821 9551 13824
rect 9493 13815 9551 13821
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 11885 13855 11943 13861
rect 10735 13824 11836 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 10042 13784 10048 13796
rect 3476 13756 10048 13784
rect 3476 13744 3482 13756
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 10965 13787 11023 13793
rect 10965 13753 10977 13787
rect 11011 13784 11023 13787
rect 11606 13784 11612 13796
rect 11011 13756 11612 13784
rect 11011 13753 11023 13756
rect 10965 13747 11023 13753
rect 11606 13744 11612 13756
rect 11664 13744 11670 13796
rect 11146 13676 11152 13728
rect 11204 13676 11210 13728
rect 11808 13716 11836 13824
rect 11885 13821 11897 13855
rect 11931 13821 11943 13855
rect 11885 13815 11943 13821
rect 11977 13855 12035 13861
rect 11977 13821 11989 13855
rect 12023 13852 12035 13855
rect 12250 13852 12256 13864
rect 12023 13824 12256 13852
rect 12023 13821 12035 13824
rect 11977 13815 12035 13821
rect 11900 13784 11928 13815
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 13449 13855 13507 13861
rect 13449 13821 13461 13855
rect 13495 13852 13507 13855
rect 14384 13852 14412 13892
rect 14550 13880 14556 13892
rect 14608 13920 14614 13932
rect 15120 13920 15148 13960
rect 14608 13892 15148 13920
rect 14608 13880 14614 13892
rect 16758 13880 16764 13932
rect 16816 13920 16822 13932
rect 16853 13923 16911 13929
rect 16853 13920 16865 13923
rect 16816 13892 16865 13920
rect 16816 13880 16822 13892
rect 16853 13889 16865 13892
rect 16899 13889 16911 13923
rect 16853 13883 16911 13889
rect 17120 13923 17178 13929
rect 17120 13889 17132 13923
rect 17166 13920 17178 13923
rect 17402 13920 17408 13932
rect 17166 13892 17408 13920
rect 17166 13889 17178 13892
rect 17120 13883 17178 13889
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 17512 13920 17540 13960
rect 19061 13957 19073 13991
rect 19107 13957 19119 13991
rect 19061 13951 19119 13957
rect 19245 13991 19303 13997
rect 19245 13957 19257 13991
rect 19291 13988 19303 13991
rect 20346 13988 20352 14000
rect 19291 13960 20352 13988
rect 19291 13957 19303 13960
rect 19245 13951 19303 13957
rect 20346 13948 20352 13960
rect 20404 13948 20410 14000
rect 21468 13988 21496 14028
rect 22005 14025 22017 14028
rect 22051 14025 22063 14059
rect 22005 14019 22063 14025
rect 22370 14016 22376 14068
rect 22428 14016 22434 14068
rect 22462 14016 22468 14068
rect 22520 14016 22526 14068
rect 22554 14016 22560 14068
rect 22612 14056 22618 14068
rect 25958 14056 25964 14068
rect 22612 14028 25964 14056
rect 22612 14016 22618 14028
rect 25958 14016 25964 14028
rect 26016 14016 26022 14068
rect 26142 14016 26148 14068
rect 26200 14016 26206 14068
rect 28813 14059 28871 14065
rect 28813 14025 28825 14059
rect 28859 14056 28871 14059
rect 29086 14056 29092 14068
rect 28859 14028 29092 14056
rect 28859 14025 28871 14028
rect 28813 14019 28871 14025
rect 29086 14016 29092 14028
rect 29144 14016 29150 14068
rect 29362 14016 29368 14068
rect 29420 14016 29426 14068
rect 29914 14016 29920 14068
rect 29972 14056 29978 14068
rect 30834 14056 30840 14068
rect 29972 14028 30840 14056
rect 29972 14016 29978 14028
rect 30834 14016 30840 14028
rect 30892 14016 30898 14068
rect 32585 14059 32643 14065
rect 32585 14025 32597 14059
rect 32631 14056 32643 14059
rect 32858 14056 32864 14068
rect 32631 14028 32864 14056
rect 32631 14025 32643 14028
rect 32585 14019 32643 14025
rect 32858 14016 32864 14028
rect 32916 14016 32922 14068
rect 34885 14059 34943 14065
rect 34885 14025 34897 14059
rect 34931 14056 34943 14059
rect 36354 14056 36360 14068
rect 34931 14028 36360 14056
rect 34931 14025 34943 14028
rect 34885 14019 34943 14025
rect 36354 14016 36360 14028
rect 36412 14016 36418 14068
rect 37366 14016 37372 14068
rect 37424 14056 37430 14068
rect 37829 14059 37887 14065
rect 37829 14056 37841 14059
rect 37424 14028 37841 14056
rect 37424 14016 37430 14028
rect 37829 14025 37841 14028
rect 37875 14025 37887 14059
rect 37829 14019 37887 14025
rect 37918 14016 37924 14068
rect 37976 14056 37982 14068
rect 38013 14059 38071 14065
rect 38013 14056 38025 14059
rect 37976 14028 38025 14056
rect 37976 14016 37982 14028
rect 38013 14025 38025 14028
rect 38059 14056 38071 14059
rect 38059 14028 38654 14056
rect 38059 14025 38071 14028
rect 38013 14019 38071 14025
rect 31294 13988 31300 14000
rect 21192 13960 21496 13988
rect 23860 13960 31300 13988
rect 17512 13892 20116 13920
rect 13495 13824 14412 13852
rect 14461 13855 14519 13861
rect 13495 13821 13507 13824
rect 13449 13815 13507 13821
rect 14461 13821 14473 13855
rect 14507 13852 14519 13855
rect 14826 13852 14832 13864
rect 14507 13824 14832 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 14826 13812 14832 13824
rect 14884 13812 14890 13864
rect 15841 13855 15899 13861
rect 15841 13821 15853 13855
rect 15887 13852 15899 13855
rect 16022 13852 16028 13864
rect 15887 13824 16028 13852
rect 15887 13821 15899 13824
rect 15841 13815 15899 13821
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 19337 13855 19395 13861
rect 18248 13824 19288 13852
rect 12342 13784 12348 13796
rect 11900 13756 12348 13784
rect 12342 13744 12348 13756
rect 12400 13744 12406 13796
rect 16574 13784 16580 13796
rect 15396 13756 16580 13784
rect 12618 13716 12624 13728
rect 11808 13688 12624 13716
rect 12618 13676 12624 13688
rect 12676 13716 12682 13728
rect 15396 13716 15424 13756
rect 16574 13744 16580 13756
rect 16632 13744 16638 13796
rect 18248 13793 18276 13824
rect 18233 13787 18291 13793
rect 18233 13753 18245 13787
rect 18279 13753 18291 13787
rect 19260 13784 19288 13824
rect 19337 13821 19349 13855
rect 19383 13852 19395 13855
rect 19426 13852 19432 13864
rect 19383 13824 19432 13852
rect 19383 13821 19395 13824
rect 19337 13815 19395 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 20088 13852 20116 13892
rect 20162 13880 20168 13932
rect 20220 13920 20226 13932
rect 21192 13929 21220 13960
rect 20257 13923 20315 13929
rect 20257 13920 20269 13923
rect 20220 13892 20269 13920
rect 20220 13880 20226 13892
rect 20257 13889 20269 13892
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13889 21235 13923
rect 23860 13920 23888 13960
rect 31294 13948 31300 13960
rect 31352 13948 31358 14000
rect 34698 13988 34704 14000
rect 31404 13960 34704 13988
rect 21177 13883 21235 13889
rect 21275 13892 23888 13920
rect 20088 13824 20760 13852
rect 19518 13784 19524 13796
rect 19260 13756 19524 13784
rect 18233 13747 18291 13753
rect 19518 13744 19524 13756
rect 19576 13744 19582 13796
rect 19702 13744 19708 13796
rect 19760 13784 19766 13796
rect 20622 13784 20628 13796
rect 19760 13756 20628 13784
rect 19760 13744 19766 13756
rect 20622 13744 20628 13756
rect 20680 13744 20686 13796
rect 20732 13784 20760 13824
rect 20990 13812 20996 13864
rect 21048 13812 21054 13864
rect 21275 13784 21303 13892
rect 23934 13880 23940 13932
rect 23992 13920 23998 13932
rect 24210 13920 24216 13932
rect 23992 13892 24216 13920
rect 23992 13880 23998 13892
rect 24210 13880 24216 13892
rect 24268 13880 24274 13932
rect 24762 13880 24768 13932
rect 24820 13880 24826 13932
rect 24946 13880 24952 13932
rect 25004 13880 25010 13932
rect 25038 13880 25044 13932
rect 25096 13880 25102 13932
rect 25222 13880 25228 13932
rect 25280 13880 25286 13932
rect 25317 13923 25375 13929
rect 25317 13889 25329 13923
rect 25363 13920 25375 13923
rect 25498 13920 25504 13932
rect 25363 13892 25504 13920
rect 25363 13889 25375 13892
rect 25317 13883 25375 13889
rect 25498 13880 25504 13892
rect 25556 13880 25562 13932
rect 25958 13880 25964 13932
rect 26016 13920 26022 13932
rect 28721 13923 28779 13929
rect 26016 13892 28672 13920
rect 26016 13880 26022 13892
rect 22557 13855 22615 13861
rect 22557 13821 22569 13855
rect 22603 13821 22615 13855
rect 24964 13852 24992 13880
rect 25866 13852 25872 13864
rect 24964 13824 25872 13852
rect 22557 13815 22615 13821
rect 20732 13756 21303 13784
rect 22572 13784 22600 13815
rect 25866 13812 25872 13824
rect 25924 13812 25930 13864
rect 26142 13812 26148 13864
rect 26200 13852 26206 13864
rect 26237 13855 26295 13861
rect 26237 13852 26249 13855
rect 26200 13824 26249 13852
rect 26200 13812 26206 13824
rect 26237 13821 26249 13824
rect 26283 13821 26295 13855
rect 26237 13815 26295 13821
rect 26421 13855 26479 13861
rect 26421 13821 26433 13855
rect 26467 13852 26479 13855
rect 28166 13852 28172 13864
rect 26467 13824 28172 13852
rect 26467 13821 26479 13824
rect 26421 13815 26479 13821
rect 28166 13812 28172 13824
rect 28224 13812 28230 13864
rect 28644 13852 28672 13892
rect 28721 13889 28733 13923
rect 28767 13920 28779 13923
rect 28810 13920 28816 13932
rect 28767 13892 28816 13920
rect 28767 13889 28779 13892
rect 28721 13883 28779 13889
rect 28810 13880 28816 13892
rect 28868 13920 28874 13932
rect 29546 13920 29552 13932
rect 28868 13892 29552 13920
rect 28868 13880 28874 13892
rect 29546 13880 29552 13892
rect 29604 13880 29610 13932
rect 29733 13923 29791 13929
rect 29733 13889 29745 13923
rect 29779 13920 29791 13923
rect 31018 13920 31024 13932
rect 29779 13892 31024 13920
rect 29779 13889 29791 13892
rect 29733 13883 29791 13889
rect 29748 13852 29776 13883
rect 31018 13880 31024 13892
rect 31076 13880 31082 13932
rect 31205 13923 31263 13929
rect 31205 13889 31217 13923
rect 31251 13920 31263 13923
rect 31404 13920 31432 13960
rect 34698 13948 34704 13960
rect 34756 13948 34762 14000
rect 37550 13948 37556 14000
rect 37608 13988 37614 14000
rect 38626 13988 38654 14028
rect 39022 14016 39028 14068
rect 39080 14016 39086 14068
rect 42061 14059 42119 14065
rect 42061 14025 42073 14059
rect 42107 14056 42119 14059
rect 42978 14056 42984 14068
rect 42107 14028 42984 14056
rect 42107 14025 42119 14028
rect 42061 14019 42119 14025
rect 42978 14016 42984 14028
rect 43036 14016 43042 14068
rect 43990 14016 43996 14068
rect 44048 14056 44054 14068
rect 56686 14056 56692 14068
rect 44048 14028 56692 14056
rect 44048 14016 44054 14028
rect 56686 14016 56692 14028
rect 56744 14016 56750 14068
rect 41322 13988 41328 14000
rect 37608 13960 38148 13988
rect 38626 13960 41328 13988
rect 37608 13948 37614 13960
rect 31251 13892 31432 13920
rect 31251 13889 31263 13892
rect 31205 13883 31263 13889
rect 31570 13880 31576 13932
rect 31628 13880 31634 13932
rect 31754 13880 31760 13932
rect 31812 13880 31818 13932
rect 31938 13880 31944 13932
rect 31996 13920 32002 13932
rect 32309 13923 32367 13929
rect 32309 13920 32321 13923
rect 31996 13892 32321 13920
rect 31996 13880 32002 13892
rect 32309 13889 32321 13892
rect 32355 13889 32367 13923
rect 32309 13883 32367 13889
rect 32490 13880 32496 13932
rect 32548 13920 32554 13932
rect 32769 13923 32827 13929
rect 32769 13920 32781 13923
rect 32548 13892 32781 13920
rect 32548 13880 32554 13892
rect 32769 13889 32781 13892
rect 32815 13889 32827 13923
rect 36722 13920 36728 13932
rect 32769 13883 32827 13889
rect 32876 13892 36728 13920
rect 28644 13824 29776 13852
rect 29822 13812 29828 13864
rect 29880 13812 29886 13864
rect 30009 13855 30067 13861
rect 30009 13821 30021 13855
rect 30055 13821 30067 13855
rect 30009 13815 30067 13821
rect 25130 13784 25136 13796
rect 22572 13756 25136 13784
rect 12676 13688 15424 13716
rect 12676 13676 12682 13688
rect 15470 13676 15476 13728
rect 15528 13716 15534 13728
rect 18414 13716 18420 13728
rect 15528 13688 18420 13716
rect 15528 13676 15534 13688
rect 18414 13676 18420 13688
rect 18472 13676 18478 13728
rect 19610 13676 19616 13728
rect 19668 13716 19674 13728
rect 20441 13719 20499 13725
rect 20441 13716 20453 13719
rect 19668 13688 20453 13716
rect 19668 13676 19674 13688
rect 20441 13685 20453 13688
rect 20487 13685 20499 13719
rect 20441 13679 20499 13685
rect 21266 13676 21272 13728
rect 21324 13716 21330 13728
rect 21361 13719 21419 13725
rect 21361 13716 21373 13719
rect 21324 13688 21373 13716
rect 21324 13676 21330 13688
rect 21361 13685 21373 13688
rect 21407 13685 21419 13719
rect 21361 13679 21419 13685
rect 21450 13676 21456 13728
rect 21508 13716 21514 13728
rect 22572 13716 22600 13756
rect 25130 13744 25136 13756
rect 25188 13744 25194 13796
rect 29454 13744 29460 13796
rect 29512 13784 29518 13796
rect 30024 13784 30052 13815
rect 30374 13812 30380 13864
rect 30432 13852 30438 13864
rect 30558 13852 30564 13864
rect 30432 13824 30564 13852
rect 30432 13812 30438 13824
rect 30558 13812 30564 13824
rect 30616 13812 30622 13864
rect 30834 13812 30840 13864
rect 30892 13852 30898 13864
rect 31113 13855 31171 13861
rect 31113 13852 31125 13855
rect 30892 13824 31125 13852
rect 30892 13812 30898 13824
rect 31113 13821 31125 13824
rect 31159 13821 31171 13855
rect 31772 13852 31800 13880
rect 32876 13852 32904 13892
rect 36722 13880 36728 13892
rect 36780 13880 36786 13932
rect 38010 13920 38016 13932
rect 37971 13892 38016 13920
rect 38010 13880 38016 13892
rect 38068 13880 38074 13932
rect 38120 13920 38148 13960
rect 41322 13948 41328 13960
rect 41380 13948 41386 14000
rect 46198 13948 46204 14000
rect 46256 13988 46262 14000
rect 57790 13988 57796 14000
rect 46256 13960 57796 13988
rect 46256 13948 46262 13960
rect 57790 13948 57796 13960
rect 57848 13948 57854 14000
rect 38654 13920 38660 13932
rect 38120 13892 38660 13920
rect 38654 13880 38660 13892
rect 38712 13880 38718 13932
rect 38930 13880 38936 13932
rect 38988 13880 38994 13932
rect 39117 13923 39175 13929
rect 39117 13889 39129 13923
rect 39163 13889 39175 13923
rect 39117 13883 39175 13889
rect 31772 13824 32904 13852
rect 31113 13815 31171 13821
rect 34790 13812 34796 13864
rect 34848 13852 34854 13864
rect 34977 13855 35035 13861
rect 34977 13852 34989 13855
rect 34848 13824 34989 13852
rect 34848 13812 34854 13824
rect 34977 13821 34989 13824
rect 35023 13821 35035 13855
rect 34977 13815 35035 13821
rect 35161 13855 35219 13861
rect 35161 13821 35173 13855
rect 35207 13852 35219 13855
rect 35342 13852 35348 13864
rect 35207 13824 35348 13852
rect 35207 13821 35219 13824
rect 35161 13815 35219 13821
rect 35342 13812 35348 13824
rect 35400 13852 35406 13864
rect 35710 13852 35716 13864
rect 35400 13824 35716 13852
rect 35400 13812 35406 13824
rect 35710 13812 35716 13824
rect 35768 13812 35774 13864
rect 38473 13855 38531 13861
rect 38473 13821 38485 13855
rect 38519 13852 38531 13855
rect 38746 13852 38752 13864
rect 38519 13824 38752 13852
rect 38519 13821 38531 13824
rect 38473 13815 38531 13821
rect 38746 13812 38752 13824
rect 38804 13812 38810 13864
rect 39132 13852 39160 13883
rect 40494 13880 40500 13932
rect 40552 13920 40558 13932
rect 41509 13923 41567 13929
rect 41509 13920 41521 13923
rect 40552 13892 41521 13920
rect 40552 13880 40558 13892
rect 41509 13889 41521 13892
rect 41555 13889 41567 13923
rect 41509 13883 41567 13889
rect 41690 13880 41696 13932
rect 41748 13880 41754 13932
rect 41782 13880 41788 13932
rect 41840 13880 41846 13932
rect 41877 13923 41935 13929
rect 41877 13889 41889 13923
rect 41923 13889 41935 13923
rect 41877 13883 41935 13889
rect 41414 13852 41420 13864
rect 39132 13824 41420 13852
rect 41414 13812 41420 13824
rect 41472 13812 41478 13864
rect 41892 13852 41920 13883
rect 43070 13880 43076 13932
rect 43128 13880 43134 13932
rect 41520 13824 41920 13852
rect 30926 13784 30932 13796
rect 29512 13756 30932 13784
rect 29512 13744 29518 13756
rect 30926 13744 30932 13756
rect 30984 13744 30990 13796
rect 38381 13787 38439 13793
rect 38381 13784 38393 13787
rect 31726 13756 38393 13784
rect 21508 13688 22600 13716
rect 21508 13676 21514 13688
rect 25774 13676 25780 13728
rect 25832 13676 25838 13728
rect 26050 13676 26056 13728
rect 26108 13716 26114 13728
rect 31726 13716 31754 13756
rect 38381 13753 38393 13756
rect 38427 13753 38439 13787
rect 41520 13784 41548 13824
rect 43346 13812 43352 13864
rect 43404 13812 43410 13864
rect 43530 13812 43536 13864
rect 43588 13852 43594 13864
rect 44729 13855 44787 13861
rect 44729 13852 44741 13855
rect 43588 13824 44741 13852
rect 43588 13812 43594 13824
rect 44729 13821 44741 13824
rect 44775 13852 44787 13855
rect 57514 13852 57520 13864
rect 44775 13824 57520 13852
rect 44775 13821 44787 13824
rect 44729 13815 44787 13821
rect 57514 13812 57520 13824
rect 57572 13812 57578 13864
rect 38381 13747 38439 13753
rect 38488 13756 41548 13784
rect 26108 13688 31754 13716
rect 26108 13676 26114 13688
rect 31846 13676 31852 13728
rect 31904 13716 31910 13728
rect 33502 13716 33508 13728
rect 31904 13688 33508 13716
rect 31904 13676 31910 13688
rect 33502 13676 33508 13688
rect 33560 13676 33566 13728
rect 34514 13676 34520 13728
rect 34572 13676 34578 13728
rect 37274 13676 37280 13728
rect 37332 13716 37338 13728
rect 38488 13716 38516 13756
rect 37332 13688 38516 13716
rect 37332 13676 37338 13688
rect 41322 13676 41328 13728
rect 41380 13716 41386 13728
rect 42518 13716 42524 13728
rect 41380 13688 42524 13716
rect 41380 13676 41386 13688
rect 42518 13676 42524 13688
rect 42576 13716 42582 13728
rect 44450 13716 44456 13728
rect 42576 13688 44456 13716
rect 42576 13676 42582 13688
rect 44450 13676 44456 13688
rect 44508 13676 44514 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 9858 13472 9864 13524
rect 9916 13472 9922 13524
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10873 13515 10931 13521
rect 10873 13512 10885 13515
rect 10192 13484 10885 13512
rect 10192 13472 10198 13484
rect 10873 13481 10885 13484
rect 10919 13481 10931 13515
rect 10873 13475 10931 13481
rect 13633 13515 13691 13521
rect 13633 13481 13645 13515
rect 13679 13512 13691 13515
rect 14274 13512 14280 13524
rect 13679 13484 14280 13512
rect 13679 13481 13691 13484
rect 13633 13475 13691 13481
rect 14274 13472 14280 13484
rect 14332 13472 14338 13524
rect 15013 13515 15071 13521
rect 15013 13481 15025 13515
rect 15059 13512 15071 13515
rect 15746 13512 15752 13524
rect 15059 13484 15752 13512
rect 15059 13481 15071 13484
rect 15013 13475 15071 13481
rect 15746 13472 15752 13484
rect 15804 13472 15810 13524
rect 16500 13484 22324 13512
rect 14461 13447 14519 13453
rect 14461 13413 14473 13447
rect 14507 13444 14519 13447
rect 16301 13447 16359 13453
rect 16301 13444 16313 13447
rect 14507 13416 16313 13444
rect 14507 13413 14519 13416
rect 14461 13407 14519 13413
rect 16301 13413 16313 13416
rect 16347 13413 16359 13447
rect 16301 13407 16359 13413
rect 11885 13379 11943 13385
rect 11885 13345 11897 13379
rect 11931 13376 11943 13379
rect 13722 13376 13728 13388
rect 11931 13348 13728 13376
rect 11931 13345 11943 13348
rect 11885 13339 11943 13345
rect 13722 13336 13728 13348
rect 13780 13336 13786 13388
rect 15197 13379 15255 13385
rect 15197 13345 15209 13379
rect 15243 13376 15255 13379
rect 16500 13376 16528 13484
rect 16574 13404 16580 13456
rect 16632 13444 16638 13456
rect 18506 13444 18512 13456
rect 16632 13416 18512 13444
rect 16632 13404 16638 13416
rect 18506 13404 18512 13416
rect 18564 13444 18570 13456
rect 18874 13444 18880 13456
rect 18564 13416 18880 13444
rect 18564 13404 18570 13416
rect 18874 13404 18880 13416
rect 18932 13404 18938 13456
rect 19613 13447 19671 13453
rect 19613 13413 19625 13447
rect 19659 13444 19671 13447
rect 20254 13444 20260 13456
rect 19659 13416 20260 13444
rect 19659 13413 19671 13416
rect 19613 13407 19671 13413
rect 20254 13404 20260 13416
rect 20312 13404 20318 13456
rect 20898 13444 20904 13456
rect 20732 13416 20904 13444
rect 15243 13348 16528 13376
rect 15243 13345 15255 13348
rect 15197 13339 15255 13345
rect 17310 13336 17316 13388
rect 17368 13376 17374 13388
rect 17770 13376 17776 13388
rect 17368 13348 17776 13376
rect 17368 13336 17374 13348
rect 17770 13336 17776 13348
rect 17828 13336 17834 13388
rect 19334 13376 19340 13388
rect 18248 13348 19340 13376
rect 1578 13268 1584 13320
rect 1636 13268 1642 13320
rect 9674 13268 9680 13320
rect 9732 13268 9738 13320
rect 10612 13280 12296 13308
rect 10612 13252 10640 13280
rect 934 13200 940 13252
rect 992 13240 998 13252
rect 1857 13243 1915 13249
rect 1857 13240 1869 13243
rect 992 13212 1869 13240
rect 992 13200 998 13212
rect 1857 13209 1869 13212
rect 1903 13209 1915 13243
rect 1857 13203 1915 13209
rect 10505 13243 10563 13249
rect 10505 13209 10517 13243
rect 10551 13240 10563 13243
rect 10594 13240 10600 13252
rect 10551 13212 10600 13240
rect 10551 13209 10563 13212
rect 10505 13203 10563 13209
rect 10594 13200 10600 13212
rect 10652 13200 10658 13252
rect 10686 13200 10692 13252
rect 10744 13200 10750 13252
rect 12268 13249 12296 13280
rect 12618 13268 12624 13320
rect 12676 13268 12682 13320
rect 13446 13268 13452 13320
rect 13504 13268 13510 13320
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 15102 13308 15108 13320
rect 14323 13280 15108 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 15286 13268 15292 13320
rect 15344 13268 15350 13320
rect 15378 13268 15384 13320
rect 15436 13268 15442 13320
rect 15470 13268 15476 13320
rect 15528 13268 15534 13320
rect 18248 13317 18276 13348
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 20165 13379 20223 13385
rect 20165 13345 20177 13379
rect 20211 13376 20223 13379
rect 20732 13376 20760 13416
rect 20898 13404 20904 13416
rect 20956 13404 20962 13456
rect 22296 13444 22324 13484
rect 22370 13472 22376 13524
rect 22428 13472 22434 13524
rect 24578 13472 24584 13524
rect 24636 13512 24642 13524
rect 27341 13515 27399 13521
rect 27341 13512 27353 13515
rect 24636 13484 27353 13512
rect 24636 13472 24642 13484
rect 27341 13481 27353 13484
rect 27387 13512 27399 13515
rect 27522 13512 27528 13524
rect 27387 13484 27528 13512
rect 27387 13481 27399 13484
rect 27341 13475 27399 13481
rect 27522 13472 27528 13484
rect 27580 13472 27586 13524
rect 27706 13472 27712 13524
rect 27764 13512 27770 13524
rect 30834 13512 30840 13524
rect 27764 13484 30840 13512
rect 27764 13472 27770 13484
rect 30834 13472 30840 13484
rect 30892 13472 30898 13524
rect 32493 13515 32551 13521
rect 31588 13484 32076 13512
rect 24026 13444 24032 13456
rect 22296 13416 24032 13444
rect 24026 13404 24032 13416
rect 24084 13444 24090 13456
rect 28810 13444 28816 13456
rect 24084 13416 28816 13444
rect 24084 13404 24090 13416
rect 28810 13404 28816 13416
rect 28868 13404 28874 13456
rect 20211 13348 20760 13376
rect 20211 13345 20223 13348
rect 20165 13339 20223 13345
rect 20272 13320 20300 13348
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 20990 13376 20996 13388
rect 20864 13348 20996 13376
rect 20864 13336 20870 13348
rect 20990 13336 20996 13348
rect 21048 13336 21054 13388
rect 24670 13336 24676 13388
rect 24728 13376 24734 13388
rect 26326 13376 26332 13388
rect 24728 13348 26332 13376
rect 24728 13336 24734 13348
rect 26326 13336 26332 13348
rect 26384 13336 26390 13388
rect 16025 13311 16083 13317
rect 16025 13308 16037 13311
rect 15580 13280 16037 13308
rect 12253 13243 12311 13249
rect 12253 13209 12265 13243
rect 12299 13240 12311 13243
rect 12342 13240 12348 13252
rect 12299 13212 12348 13240
rect 12299 13209 12311 13212
rect 12253 13203 12311 13209
rect 12342 13200 12348 13212
rect 12400 13240 12406 13252
rect 12400 13200 12434 13240
rect 11974 13132 11980 13184
rect 12032 13172 12038 13184
rect 12069 13175 12127 13181
rect 12069 13172 12081 13175
rect 12032 13144 12081 13172
rect 12032 13132 12038 13144
rect 12069 13141 12081 13144
rect 12115 13141 12127 13175
rect 12069 13135 12127 13141
rect 12158 13132 12164 13184
rect 12216 13132 12222 13184
rect 12406 13172 12434 13200
rect 15194 13172 15200 13184
rect 12406 13144 15200 13172
rect 15194 13132 15200 13144
rect 15252 13172 15258 13184
rect 15580 13172 15608 13280
rect 16025 13277 16037 13280
rect 16071 13277 16083 13311
rect 16025 13271 16083 13277
rect 17221 13311 17279 13317
rect 17221 13277 17233 13311
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 18233 13311 18291 13317
rect 18233 13277 18245 13311
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 17236 13240 17264 13271
rect 18414 13268 18420 13320
rect 18472 13268 18478 13320
rect 18506 13268 18512 13320
rect 18564 13268 18570 13320
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13308 19487 13311
rect 19610 13308 19616 13320
rect 19475 13280 19616 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 19610 13268 19616 13280
rect 19668 13268 19674 13320
rect 20254 13268 20260 13320
rect 20312 13268 20318 13320
rect 20349 13311 20407 13317
rect 20349 13277 20361 13311
rect 20395 13308 20407 13311
rect 20714 13308 20720 13320
rect 20395 13280 20720 13308
rect 20395 13277 20407 13280
rect 20349 13271 20407 13277
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 21266 13317 21272 13320
rect 21260 13308 21272 13317
rect 21227 13280 21272 13308
rect 21260 13271 21272 13280
rect 21266 13268 21272 13271
rect 21324 13268 21330 13320
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13308 24823 13311
rect 24854 13308 24860 13320
rect 24811 13280 24860 13308
rect 24811 13277 24823 13280
rect 24765 13271 24823 13277
rect 24854 13268 24860 13280
rect 24912 13268 24918 13320
rect 28534 13308 28540 13320
rect 24964 13280 28540 13308
rect 19702 13240 19708 13252
rect 17236 13212 19708 13240
rect 19702 13200 19708 13212
rect 19760 13200 19766 13252
rect 20898 13200 20904 13252
rect 20956 13240 20962 13252
rect 23566 13240 23572 13252
rect 20956 13212 23572 13240
rect 20956 13200 20962 13212
rect 23566 13200 23572 13212
rect 23624 13200 23630 13252
rect 24964 13240 24992 13280
rect 28534 13268 28540 13280
rect 28592 13268 28598 13320
rect 30098 13268 30104 13320
rect 30156 13308 30162 13320
rect 31588 13317 31616 13484
rect 31938 13444 31944 13456
rect 31680 13416 31944 13444
rect 30837 13311 30895 13317
rect 30837 13308 30849 13311
rect 30156 13280 30849 13308
rect 30156 13268 30162 13280
rect 30837 13277 30849 13280
rect 30883 13308 30895 13311
rect 31573 13311 31631 13317
rect 30883 13280 31524 13308
rect 30883 13277 30895 13280
rect 30837 13271 30895 13277
rect 23667 13212 24992 13240
rect 26053 13243 26111 13249
rect 15252 13144 15608 13172
rect 15252 13132 15258 13144
rect 15838 13132 15844 13184
rect 15896 13172 15902 13184
rect 16485 13175 16543 13181
rect 16485 13172 16497 13175
rect 15896 13144 16497 13172
rect 15896 13132 15902 13144
rect 16485 13141 16497 13144
rect 16531 13141 16543 13175
rect 16485 13135 16543 13141
rect 16942 13132 16948 13184
rect 17000 13172 17006 13184
rect 17589 13175 17647 13181
rect 17589 13172 17601 13175
rect 17000 13144 17601 13172
rect 17000 13132 17006 13144
rect 17589 13141 17601 13144
rect 17635 13141 17647 13175
rect 17589 13135 17647 13141
rect 18049 13175 18107 13181
rect 18049 13141 18061 13175
rect 18095 13172 18107 13175
rect 18138 13172 18144 13184
rect 18095 13144 18144 13172
rect 18095 13141 18107 13144
rect 18049 13135 18107 13141
rect 18138 13132 18144 13144
rect 18196 13132 18202 13184
rect 20533 13175 20591 13181
rect 20533 13141 20545 13175
rect 20579 13172 20591 13175
rect 21082 13172 21088 13184
rect 20579 13144 21088 13172
rect 20579 13141 20591 13144
rect 20533 13135 20591 13141
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 21910 13132 21916 13184
rect 21968 13172 21974 13184
rect 23667 13172 23695 13212
rect 26053 13209 26065 13243
rect 26099 13240 26111 13243
rect 28626 13240 28632 13252
rect 26099 13212 28632 13240
rect 26099 13209 26111 13212
rect 26053 13203 26111 13209
rect 28626 13200 28632 13212
rect 28684 13200 28690 13252
rect 31113 13243 31171 13249
rect 31113 13209 31125 13243
rect 31159 13240 31171 13243
rect 31386 13240 31392 13252
rect 31159 13212 31392 13240
rect 31159 13209 31171 13212
rect 31113 13203 31171 13209
rect 31386 13200 31392 13212
rect 31444 13200 31450 13252
rect 31496 13240 31524 13280
rect 31573 13277 31585 13311
rect 31619 13277 31631 13311
rect 31573 13271 31631 13277
rect 31680 13240 31708 13416
rect 31938 13404 31944 13416
rect 31996 13404 32002 13456
rect 31846 13336 31852 13388
rect 31904 13336 31910 13388
rect 32048 13376 32076 13484
rect 32493 13481 32505 13515
rect 32539 13512 32551 13515
rect 32582 13512 32588 13524
rect 32539 13484 32588 13512
rect 32539 13481 32551 13484
rect 32493 13475 32551 13481
rect 32582 13472 32588 13484
rect 32640 13512 32646 13524
rect 32769 13515 32827 13521
rect 32769 13512 32781 13515
rect 32640 13484 32781 13512
rect 32640 13472 32646 13484
rect 32769 13481 32781 13484
rect 32815 13481 32827 13515
rect 32769 13475 32827 13481
rect 38010 13472 38016 13524
rect 38068 13512 38074 13524
rect 38068 13484 41414 13512
rect 38068 13472 38074 13484
rect 32125 13447 32183 13453
rect 32125 13413 32137 13447
rect 32171 13444 32183 13447
rect 32171 13416 32904 13444
rect 32171 13413 32183 13416
rect 32125 13407 32183 13413
rect 32876 13385 32904 13416
rect 33594 13404 33600 13456
rect 33652 13444 33658 13456
rect 38838 13444 38844 13456
rect 33652 13416 38844 13444
rect 33652 13404 33658 13416
rect 38838 13404 38844 13416
rect 38896 13404 38902 13456
rect 41386 13444 41414 13484
rect 43254 13472 43260 13524
rect 43312 13512 43318 13524
rect 43533 13515 43591 13521
rect 43533 13512 43545 13515
rect 43312 13484 43545 13512
rect 43312 13472 43318 13484
rect 43533 13481 43545 13484
rect 43579 13481 43591 13515
rect 43533 13475 43591 13481
rect 57330 13444 57336 13456
rect 41386 13416 57336 13444
rect 57330 13404 57336 13416
rect 57388 13404 57394 13456
rect 32861 13379 32919 13385
rect 32048 13348 32536 13376
rect 31864 13308 31892 13336
rect 31941 13311 31999 13317
rect 31941 13308 31953 13311
rect 31864 13280 31953 13308
rect 31941 13277 31953 13280
rect 31987 13308 31999 13311
rect 32398 13308 32404 13320
rect 31987 13280 32404 13308
rect 31987 13277 31999 13280
rect 31941 13271 31999 13277
rect 32398 13268 32404 13280
rect 32456 13268 32462 13320
rect 32508 13308 32536 13348
rect 32861 13345 32873 13379
rect 32907 13345 32919 13379
rect 35986 13376 35992 13388
rect 32861 13339 32919 13345
rect 32968 13348 35992 13376
rect 32968 13308 32996 13348
rect 35986 13336 35992 13348
rect 36044 13336 36050 13388
rect 36078 13336 36084 13388
rect 36136 13376 36142 13388
rect 38657 13379 38715 13385
rect 38657 13376 38669 13379
rect 36136 13348 38669 13376
rect 36136 13336 36142 13348
rect 38657 13345 38669 13348
rect 38703 13376 38715 13379
rect 41690 13376 41696 13388
rect 38703 13348 41696 13376
rect 38703 13345 38715 13348
rect 38657 13339 38715 13345
rect 41690 13336 41696 13348
rect 41748 13376 41754 13388
rect 44542 13376 44548 13388
rect 41748 13348 42380 13376
rect 41748 13336 41754 13348
rect 32508 13280 32996 13308
rect 33042 13268 33048 13320
rect 33100 13268 33106 13320
rect 36357 13311 36415 13317
rect 36357 13277 36369 13311
rect 36403 13277 36415 13311
rect 36357 13271 36415 13277
rect 31496 13212 31708 13240
rect 31757 13243 31815 13249
rect 31757 13209 31769 13243
rect 31803 13209 31815 13243
rect 31757 13203 31815 13209
rect 21968 13144 23695 13172
rect 24857 13175 24915 13181
rect 21968 13132 21974 13144
rect 24857 13141 24869 13175
rect 24903 13172 24915 13175
rect 24946 13172 24952 13184
rect 24903 13144 24952 13172
rect 24903 13141 24915 13144
rect 24857 13135 24915 13141
rect 24946 13132 24952 13144
rect 25004 13132 25010 13184
rect 31772 13172 31800 13203
rect 31846 13200 31852 13252
rect 31904 13200 31910 13252
rect 32769 13243 32827 13249
rect 32769 13209 32781 13243
rect 32815 13240 32827 13243
rect 35802 13240 35808 13252
rect 32815 13212 35808 13240
rect 32815 13209 32827 13212
rect 32769 13203 32827 13209
rect 35802 13200 35808 13212
rect 35860 13200 35866 13252
rect 36372 13240 36400 13271
rect 36446 13268 36452 13320
rect 36504 13268 36510 13320
rect 38286 13268 38292 13320
rect 38344 13268 38350 13320
rect 38746 13268 38752 13320
rect 38804 13308 38810 13320
rect 39114 13308 39120 13320
rect 38804 13280 39120 13308
rect 38804 13268 38810 13280
rect 39114 13268 39120 13280
rect 39172 13268 39178 13320
rect 42352 13317 42380 13348
rect 42444 13348 44548 13376
rect 42444 13317 42472 13348
rect 44542 13336 44548 13348
rect 44600 13336 44606 13388
rect 58158 13336 58164 13388
rect 58216 13336 58222 13388
rect 42153 13311 42211 13317
rect 42153 13277 42165 13311
rect 42199 13277 42211 13311
rect 42153 13271 42211 13277
rect 42337 13311 42395 13317
rect 42337 13277 42349 13311
rect 42383 13277 42395 13311
rect 42337 13271 42395 13277
rect 42429 13311 42487 13317
rect 42429 13277 42441 13311
rect 42475 13277 42487 13311
rect 42429 13271 42487 13277
rect 41966 13240 41972 13252
rect 36372 13212 41972 13240
rect 41966 13200 41972 13212
rect 42024 13200 42030 13252
rect 31938 13172 31944 13184
rect 31772 13144 31944 13172
rect 31938 13132 31944 13144
rect 31996 13132 32002 13184
rect 32582 13132 32588 13184
rect 32640 13172 32646 13184
rect 33229 13175 33287 13181
rect 33229 13172 33241 13175
rect 32640 13144 33241 13172
rect 32640 13132 32646 13144
rect 33229 13141 33241 13144
rect 33275 13141 33287 13175
rect 33229 13135 33287 13141
rect 36630 13132 36636 13184
rect 36688 13132 36694 13184
rect 42168 13172 42196 13271
rect 42518 13268 42524 13320
rect 42576 13268 42582 13320
rect 42702 13268 42708 13320
rect 42760 13308 42766 13320
rect 43165 13311 43223 13317
rect 43165 13308 43177 13311
rect 42760 13280 43177 13308
rect 42760 13268 42766 13280
rect 43165 13277 43177 13280
rect 43211 13277 43223 13311
rect 43165 13271 43223 13277
rect 43349 13311 43407 13317
rect 43349 13277 43361 13311
rect 43395 13277 43407 13311
rect 43349 13271 43407 13277
rect 43364 13240 43392 13271
rect 46566 13268 46572 13320
rect 46624 13308 46630 13320
rect 57885 13311 57943 13317
rect 57885 13308 57897 13311
rect 46624 13280 57897 13308
rect 46624 13268 46630 13280
rect 57885 13277 57897 13280
rect 57931 13277 57943 13311
rect 57885 13271 57943 13277
rect 42720 13212 43392 13240
rect 57057 13243 57115 13249
rect 42518 13172 42524 13184
rect 42168 13144 42524 13172
rect 42518 13132 42524 13144
rect 42576 13132 42582 13184
rect 42720 13181 42748 13212
rect 57057 13209 57069 13243
rect 57103 13240 57115 13243
rect 58986 13240 58992 13252
rect 57103 13212 58992 13240
rect 57103 13209 57115 13212
rect 57057 13203 57115 13209
rect 58986 13200 58992 13212
rect 59044 13200 59050 13252
rect 42705 13175 42763 13181
rect 42705 13141 42717 13175
rect 42751 13141 42763 13175
rect 42705 13135 42763 13141
rect 57146 13132 57152 13184
rect 57204 13132 57210 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 10689 12971 10747 12977
rect 10689 12968 10701 12971
rect 9824 12940 10701 12968
rect 9824 12928 9830 12940
rect 10689 12937 10701 12940
rect 10735 12937 10747 12971
rect 10689 12931 10747 12937
rect 11882 12928 11888 12980
rect 11940 12928 11946 12980
rect 13998 12928 14004 12980
rect 14056 12928 14062 12980
rect 15194 12928 15200 12980
rect 15252 12928 15258 12980
rect 15470 12928 15476 12980
rect 15528 12968 15534 12980
rect 15528 12940 19196 12968
rect 15528 12928 15534 12940
rect 14550 12860 14556 12912
rect 14608 12860 14614 12912
rect 14921 12903 14979 12909
rect 14921 12869 14933 12903
rect 14967 12900 14979 12903
rect 15378 12900 15384 12912
rect 14967 12872 15384 12900
rect 14967 12869 14979 12872
rect 14921 12863 14979 12869
rect 15378 12860 15384 12872
rect 15436 12860 15442 12912
rect 17681 12903 17739 12909
rect 17681 12900 17693 12903
rect 16046 12872 17693 12900
rect 10502 12792 10508 12844
rect 10560 12792 10566 12844
rect 11146 12792 11152 12844
rect 11204 12832 11210 12844
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 11204 12804 11713 12832
rect 11204 12792 11210 12804
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 12434 12792 12440 12844
rect 12492 12792 12498 12844
rect 13814 12792 13820 12844
rect 13872 12792 13878 12844
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15102 12832 15108 12844
rect 14875 12804 15108 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 16046 12841 16074 12872
rect 17681 12869 17693 12872
rect 17727 12869 17739 12903
rect 17681 12863 17739 12869
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 17310 12792 17316 12844
rect 17368 12792 17374 12844
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12832 17555 12835
rect 18046 12832 18052 12844
rect 17543 12804 18052 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 18138 12792 18144 12844
rect 18196 12792 18202 12844
rect 15013 12767 15071 12773
rect 15013 12733 15025 12767
rect 15059 12764 15071 12767
rect 19168 12764 19196 12940
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19429 12971 19487 12977
rect 19429 12968 19441 12971
rect 19392 12940 19441 12968
rect 19392 12928 19398 12940
rect 19429 12937 19441 12940
rect 19475 12937 19487 12971
rect 19429 12931 19487 12937
rect 20165 12971 20223 12977
rect 20165 12937 20177 12971
rect 20211 12937 20223 12971
rect 20165 12931 20223 12937
rect 20180 12900 20208 12931
rect 20714 12928 20720 12980
rect 20772 12928 20778 12980
rect 22925 12971 22983 12977
rect 22925 12968 22937 12971
rect 20916 12940 22937 12968
rect 19720 12872 20208 12900
rect 19270 12835 19328 12841
rect 19270 12801 19282 12835
rect 19316 12832 19328 12835
rect 19720 12832 19748 12872
rect 19316 12804 19748 12832
rect 19981 12835 20039 12841
rect 19316 12801 19328 12804
rect 19270 12795 19328 12801
rect 19981 12801 19993 12835
rect 20027 12832 20039 12835
rect 20916 12832 20944 12940
rect 22925 12937 22937 12940
rect 22971 12937 22983 12971
rect 22925 12931 22983 12937
rect 23382 12928 23388 12980
rect 23440 12968 23446 12980
rect 27341 12971 27399 12977
rect 23440 12940 25912 12968
rect 23440 12928 23446 12940
rect 20990 12860 20996 12912
rect 21048 12900 21054 12912
rect 24578 12900 24584 12912
rect 21048 12872 24584 12900
rect 21048 12860 21054 12872
rect 24578 12860 24584 12872
rect 24636 12900 24642 12912
rect 25124 12903 25182 12909
rect 24636 12872 24900 12900
rect 24636 12860 24642 12872
rect 20027 12804 20944 12832
rect 21085 12835 21143 12841
rect 20027 12801 20039 12804
rect 19981 12795 20039 12801
rect 21085 12801 21097 12835
rect 21131 12832 21143 12835
rect 21634 12832 21640 12844
rect 21131 12804 21640 12832
rect 21131 12801 21143 12804
rect 21085 12795 21143 12801
rect 21634 12792 21640 12804
rect 21692 12792 21698 12844
rect 22005 12835 22063 12841
rect 22005 12801 22017 12835
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 15059 12736 19012 12764
rect 19168 12736 19334 12764
rect 15059 12733 15071 12736
rect 15013 12727 15071 12733
rect 15378 12656 15384 12708
rect 15436 12696 15442 12708
rect 18230 12696 18236 12708
rect 15436 12668 18236 12696
rect 15436 12656 15442 12668
rect 18230 12656 18236 12668
rect 18288 12656 18294 12708
rect 18984 12696 19012 12736
rect 19150 12696 19156 12708
rect 18984 12668 19156 12696
rect 19150 12656 19156 12668
rect 19208 12656 19214 12708
rect 19306 12696 19334 12736
rect 21174 12724 21180 12776
rect 21232 12724 21238 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 21450 12764 21456 12776
rect 21407 12736 21456 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 20806 12696 20812 12708
rect 19306 12668 20812 12696
rect 20806 12656 20812 12668
rect 20864 12656 20870 12708
rect 22020 12696 22048 12795
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 22741 12835 22799 12841
rect 22741 12832 22753 12835
rect 22244 12804 22753 12832
rect 22244 12792 22250 12804
rect 22741 12801 22753 12804
rect 22787 12832 22799 12835
rect 23014 12832 23020 12844
rect 22787 12804 23020 12832
rect 22787 12801 22799 12804
rect 22741 12795 22799 12801
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 24872 12841 24900 12872
rect 25124 12869 25136 12903
rect 25170 12900 25182 12903
rect 25774 12900 25780 12912
rect 25170 12872 25780 12900
rect 25170 12869 25182 12872
rect 25124 12863 25182 12869
rect 25774 12860 25780 12872
rect 25832 12860 25838 12912
rect 25884 12900 25912 12940
rect 27341 12937 27353 12971
rect 27387 12968 27399 12971
rect 27798 12968 27804 12980
rect 27387 12940 27804 12968
rect 27387 12937 27399 12940
rect 27341 12931 27399 12937
rect 27798 12928 27804 12940
rect 27856 12928 27862 12980
rect 27908 12940 28764 12968
rect 27908 12900 27936 12940
rect 25884 12872 27936 12900
rect 28626 12860 28632 12912
rect 28684 12860 28690 12912
rect 28736 12900 28764 12940
rect 29730 12928 29736 12980
rect 29788 12968 29794 12980
rect 29917 12971 29975 12977
rect 29917 12968 29929 12971
rect 29788 12940 29929 12968
rect 29788 12928 29794 12940
rect 29917 12937 29929 12940
rect 29963 12937 29975 12971
rect 31205 12971 31263 12977
rect 31205 12968 31217 12971
rect 29917 12931 29975 12937
rect 30024 12940 31217 12968
rect 30024 12900 30052 12940
rect 31205 12937 31217 12940
rect 31251 12937 31263 12971
rect 31205 12931 31263 12937
rect 31478 12928 31484 12980
rect 31536 12968 31542 12980
rect 34790 12968 34796 12980
rect 31536 12940 34796 12968
rect 31536 12928 31542 12940
rect 34790 12928 34796 12940
rect 34848 12968 34854 12980
rect 35161 12971 35219 12977
rect 35161 12968 35173 12971
rect 34848 12940 35173 12968
rect 34848 12928 34854 12940
rect 35161 12937 35173 12940
rect 35207 12937 35219 12971
rect 35161 12931 35219 12937
rect 35250 12928 35256 12980
rect 35308 12968 35314 12980
rect 39666 12968 39672 12980
rect 35308 12940 39672 12968
rect 35308 12928 35314 12940
rect 39666 12928 39672 12940
rect 39724 12928 39730 12980
rect 41969 12971 42027 12977
rect 41969 12937 41981 12971
rect 42015 12968 42027 12971
rect 42794 12968 42800 12980
rect 42015 12940 42800 12968
rect 42015 12937 42027 12940
rect 41969 12931 42027 12937
rect 42794 12928 42800 12940
rect 42852 12928 42858 12980
rect 43165 12971 43223 12977
rect 43165 12937 43177 12971
rect 43211 12968 43223 12971
rect 43346 12968 43352 12980
rect 43211 12940 43352 12968
rect 43211 12937 43223 12940
rect 43165 12931 43223 12937
rect 43346 12928 43352 12940
rect 43404 12928 43410 12980
rect 32306 12900 32312 12912
rect 28736 12872 30052 12900
rect 30208 12872 32312 12900
rect 24857 12835 24915 12841
rect 24857 12801 24869 12835
rect 24903 12801 24915 12835
rect 26142 12832 26148 12844
rect 24857 12795 24915 12801
rect 24964 12804 26148 12832
rect 24762 12724 24768 12776
rect 24820 12764 24826 12776
rect 24964 12764 24992 12804
rect 26142 12792 26148 12804
rect 26200 12832 26206 12844
rect 26200 12804 26280 12832
rect 26200 12792 26206 12804
rect 24820 12736 24992 12764
rect 24820 12724 24826 12736
rect 26252 12705 26280 12804
rect 26878 12792 26884 12844
rect 26936 12832 26942 12844
rect 27249 12835 27307 12841
rect 27249 12832 27261 12835
rect 26936 12804 27261 12832
rect 26936 12792 26942 12804
rect 27249 12801 27261 12804
rect 27295 12801 27307 12835
rect 27249 12795 27307 12801
rect 27433 12835 27491 12841
rect 27433 12801 27445 12835
rect 27479 12832 27491 12835
rect 27798 12832 27804 12844
rect 27479 12804 27804 12832
rect 27479 12801 27491 12804
rect 27433 12795 27491 12801
rect 27798 12792 27804 12804
rect 27856 12792 27862 12844
rect 29730 12724 29736 12776
rect 29788 12764 29794 12776
rect 30208 12764 30236 12872
rect 32306 12860 32312 12872
rect 32364 12900 32370 12912
rect 34048 12903 34106 12909
rect 32364 12872 33824 12900
rect 32364 12860 32370 12872
rect 33796 12844 33824 12872
rect 34048 12869 34060 12903
rect 34094 12900 34106 12903
rect 34514 12900 34520 12912
rect 34094 12872 34520 12900
rect 34094 12869 34106 12872
rect 34048 12863 34106 12869
rect 34514 12860 34520 12872
rect 34572 12860 34578 12912
rect 36078 12860 36084 12912
rect 36136 12860 36142 12912
rect 36173 12903 36231 12909
rect 36173 12869 36185 12903
rect 36219 12900 36231 12903
rect 38010 12900 38016 12912
rect 36219 12872 38016 12900
rect 36219 12869 36231 12872
rect 36173 12863 36231 12869
rect 38010 12860 38016 12872
rect 38068 12860 38074 12912
rect 41892 12872 51074 12900
rect 30742 12792 30748 12844
rect 30800 12832 30806 12844
rect 31021 12835 31079 12841
rect 31021 12832 31033 12835
rect 30800 12804 31033 12832
rect 30800 12792 30806 12804
rect 31021 12801 31033 12804
rect 31067 12801 31079 12835
rect 31021 12795 31079 12801
rect 31297 12835 31355 12841
rect 31297 12801 31309 12835
rect 31343 12801 31355 12835
rect 31297 12795 31355 12801
rect 29788 12736 30236 12764
rect 29788 12724 29794 12736
rect 31110 12724 31116 12776
rect 31168 12764 31174 12776
rect 31312 12764 31340 12795
rect 32582 12792 32588 12844
rect 32640 12792 32646 12844
rect 32766 12792 32772 12844
rect 32824 12832 32830 12844
rect 32861 12835 32919 12841
rect 32861 12832 32873 12835
rect 32824 12804 32873 12832
rect 32824 12792 32830 12804
rect 32861 12801 32873 12804
rect 32907 12801 32919 12835
rect 32861 12795 32919 12801
rect 33778 12792 33784 12844
rect 33836 12792 33842 12844
rect 34790 12792 34796 12844
rect 34848 12832 34854 12844
rect 35897 12835 35955 12841
rect 35897 12832 35909 12835
rect 34848 12804 35909 12832
rect 34848 12792 34854 12804
rect 35897 12801 35909 12804
rect 35943 12801 35955 12835
rect 35897 12795 35955 12801
rect 36265 12835 36323 12841
rect 36265 12801 36277 12835
rect 36311 12832 36323 12835
rect 37274 12832 37280 12844
rect 36311 12804 37280 12832
rect 36311 12801 36323 12804
rect 36265 12795 36323 12801
rect 37274 12792 37280 12804
rect 37332 12792 37338 12844
rect 38654 12792 38660 12844
rect 38712 12832 38718 12844
rect 39666 12832 39672 12844
rect 38712 12804 39672 12832
rect 38712 12792 38718 12804
rect 39666 12792 39672 12804
rect 39724 12832 39730 12844
rect 41892 12841 41920 12872
rect 41877 12835 41935 12841
rect 41877 12832 41889 12835
rect 39724 12804 41889 12832
rect 39724 12792 39730 12804
rect 41877 12801 41889 12804
rect 41923 12801 41935 12835
rect 41877 12795 41935 12801
rect 42702 12792 42708 12844
rect 42760 12832 42766 12844
rect 42797 12835 42855 12841
rect 42797 12832 42809 12835
rect 42760 12804 42809 12832
rect 42760 12792 42766 12804
rect 42797 12801 42809 12804
rect 42843 12801 42855 12835
rect 42797 12795 42855 12801
rect 42978 12792 42984 12844
rect 43036 12792 43042 12844
rect 51046 12832 51074 12872
rect 56134 12832 56140 12844
rect 51046 12804 56140 12832
rect 56134 12792 56140 12804
rect 56192 12792 56198 12844
rect 31168 12736 31340 12764
rect 31168 12724 31174 12736
rect 32398 12724 32404 12776
rect 32456 12764 32462 12776
rect 33042 12764 33048 12776
rect 32456 12736 33048 12764
rect 32456 12724 32462 12736
rect 33042 12724 33048 12736
rect 33100 12724 33106 12776
rect 33226 12724 33232 12776
rect 33284 12724 33290 12776
rect 35986 12724 35992 12776
rect 36044 12764 36050 12776
rect 42150 12764 42156 12776
rect 36044 12736 42156 12764
rect 36044 12724 36050 12736
rect 42150 12724 42156 12736
rect 42208 12724 42214 12776
rect 26237 12699 26295 12705
rect 22020 12668 24900 12696
rect 11974 12588 11980 12640
rect 12032 12628 12038 12640
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 12032 12600 12633 12628
rect 12032 12588 12038 12600
rect 12621 12597 12633 12600
rect 12667 12597 12679 12631
rect 12621 12591 12679 12597
rect 16209 12631 16267 12637
rect 16209 12597 16221 12631
rect 16255 12628 16267 12631
rect 17218 12628 17224 12640
rect 16255 12600 17224 12628
rect 16255 12597 16267 12600
rect 16209 12591 16267 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 18325 12631 18383 12637
rect 18325 12597 18337 12631
rect 18371 12628 18383 12631
rect 18414 12628 18420 12640
rect 18371 12600 18420 12628
rect 18371 12597 18383 12600
rect 18325 12591 18383 12597
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 18506 12588 18512 12640
rect 18564 12628 18570 12640
rect 22189 12631 22247 12637
rect 22189 12628 22201 12631
rect 18564 12600 22201 12628
rect 18564 12588 18570 12600
rect 22189 12597 22201 12600
rect 22235 12597 22247 12631
rect 24872 12628 24900 12668
rect 26237 12665 26249 12699
rect 26283 12665 26295 12699
rect 26237 12659 26295 12665
rect 27982 12656 27988 12708
rect 28040 12696 28046 12708
rect 32490 12696 32496 12708
rect 28040 12668 32496 12696
rect 28040 12656 28046 12668
rect 32490 12656 32496 12668
rect 32548 12656 32554 12708
rect 32677 12699 32735 12705
rect 32677 12665 32689 12699
rect 32723 12696 32735 12699
rect 32723 12668 33824 12696
rect 32723 12665 32735 12668
rect 32677 12659 32735 12665
rect 26418 12628 26424 12640
rect 24872 12600 26424 12628
rect 22189 12591 22247 12597
rect 26418 12588 26424 12600
rect 26476 12588 26482 12640
rect 30837 12631 30895 12637
rect 30837 12597 30849 12631
rect 30883 12628 30895 12631
rect 31018 12628 31024 12640
rect 30883 12600 31024 12628
rect 30883 12597 30895 12600
rect 30837 12591 30895 12597
rect 31018 12588 31024 12600
rect 31076 12588 31082 12640
rect 33796 12628 33824 12668
rect 36446 12656 36452 12708
rect 36504 12656 36510 12708
rect 40862 12656 40868 12708
rect 40920 12696 40926 12708
rect 41138 12696 41144 12708
rect 40920 12668 41144 12696
rect 40920 12656 40926 12668
rect 41138 12656 41144 12668
rect 41196 12696 41202 12708
rect 41414 12696 41420 12708
rect 41196 12668 41420 12696
rect 41196 12656 41202 12668
rect 41414 12656 41420 12668
rect 41472 12656 41478 12708
rect 41966 12656 41972 12708
rect 42024 12696 42030 12708
rect 42024 12668 43116 12696
rect 42024 12656 42030 12668
rect 43088 12640 43116 12668
rect 35894 12628 35900 12640
rect 33796 12600 35900 12628
rect 35894 12588 35900 12600
rect 35952 12588 35958 12640
rect 36170 12588 36176 12640
rect 36228 12628 36234 12640
rect 42794 12628 42800 12640
rect 36228 12600 42800 12628
rect 36228 12588 36234 12600
rect 42794 12588 42800 12600
rect 42852 12588 42858 12640
rect 43070 12588 43076 12640
rect 43128 12588 43134 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 10502 12384 10508 12436
rect 10560 12424 10566 12436
rect 10597 12427 10655 12433
rect 10597 12424 10609 12427
rect 10560 12396 10609 12424
rect 10560 12384 10566 12396
rect 10597 12393 10609 12396
rect 10643 12393 10655 12427
rect 10597 12387 10655 12393
rect 11606 12384 11612 12436
rect 11664 12384 11670 12436
rect 14182 12424 14188 12436
rect 12406 12396 14188 12424
rect 2314 12316 2320 12368
rect 2372 12316 2378 12368
rect 6178 12316 6184 12368
rect 6236 12356 6242 12368
rect 12406 12356 12434 12396
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 14826 12384 14832 12436
rect 14884 12424 14890 12436
rect 16025 12427 16083 12433
rect 16025 12424 16037 12427
rect 14884 12396 16037 12424
rect 14884 12384 14890 12396
rect 16025 12393 16037 12396
rect 16071 12393 16083 12427
rect 16025 12387 16083 12393
rect 16114 12384 16120 12436
rect 16172 12424 16178 12436
rect 17129 12427 17187 12433
rect 17129 12424 17141 12427
rect 16172 12396 17141 12424
rect 16172 12384 16178 12396
rect 17129 12393 17141 12396
rect 17175 12393 17187 12427
rect 17129 12387 17187 12393
rect 18046 12384 18052 12436
rect 18104 12424 18110 12436
rect 18601 12427 18659 12433
rect 18601 12424 18613 12427
rect 18104 12396 18613 12424
rect 18104 12384 18110 12396
rect 18601 12393 18613 12396
rect 18647 12393 18659 12427
rect 18601 12387 18659 12393
rect 19242 12384 19248 12436
rect 19300 12424 19306 12436
rect 21818 12424 21824 12436
rect 19300 12396 21824 12424
rect 19300 12384 19306 12396
rect 21818 12384 21824 12396
rect 21876 12384 21882 12436
rect 22186 12384 22192 12436
rect 22244 12384 22250 12436
rect 27062 12424 27068 12436
rect 25700 12396 27068 12424
rect 20254 12356 20260 12368
rect 6236 12328 12434 12356
rect 13556 12328 20260 12356
rect 6236 12316 6242 12328
rect 9950 12288 9956 12300
rect 2148 12260 9956 12288
rect 2148 12229 2176 12260
rect 9950 12248 9956 12260
rect 10008 12288 10014 12300
rect 10008 12260 12434 12288
rect 10008 12248 10014 12260
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 2590 12180 2596 12232
rect 2648 12180 2654 12232
rect 10505 12223 10563 12229
rect 10505 12189 10517 12223
rect 10551 12220 10563 12223
rect 10594 12220 10600 12232
rect 10551 12192 10600 12220
rect 10551 12189 10563 12192
rect 10505 12183 10563 12189
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 10686 12180 10692 12232
rect 10744 12180 10750 12232
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12220 11483 12223
rect 11974 12220 11980 12232
rect 11471 12192 11980 12220
rect 11471 12189 11483 12192
rect 11425 12183 11483 12189
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 12406 12152 12434 12260
rect 13556 12229 13584 12328
rect 20254 12316 20260 12328
rect 20312 12316 20318 12368
rect 24854 12316 24860 12368
rect 24912 12356 24918 12368
rect 25133 12359 25191 12365
rect 25133 12356 25145 12359
rect 24912 12328 25145 12356
rect 24912 12316 24918 12328
rect 25133 12325 25145 12328
rect 25179 12325 25191 12359
rect 25133 12319 25191 12325
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 14369 12291 14427 12297
rect 14369 12288 14381 12291
rect 13679 12260 14381 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 14369 12257 14381 12260
rect 14415 12257 14427 12291
rect 14369 12251 14427 12257
rect 15010 12248 15016 12300
rect 15068 12288 15074 12300
rect 17954 12288 17960 12300
rect 15068 12260 17960 12288
rect 15068 12248 15074 12260
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 18506 12288 18512 12300
rect 18064 12260 18512 12288
rect 13541 12223 13599 12229
rect 13541 12189 13553 12223
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12220 14519 12223
rect 15746 12220 15752 12232
rect 14507 12192 15752 12220
rect 14507 12189 14519 12192
rect 14461 12183 14519 12189
rect 13170 12152 13176 12164
rect 12406 12124 13176 12152
rect 13170 12112 13176 12124
rect 13228 12112 13234 12164
rect 13354 12112 13360 12164
rect 13412 12152 13418 12164
rect 13740 12152 13768 12183
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15838 12180 15844 12232
rect 15896 12180 15902 12232
rect 16942 12180 16948 12232
rect 17000 12180 17006 12232
rect 17678 12180 17684 12232
rect 17736 12220 17742 12232
rect 18064 12220 18092 12260
rect 18506 12248 18512 12260
rect 18564 12248 18570 12300
rect 20070 12248 20076 12300
rect 20128 12288 20134 12300
rect 20530 12288 20536 12300
rect 20128 12260 20536 12288
rect 20128 12248 20134 12260
rect 20530 12248 20536 12260
rect 20588 12248 20594 12300
rect 25700 12297 25728 12396
rect 27062 12384 27068 12396
rect 27120 12384 27126 12436
rect 27614 12384 27620 12436
rect 27672 12384 27678 12436
rect 30006 12384 30012 12436
rect 30064 12384 30070 12436
rect 30116 12396 31984 12424
rect 26510 12316 26516 12368
rect 26568 12356 26574 12368
rect 29914 12356 29920 12368
rect 26568 12328 29920 12356
rect 26568 12316 26574 12328
rect 29914 12316 29920 12328
rect 29972 12316 29978 12368
rect 25685 12291 25743 12297
rect 25685 12257 25697 12291
rect 25731 12257 25743 12291
rect 25685 12251 25743 12257
rect 26234 12248 26240 12300
rect 26292 12288 26298 12300
rect 26605 12291 26663 12297
rect 26605 12288 26617 12291
rect 26292 12260 26617 12288
rect 26292 12248 26298 12260
rect 26605 12257 26617 12260
rect 26651 12257 26663 12291
rect 26605 12251 26663 12257
rect 29086 12248 29092 12300
rect 29144 12288 29150 12300
rect 30116 12288 30144 12396
rect 31018 12316 31024 12368
rect 31076 12316 31082 12368
rect 31110 12316 31116 12368
rect 31168 12356 31174 12368
rect 31570 12356 31576 12368
rect 31168 12328 31576 12356
rect 31168 12316 31174 12328
rect 31570 12316 31576 12328
rect 31628 12316 31634 12368
rect 29144 12260 30144 12288
rect 30300 12260 31800 12288
rect 29144 12248 29150 12260
rect 17736 12192 18092 12220
rect 17736 12180 17742 12192
rect 18414 12180 18420 12232
rect 18472 12180 18478 12232
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 20622 12220 20628 12232
rect 20312 12192 20628 12220
rect 20312 12180 20318 12192
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 20809 12223 20867 12229
rect 20809 12189 20821 12223
rect 20855 12220 20867 12223
rect 20898 12220 20904 12232
rect 20855 12192 20904 12220
rect 20855 12189 20867 12192
rect 20809 12183 20867 12189
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 21082 12229 21088 12232
rect 21076 12183 21088 12229
rect 21082 12180 21088 12183
rect 21140 12180 21146 12232
rect 24670 12180 24676 12232
rect 24728 12220 24734 12232
rect 24857 12223 24915 12229
rect 24857 12220 24869 12223
rect 24728 12192 24869 12220
rect 24728 12180 24734 12192
rect 24857 12189 24869 12192
rect 24903 12189 24915 12223
rect 24857 12183 24915 12189
rect 25133 12223 25191 12229
rect 25133 12189 25145 12223
rect 25179 12220 25191 12223
rect 25869 12223 25927 12229
rect 25179 12192 25268 12220
rect 25179 12189 25191 12192
rect 25133 12183 25191 12189
rect 13412 12124 14964 12152
rect 13412 12112 13418 12124
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 14829 12087 14887 12093
rect 14829 12084 14841 12087
rect 14516 12056 14841 12084
rect 14516 12044 14522 12056
rect 14829 12053 14841 12056
rect 14875 12053 14887 12087
rect 14936 12084 14964 12124
rect 15194 12112 15200 12164
rect 15252 12152 15258 12164
rect 24762 12152 24768 12164
rect 15252 12124 24768 12152
rect 15252 12112 15258 12124
rect 24762 12112 24768 12124
rect 24820 12112 24826 12164
rect 25240 12096 25268 12192
rect 25869 12189 25881 12223
rect 25915 12189 25927 12223
rect 25869 12183 25927 12189
rect 25314 12112 25320 12164
rect 25372 12152 25378 12164
rect 25884 12152 25912 12183
rect 25958 12180 25964 12232
rect 26016 12220 26022 12232
rect 26513 12223 26571 12229
rect 26513 12220 26525 12223
rect 26016 12192 26525 12220
rect 26016 12180 26022 12192
rect 26513 12189 26525 12192
rect 26559 12189 26571 12223
rect 26513 12183 26571 12189
rect 27617 12223 27675 12229
rect 27617 12189 27629 12223
rect 27663 12189 27675 12223
rect 27617 12183 27675 12189
rect 25372 12124 25912 12152
rect 25976 12124 26648 12152
rect 25372 12112 25378 12124
rect 17865 12087 17923 12093
rect 17865 12084 17877 12087
rect 14936 12056 17877 12084
rect 14829 12047 14887 12053
rect 17865 12053 17877 12056
rect 17911 12053 17923 12087
rect 17865 12047 17923 12053
rect 17954 12044 17960 12096
rect 18012 12084 18018 12096
rect 25130 12084 25136 12096
rect 18012 12056 25136 12084
rect 18012 12044 18018 12056
rect 25130 12044 25136 12056
rect 25188 12044 25194 12096
rect 25222 12044 25228 12096
rect 25280 12084 25286 12096
rect 25976 12084 26004 12124
rect 25280 12056 26004 12084
rect 25280 12044 25286 12056
rect 26050 12044 26056 12096
rect 26108 12044 26114 12096
rect 26510 12044 26516 12096
rect 26568 12044 26574 12096
rect 26620 12084 26648 12124
rect 26694 12112 26700 12164
rect 26752 12152 26758 12164
rect 26789 12155 26847 12161
rect 26789 12152 26801 12155
rect 26752 12124 26801 12152
rect 26752 12112 26758 12124
rect 26789 12121 26801 12124
rect 26835 12121 26847 12155
rect 27632 12152 27660 12183
rect 27798 12180 27804 12232
rect 27856 12220 27862 12232
rect 28258 12220 28264 12232
rect 27856 12192 28264 12220
rect 27856 12180 27862 12192
rect 28258 12180 28264 12192
rect 28316 12180 28322 12232
rect 30098 12180 30104 12232
rect 30156 12220 30162 12232
rect 30193 12223 30251 12229
rect 30193 12220 30205 12223
rect 30156 12192 30205 12220
rect 30156 12180 30162 12192
rect 30193 12189 30205 12192
rect 30239 12189 30251 12223
rect 30193 12183 30251 12189
rect 28442 12152 28448 12164
rect 27632 12124 28448 12152
rect 26789 12115 26847 12121
rect 28442 12112 28448 12124
rect 28500 12152 28506 12164
rect 30300 12152 30328 12260
rect 30469 12223 30527 12229
rect 30469 12189 30481 12223
rect 30515 12220 30527 12223
rect 31110 12220 31116 12232
rect 30515 12192 31116 12220
rect 30515 12189 30527 12192
rect 30469 12183 30527 12189
rect 31110 12180 31116 12192
rect 31168 12180 31174 12232
rect 31202 12180 31208 12232
rect 31260 12180 31266 12232
rect 31297 12223 31355 12229
rect 31297 12189 31309 12223
rect 31343 12220 31355 12223
rect 31386 12220 31392 12232
rect 31343 12192 31392 12220
rect 31343 12189 31355 12192
rect 31297 12183 31355 12189
rect 31386 12180 31392 12192
rect 31444 12180 31450 12232
rect 31772 12229 31800 12260
rect 31956 12229 31984 12396
rect 35802 12384 35808 12436
rect 35860 12384 35866 12436
rect 37829 12427 37887 12433
rect 36280 12396 37412 12424
rect 32766 12316 32772 12368
rect 32824 12356 32830 12368
rect 36280 12356 36308 12396
rect 32824 12328 36308 12356
rect 32824 12316 32830 12328
rect 33778 12248 33784 12300
rect 33836 12288 33842 12300
rect 36265 12291 36323 12297
rect 36265 12288 36277 12291
rect 33836 12260 36277 12288
rect 33836 12248 33842 12260
rect 36265 12257 36277 12260
rect 36311 12257 36323 12291
rect 36265 12251 36323 12257
rect 36541 12291 36599 12297
rect 36541 12257 36553 12291
rect 36587 12288 36599 12291
rect 36630 12288 36636 12300
rect 36587 12260 36636 12288
rect 36587 12257 36599 12260
rect 36541 12251 36599 12257
rect 36630 12248 36636 12260
rect 36688 12248 36694 12300
rect 31757 12223 31815 12229
rect 31757 12189 31769 12223
rect 31803 12189 31815 12223
rect 31757 12183 31815 12189
rect 31941 12223 31999 12229
rect 31941 12189 31953 12223
rect 31987 12189 31999 12223
rect 31941 12183 31999 12189
rect 35253 12223 35311 12229
rect 35253 12189 35265 12223
rect 35299 12220 35311 12223
rect 35342 12220 35348 12232
rect 35299 12192 35348 12220
rect 35299 12189 35311 12192
rect 35253 12183 35311 12189
rect 35342 12180 35348 12192
rect 35400 12180 35406 12232
rect 35526 12180 35532 12232
rect 35584 12180 35590 12232
rect 35621 12223 35679 12229
rect 35621 12189 35633 12223
rect 35667 12220 35679 12223
rect 35667 12192 36400 12220
rect 35667 12189 35679 12192
rect 35621 12183 35679 12189
rect 28500 12124 30328 12152
rect 31021 12155 31079 12161
rect 28500 12112 28506 12124
rect 31021 12121 31033 12155
rect 31067 12152 31079 12155
rect 31067 12124 31340 12152
rect 31067 12121 31079 12124
rect 31021 12115 31079 12121
rect 31312 12096 31340 12124
rect 31570 12112 31576 12164
rect 31628 12152 31634 12164
rect 31849 12155 31907 12161
rect 31849 12152 31861 12155
rect 31628 12124 31861 12152
rect 31628 12112 31634 12124
rect 31849 12121 31861 12124
rect 31895 12121 31907 12155
rect 31849 12115 31907 12121
rect 34330 12112 34336 12164
rect 34388 12152 34394 12164
rect 35437 12155 35495 12161
rect 35437 12152 35449 12155
rect 34388 12124 35449 12152
rect 34388 12112 34394 12124
rect 35437 12121 35449 12124
rect 35483 12121 35495 12155
rect 35437 12115 35495 12121
rect 26878 12084 26884 12096
rect 26620 12056 26884 12084
rect 26878 12044 26884 12056
rect 26936 12044 26942 12096
rect 30282 12044 30288 12096
rect 30340 12084 30346 12096
rect 30377 12087 30435 12093
rect 30377 12084 30389 12087
rect 30340 12056 30389 12084
rect 30340 12044 30346 12056
rect 30377 12053 30389 12056
rect 30423 12053 30435 12087
rect 30377 12047 30435 12053
rect 31294 12044 31300 12096
rect 31352 12044 31358 12096
rect 32858 12044 32864 12096
rect 32916 12084 32922 12096
rect 35728 12084 35756 12192
rect 32916 12056 35756 12084
rect 36372 12084 36400 12192
rect 37384 12152 37412 12396
rect 37829 12393 37841 12427
rect 37875 12424 37887 12427
rect 38010 12424 38016 12436
rect 37875 12396 38016 12424
rect 37875 12393 37887 12396
rect 37829 12387 37887 12393
rect 38010 12384 38016 12396
rect 38068 12384 38074 12436
rect 38378 12384 38384 12436
rect 38436 12424 38442 12436
rect 38436 12396 46244 12424
rect 38436 12384 38442 12396
rect 41598 12356 41604 12368
rect 40328 12328 41604 12356
rect 40034 12180 40040 12232
rect 40092 12180 40098 12232
rect 40185 12223 40243 12229
rect 40185 12189 40197 12223
rect 40231 12220 40243 12223
rect 40328 12220 40356 12328
rect 41598 12316 41604 12328
rect 41656 12316 41662 12368
rect 41690 12316 41696 12368
rect 41748 12316 41754 12368
rect 46216 12356 46244 12396
rect 46290 12384 46296 12436
rect 46348 12424 46354 12436
rect 53190 12424 53196 12436
rect 46348 12396 53196 12424
rect 46348 12384 46354 12396
rect 53190 12384 53196 12396
rect 53248 12424 53254 12436
rect 54386 12424 54392 12436
rect 53248 12396 54392 12424
rect 53248 12384 53254 12396
rect 54386 12384 54392 12396
rect 54444 12384 54450 12436
rect 53466 12356 53472 12368
rect 46216 12328 53472 12356
rect 53466 12316 53472 12328
rect 53524 12316 53530 12368
rect 41708 12288 41736 12316
rect 40558 12260 41736 12288
rect 40231 12192 40356 12220
rect 40231 12189 40243 12192
rect 40185 12183 40243 12189
rect 40402 12180 40408 12232
rect 40460 12180 40466 12232
rect 40558 12229 40586 12260
rect 40543 12223 40601 12229
rect 40543 12189 40555 12223
rect 40589 12189 40601 12223
rect 40543 12183 40601 12189
rect 41138 12180 41144 12232
rect 41196 12180 41202 12232
rect 41322 12229 41328 12232
rect 41279 12223 41328 12229
rect 41279 12189 41291 12223
rect 41325 12189 41328 12223
rect 41279 12183 41328 12189
rect 41322 12180 41328 12183
rect 41380 12180 41386 12232
rect 41414 12180 41420 12232
rect 41472 12180 41478 12232
rect 41506 12180 41512 12232
rect 41564 12180 41570 12232
rect 41621 12229 41649 12260
rect 43438 12248 43444 12300
rect 43496 12288 43502 12300
rect 53558 12288 53564 12300
rect 43496 12260 53564 12288
rect 43496 12248 43502 12260
rect 53558 12248 53564 12260
rect 53616 12248 53622 12300
rect 41621 12223 41683 12229
rect 41621 12192 41637 12223
rect 41625 12189 41637 12192
rect 41671 12189 41683 12223
rect 41625 12183 41683 12189
rect 57882 12180 57888 12232
rect 57940 12180 57946 12232
rect 40313 12155 40371 12161
rect 40313 12152 40325 12155
rect 37384 12124 40325 12152
rect 40313 12121 40325 12124
rect 40359 12152 40371 12155
rect 40862 12152 40868 12164
rect 40359 12124 40868 12152
rect 40359 12121 40371 12124
rect 40313 12115 40371 12121
rect 40862 12112 40868 12124
rect 40920 12112 40926 12164
rect 58158 12112 58164 12164
rect 58216 12112 58222 12164
rect 37918 12084 37924 12096
rect 36372 12056 37924 12084
rect 32916 12044 32922 12056
rect 37918 12044 37924 12056
rect 37976 12084 37982 12096
rect 38378 12084 38384 12096
rect 37976 12056 38384 12084
rect 37976 12044 37982 12056
rect 38378 12044 38384 12056
rect 38436 12044 38442 12096
rect 40681 12087 40739 12093
rect 40681 12053 40693 12087
rect 40727 12084 40739 12087
rect 41138 12084 41144 12096
rect 40727 12056 41144 12084
rect 40727 12053 40739 12056
rect 40681 12047 40739 12053
rect 41138 12044 41144 12056
rect 41196 12044 41202 12096
rect 41782 12044 41788 12096
rect 41840 12044 41846 12096
rect 46382 12044 46388 12096
rect 46440 12084 46446 12096
rect 46842 12084 46848 12096
rect 46440 12056 46848 12084
rect 46440 12044 46446 12056
rect 46842 12044 46848 12056
rect 46900 12044 46906 12096
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 2590 11840 2596 11892
rect 2648 11880 2654 11892
rect 11054 11880 11060 11892
rect 2648 11852 11060 11880
rect 2648 11840 2654 11852
rect 11054 11840 11060 11852
rect 11112 11840 11118 11892
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 13872 11852 14657 11880
rect 13872 11840 13878 11852
rect 14645 11849 14657 11852
rect 14691 11849 14703 11883
rect 14645 11843 14703 11849
rect 14918 11840 14924 11892
rect 14976 11880 14982 11892
rect 14976 11852 15516 11880
rect 14976 11840 14982 11852
rect 934 11772 940 11824
rect 992 11812 998 11824
rect 1857 11815 1915 11821
rect 1857 11812 1869 11815
rect 992 11784 1869 11812
rect 992 11772 998 11784
rect 1857 11781 1869 11784
rect 1903 11781 1915 11815
rect 1857 11775 1915 11781
rect 10686 11772 10692 11824
rect 10744 11812 10750 11824
rect 15488 11821 15516 11852
rect 17402 11840 17408 11892
rect 17460 11840 17466 11892
rect 18141 11883 18199 11889
rect 18141 11849 18153 11883
rect 18187 11849 18199 11883
rect 24026 11880 24032 11892
rect 18141 11843 18199 11849
rect 18248 11852 24032 11880
rect 15473 11815 15531 11821
rect 10744 11784 15332 11812
rect 10744 11772 10750 11784
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11744 1639 11747
rect 11977 11747 12035 11753
rect 1627 11716 2774 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 2746 11676 2774 11716
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 14366 11744 14372 11756
rect 12023 11716 14372 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 14458 11704 14464 11756
rect 14516 11704 14522 11756
rect 15304 11744 15332 11784
rect 15473 11781 15485 11815
rect 15519 11781 15531 11815
rect 15473 11775 15531 11781
rect 15562 11772 15568 11824
rect 15620 11812 15626 11824
rect 15673 11815 15731 11821
rect 15673 11812 15685 11815
rect 15620 11784 15685 11812
rect 15620 11772 15626 11784
rect 15673 11781 15685 11784
rect 15719 11781 15731 11815
rect 18156 11812 18184 11843
rect 15673 11775 15731 11781
rect 15764 11784 18184 11812
rect 15764 11744 15792 11784
rect 15304 11716 15792 11744
rect 17218 11704 17224 11756
rect 17276 11704 17282 11756
rect 17957 11747 18015 11753
rect 17957 11713 17969 11747
rect 18003 11744 18015 11747
rect 18248 11744 18276 11852
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 24486 11840 24492 11892
rect 24544 11880 24550 11892
rect 24581 11883 24639 11889
rect 24581 11880 24593 11883
rect 24544 11852 24593 11880
rect 24544 11840 24550 11852
rect 24581 11849 24593 11852
rect 24627 11849 24639 11883
rect 24581 11843 24639 11849
rect 24673 11883 24731 11889
rect 24673 11849 24685 11883
rect 24719 11880 24731 11883
rect 24762 11880 24768 11892
rect 24719 11852 24768 11880
rect 24719 11849 24731 11852
rect 24673 11843 24731 11849
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 25314 11840 25320 11892
rect 25372 11840 25378 11892
rect 25406 11840 25412 11892
rect 25464 11880 25470 11892
rect 25682 11880 25688 11892
rect 25464 11852 25688 11880
rect 25464 11840 25470 11852
rect 25682 11840 25688 11852
rect 25740 11840 25746 11892
rect 25777 11883 25835 11889
rect 25777 11849 25789 11883
rect 25823 11880 25835 11883
rect 26142 11880 26148 11892
rect 25823 11852 26148 11880
rect 25823 11849 25835 11852
rect 25777 11843 25835 11849
rect 26142 11840 26148 11852
rect 26200 11840 26206 11892
rect 26510 11840 26516 11892
rect 26568 11880 26574 11892
rect 29822 11880 29828 11892
rect 26568 11852 29828 11880
rect 26568 11840 26574 11852
rect 29822 11840 29828 11852
rect 29880 11840 29886 11892
rect 31110 11840 31116 11892
rect 31168 11880 31174 11892
rect 31389 11883 31447 11889
rect 31389 11880 31401 11883
rect 31168 11852 31401 11880
rect 31168 11840 31174 11852
rect 31389 11849 31401 11852
rect 31435 11880 31447 11883
rect 31846 11880 31852 11892
rect 31435 11852 31852 11880
rect 31435 11849 31447 11852
rect 31389 11843 31447 11849
rect 31846 11840 31852 11852
rect 31904 11840 31910 11892
rect 31938 11840 31944 11892
rect 31996 11880 32002 11892
rect 32306 11880 32312 11892
rect 31996 11852 32312 11880
rect 31996 11840 32002 11852
rect 32306 11840 32312 11852
rect 32364 11840 32370 11892
rect 33413 11883 33471 11889
rect 33413 11849 33425 11883
rect 33459 11849 33471 11883
rect 33413 11843 33471 11849
rect 18322 11772 18328 11824
rect 18380 11812 18386 11824
rect 21082 11812 21088 11824
rect 18380 11784 21088 11812
rect 18380 11772 18386 11784
rect 21082 11772 21088 11784
rect 21140 11772 21146 11824
rect 21358 11772 21364 11824
rect 21416 11812 21422 11824
rect 24857 11815 24915 11821
rect 24857 11812 24869 11815
rect 21416 11784 24869 11812
rect 21416 11772 21422 11784
rect 24857 11781 24869 11784
rect 24903 11781 24915 11815
rect 24857 11775 24915 11781
rect 26050 11772 26056 11824
rect 26108 11812 26114 11824
rect 27402 11815 27460 11821
rect 27402 11812 27414 11815
rect 26108 11784 27414 11812
rect 26108 11772 26114 11784
rect 27402 11781 27414 11784
rect 27448 11781 27460 11815
rect 27402 11775 27460 11781
rect 27522 11772 27528 11824
rect 27580 11812 27586 11824
rect 31570 11812 31576 11824
rect 27580 11784 29960 11812
rect 27580 11772 27586 11784
rect 18003 11716 18276 11744
rect 18003 11713 18015 11716
rect 17957 11707 18015 11713
rect 11701 11679 11759 11685
rect 11701 11676 11713 11679
rect 2746 11648 11713 11676
rect 11701 11645 11713 11648
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 11885 11679 11943 11685
rect 11885 11645 11897 11679
rect 11931 11645 11943 11679
rect 11885 11639 11943 11645
rect 11146 11568 11152 11620
rect 11204 11608 11210 11620
rect 11900 11608 11928 11639
rect 12066 11636 12072 11688
rect 12124 11636 12130 11688
rect 12158 11636 12164 11688
rect 12216 11636 12222 11688
rect 12250 11636 12256 11688
rect 12308 11676 12314 11688
rect 17972 11676 18000 11707
rect 20346 11704 20352 11756
rect 20404 11704 20410 11756
rect 24489 11747 24547 11753
rect 20548 11716 22094 11744
rect 12308 11648 18000 11676
rect 12308 11636 12314 11648
rect 19610 11636 19616 11688
rect 19668 11676 19674 11688
rect 20070 11676 20076 11688
rect 19668 11648 20076 11676
rect 19668 11636 19674 11648
rect 20070 11636 20076 11648
rect 20128 11636 20134 11688
rect 20254 11636 20260 11688
rect 20312 11676 20318 11688
rect 20441 11679 20499 11685
rect 20441 11676 20453 11679
rect 20312 11648 20453 11676
rect 20312 11636 20318 11648
rect 20441 11645 20453 11648
rect 20487 11645 20499 11679
rect 20441 11639 20499 11645
rect 20548 11608 20576 11716
rect 20625 11679 20683 11685
rect 20625 11645 20637 11679
rect 20671 11676 20683 11679
rect 20898 11676 20904 11688
rect 20671 11648 20904 11676
rect 20671 11645 20683 11648
rect 20625 11639 20683 11645
rect 20898 11636 20904 11648
rect 20956 11636 20962 11688
rect 22066 11676 22094 11716
rect 24489 11713 24501 11747
rect 24535 11744 24547 11747
rect 25222 11744 25228 11756
rect 24535 11716 25228 11744
rect 24535 11713 24547 11716
rect 24489 11707 24547 11713
rect 25222 11704 25228 11716
rect 25280 11704 25286 11756
rect 25682 11704 25688 11756
rect 25740 11704 25746 11756
rect 26786 11704 26792 11756
rect 26844 11744 26850 11756
rect 26844 11716 29224 11744
rect 26844 11704 26850 11716
rect 24946 11676 24952 11688
rect 22066 11648 24952 11676
rect 24946 11636 24952 11648
rect 25004 11636 25010 11688
rect 25961 11679 26019 11685
rect 25961 11645 25973 11679
rect 26007 11676 26019 11679
rect 26050 11676 26056 11688
rect 26007 11648 26056 11676
rect 26007 11645 26019 11648
rect 25961 11639 26019 11645
rect 26050 11636 26056 11648
rect 26108 11636 26114 11688
rect 27157 11679 27215 11685
rect 27157 11645 27169 11679
rect 27203 11645 27215 11679
rect 29196 11676 29224 11716
rect 29270 11704 29276 11756
rect 29328 11744 29334 11756
rect 29546 11744 29552 11756
rect 29328 11716 29552 11744
rect 29328 11704 29334 11716
rect 29546 11704 29552 11716
rect 29604 11704 29610 11756
rect 29638 11704 29644 11756
rect 29696 11704 29702 11756
rect 29822 11704 29828 11756
rect 29880 11704 29886 11756
rect 29932 11753 29960 11784
rect 30668 11784 31576 11812
rect 30668 11753 30696 11784
rect 31570 11772 31576 11784
rect 31628 11772 31634 11824
rect 31662 11772 31668 11824
rect 31720 11812 31726 11824
rect 33428 11812 33456 11843
rect 35342 11840 35348 11892
rect 35400 11880 35406 11892
rect 35618 11880 35624 11892
rect 35400 11852 35624 11880
rect 35400 11840 35406 11852
rect 35618 11840 35624 11852
rect 35676 11840 35682 11892
rect 42242 11840 42248 11892
rect 42300 11880 42306 11892
rect 56410 11880 56416 11892
rect 42300 11852 56416 11880
rect 42300 11840 42306 11852
rect 56410 11840 56416 11852
rect 56468 11840 56474 11892
rect 31720 11784 33456 11812
rect 31720 11772 31726 11784
rect 33594 11772 33600 11824
rect 33652 11812 33658 11824
rect 41046 11812 41052 11824
rect 33652 11784 41052 11812
rect 33652 11772 33658 11784
rect 41046 11772 41052 11784
rect 41104 11772 41110 11824
rect 41966 11772 41972 11824
rect 42024 11812 42030 11824
rect 46661 11815 46719 11821
rect 42024 11784 46612 11812
rect 42024 11772 42030 11784
rect 29917 11747 29975 11753
rect 29917 11713 29929 11747
rect 29963 11713 29975 11747
rect 29917 11707 29975 11713
rect 30653 11747 30711 11753
rect 30653 11713 30665 11747
rect 30699 11713 30711 11747
rect 30653 11707 30711 11713
rect 30742 11704 30748 11756
rect 30800 11744 30806 11756
rect 31297 11747 31355 11753
rect 31297 11744 31309 11747
rect 30800 11716 31309 11744
rect 30800 11704 30806 11716
rect 31297 11713 31309 11716
rect 31343 11713 31355 11747
rect 31297 11707 31355 11713
rect 31481 11747 31539 11753
rect 31481 11713 31493 11747
rect 31527 11744 31539 11747
rect 32858 11744 32864 11756
rect 31527 11716 32864 11744
rect 31527 11713 31539 11716
rect 31481 11707 31539 11713
rect 31496 11676 31524 11707
rect 32858 11704 32864 11716
rect 32916 11704 32922 11756
rect 32950 11704 32956 11756
rect 33008 11704 33014 11756
rect 33134 11704 33140 11756
rect 33192 11744 33198 11756
rect 33229 11747 33287 11753
rect 33229 11744 33241 11747
rect 33192 11716 33241 11744
rect 33192 11704 33198 11716
rect 33229 11713 33241 11716
rect 33275 11713 33287 11747
rect 33229 11707 33287 11713
rect 33778 11704 33784 11756
rect 33836 11744 33842 11756
rect 34609 11747 34667 11753
rect 34609 11744 34621 11747
rect 33836 11716 34621 11744
rect 33836 11704 33842 11716
rect 34609 11713 34621 11716
rect 34655 11713 34667 11747
rect 34609 11707 34667 11713
rect 34876 11747 34934 11753
rect 34876 11713 34888 11747
rect 34922 11744 34934 11747
rect 35342 11744 35348 11756
rect 34922 11716 35348 11744
rect 34922 11713 34934 11716
rect 34876 11707 34934 11713
rect 35342 11704 35348 11716
rect 35400 11704 35406 11756
rect 38746 11704 38752 11756
rect 38804 11704 38810 11756
rect 41138 11704 41144 11756
rect 41196 11744 41202 11756
rect 42242 11744 42248 11756
rect 41196 11716 42248 11744
rect 41196 11704 41202 11716
rect 42242 11704 42248 11716
rect 42300 11704 42306 11756
rect 42334 11704 42340 11756
rect 42392 11744 42398 11756
rect 46290 11744 46296 11756
rect 42392 11716 46296 11744
rect 42392 11704 42398 11716
rect 46290 11704 46296 11716
rect 46348 11704 46354 11756
rect 46584 11744 46612 11784
rect 46661 11781 46673 11815
rect 46707 11812 46719 11815
rect 59446 11812 59452 11824
rect 46707 11784 59452 11812
rect 46707 11781 46719 11784
rect 46661 11775 46719 11781
rect 59446 11772 59452 11784
rect 59504 11772 59510 11824
rect 48314 11744 48320 11756
rect 46584 11716 48320 11744
rect 48314 11704 48320 11716
rect 48372 11704 48378 11756
rect 57149 11747 57207 11753
rect 57149 11713 57161 11747
rect 57195 11744 57207 11747
rect 58986 11744 58992 11756
rect 57195 11716 58992 11744
rect 57195 11713 57207 11716
rect 57149 11707 57207 11713
rect 58986 11704 58992 11716
rect 59044 11704 59050 11756
rect 29196 11648 31524 11676
rect 27157 11639 27215 11645
rect 24305 11611 24363 11617
rect 24305 11608 24317 11611
rect 11204 11580 20576 11608
rect 22066 11580 24317 11608
rect 11204 11568 11210 11580
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 12066 11540 12072 11552
rect 11388 11512 12072 11540
rect 11388 11500 11394 11512
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15657 11543 15715 11549
rect 15657 11540 15669 11543
rect 15436 11512 15669 11540
rect 15436 11500 15442 11512
rect 15657 11509 15669 11512
rect 15703 11509 15715 11543
rect 15657 11503 15715 11509
rect 15841 11543 15899 11549
rect 15841 11509 15853 11543
rect 15887 11540 15899 11543
rect 16298 11540 16304 11552
rect 15887 11512 16304 11540
rect 15887 11509 15899 11512
rect 15841 11503 15899 11509
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 16482 11500 16488 11552
rect 16540 11540 16546 11552
rect 19518 11540 19524 11552
rect 16540 11512 19524 11540
rect 16540 11500 16546 11512
rect 19518 11500 19524 11512
rect 19576 11500 19582 11552
rect 19886 11500 19892 11552
rect 19944 11540 19950 11552
rect 19981 11543 20039 11549
rect 19981 11540 19993 11543
rect 19944 11512 19993 11540
rect 19944 11500 19950 11512
rect 19981 11509 19993 11512
rect 20027 11509 20039 11543
rect 19981 11503 20039 11509
rect 20070 11500 20076 11552
rect 20128 11540 20134 11552
rect 22066 11540 22094 11580
rect 24305 11577 24317 11580
rect 24351 11577 24363 11611
rect 24305 11571 24363 11577
rect 24394 11568 24400 11620
rect 24452 11608 24458 11620
rect 27172 11608 27200 11639
rect 32030 11636 32036 11688
rect 32088 11676 32094 11688
rect 33045 11679 33103 11685
rect 33045 11676 33057 11679
rect 32088 11648 33057 11676
rect 32088 11636 32094 11648
rect 33045 11645 33057 11648
rect 33091 11645 33103 11679
rect 33045 11639 33103 11645
rect 41322 11636 41328 11688
rect 41380 11676 41386 11688
rect 43438 11676 43444 11688
rect 41380 11648 43444 11676
rect 41380 11636 41386 11648
rect 43438 11636 43444 11648
rect 43496 11636 43502 11688
rect 43990 11636 43996 11688
rect 44048 11676 44054 11688
rect 46750 11676 46756 11688
rect 44048 11648 46756 11676
rect 44048 11636 44054 11648
rect 46750 11636 46756 11648
rect 46808 11636 46814 11688
rect 46845 11679 46903 11685
rect 46845 11645 46857 11679
rect 46891 11676 46903 11679
rect 46934 11676 46940 11688
rect 46891 11648 46940 11676
rect 46891 11645 46903 11648
rect 46845 11639 46903 11645
rect 46934 11636 46940 11648
rect 46992 11636 46998 11688
rect 24452 11580 27200 11608
rect 24452 11568 24458 11580
rect 28626 11568 28632 11620
rect 28684 11608 28690 11620
rect 40037 11611 40095 11617
rect 40037 11608 40049 11611
rect 28684 11580 31754 11608
rect 28684 11568 28690 11580
rect 20128 11512 22094 11540
rect 20128 11500 20134 11512
rect 25682 11500 25688 11552
rect 25740 11540 25746 11552
rect 28537 11543 28595 11549
rect 28537 11540 28549 11543
rect 25740 11512 28549 11540
rect 25740 11500 25746 11512
rect 28537 11509 28549 11512
rect 28583 11540 28595 11543
rect 29270 11540 29276 11552
rect 28583 11512 29276 11540
rect 28583 11509 28595 11512
rect 28537 11503 28595 11509
rect 29270 11500 29276 11512
rect 29328 11500 29334 11552
rect 29362 11500 29368 11552
rect 29420 11500 29426 11552
rect 30742 11500 30748 11552
rect 30800 11500 30806 11552
rect 31726 11540 31754 11580
rect 35912 11580 40049 11608
rect 35912 11540 35940 11580
rect 40037 11577 40049 11580
rect 40083 11608 40095 11611
rect 44174 11608 44180 11620
rect 40083 11580 44180 11608
rect 40083 11577 40095 11580
rect 40037 11571 40095 11577
rect 44174 11568 44180 11580
rect 44232 11568 44238 11620
rect 45462 11568 45468 11620
rect 45520 11608 45526 11620
rect 45520 11580 51074 11608
rect 45520 11568 45526 11580
rect 31726 11512 35940 11540
rect 35986 11500 35992 11552
rect 36044 11500 36050 11552
rect 36630 11500 36636 11552
rect 36688 11540 36694 11552
rect 46198 11540 46204 11552
rect 36688 11512 46204 11540
rect 36688 11500 36694 11512
rect 46198 11500 46204 11512
rect 46256 11500 46262 11552
rect 46290 11500 46296 11552
rect 46348 11500 46354 11552
rect 51046 11540 51074 11580
rect 52086 11540 52092 11552
rect 51046 11512 52092 11540
rect 52086 11500 52092 11512
rect 52144 11500 52150 11552
rect 57238 11500 57244 11552
rect 57296 11500 57302 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 15194 11336 15200 11348
rect 11256 11308 15200 11336
rect 934 11160 940 11212
rect 992 11200 998 11212
rect 1765 11203 1823 11209
rect 1765 11200 1777 11203
rect 992 11172 1777 11200
rect 992 11160 998 11172
rect 1765 11169 1777 11172
rect 1811 11169 1823 11203
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 1765 11163 1823 11169
rect 2746 11172 10977 11200
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11132 1639 11135
rect 2746 11132 2774 11172
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 11146 11160 11152 11212
rect 11204 11160 11210 11212
rect 11256 11209 11284 11308
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 15746 11296 15752 11348
rect 15804 11336 15810 11348
rect 18785 11339 18843 11345
rect 18785 11336 18797 11339
rect 15804 11308 18797 11336
rect 15804 11296 15810 11308
rect 18785 11305 18797 11308
rect 18831 11305 18843 11339
rect 18785 11299 18843 11305
rect 19150 11296 19156 11348
rect 19208 11336 19214 11348
rect 19208 11308 20760 11336
rect 19208 11296 19214 11308
rect 11790 11228 11796 11280
rect 11848 11268 11854 11280
rect 15105 11271 15163 11277
rect 15105 11268 15117 11271
rect 11848 11240 15117 11268
rect 11848 11228 11854 11240
rect 15105 11237 15117 11240
rect 15151 11237 15163 11271
rect 16482 11268 16488 11280
rect 15105 11231 15163 11237
rect 15212 11240 16488 11268
rect 11241 11203 11299 11209
rect 11241 11169 11253 11203
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11330 11160 11336 11212
rect 11388 11160 11394 11212
rect 11882 11160 11888 11212
rect 11940 11200 11946 11212
rect 11940 11172 13124 11200
rect 11940 11160 11946 11172
rect 1627 11104 2774 11132
rect 1627 11101 1639 11104
rect 1581 11095 1639 11101
rect 11422 11092 11428 11144
rect 11480 11092 11486 11144
rect 12989 11135 13047 11141
rect 12989 11132 13001 11135
rect 12406 11104 13001 11132
rect 8938 11024 8944 11076
rect 8996 11064 9002 11076
rect 12406 11064 12434 11104
rect 12989 11101 13001 11104
rect 13035 11101 13047 11135
rect 13096 11132 13124 11172
rect 13170 11160 13176 11212
rect 13228 11160 13234 11212
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 15212 11200 15240 11240
rect 16482 11228 16488 11240
rect 16540 11228 16546 11280
rect 16684 11240 16896 11268
rect 13872 11172 15240 11200
rect 16393 11203 16451 11209
rect 13872 11160 13878 11172
rect 16393 11169 16405 11203
rect 16439 11200 16451 11203
rect 16684 11200 16712 11240
rect 16439 11172 16712 11200
rect 16868 11200 16896 11240
rect 17494 11228 17500 11280
rect 17552 11268 17558 11280
rect 19426 11268 19432 11280
rect 17552 11240 19432 11268
rect 17552 11228 17558 11240
rect 19426 11228 19432 11240
rect 19484 11228 19490 11280
rect 19242 11200 19248 11212
rect 16868 11172 19248 11200
rect 16439 11169 16451 11172
rect 16393 11163 16451 11169
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 20732 11200 20760 11308
rect 20990 11296 20996 11348
rect 21048 11296 21054 11348
rect 21082 11296 21088 11348
rect 21140 11336 21146 11348
rect 25682 11336 25688 11348
rect 21140 11308 25688 11336
rect 21140 11296 21146 11308
rect 25682 11296 25688 11308
rect 25740 11296 25746 11348
rect 26418 11296 26424 11348
rect 26476 11296 26482 11348
rect 29638 11336 29644 11348
rect 26896 11308 29644 11336
rect 20806 11228 20812 11280
rect 20864 11268 20870 11280
rect 21637 11271 21695 11277
rect 21637 11268 21649 11271
rect 20864 11240 21649 11268
rect 20864 11228 20870 11240
rect 21637 11237 21649 11240
rect 21683 11237 21695 11271
rect 21637 11231 21695 11237
rect 23934 11228 23940 11280
rect 23992 11268 23998 11280
rect 24762 11268 24768 11280
rect 23992 11240 24768 11268
rect 23992 11228 23998 11240
rect 24762 11228 24768 11240
rect 24820 11228 24826 11280
rect 24946 11228 24952 11280
rect 25004 11268 25010 11280
rect 26896 11268 26924 11308
rect 29638 11296 29644 11308
rect 29696 11296 29702 11348
rect 31202 11296 31208 11348
rect 31260 11336 31266 11348
rect 31662 11336 31668 11348
rect 31260 11308 31668 11336
rect 31260 11296 31266 11308
rect 31662 11296 31668 11308
rect 31720 11296 31726 11348
rect 33410 11296 33416 11348
rect 33468 11336 33474 11348
rect 34146 11336 34152 11348
rect 33468 11308 34152 11336
rect 33468 11296 33474 11308
rect 34146 11296 34152 11308
rect 34204 11296 34210 11348
rect 35253 11339 35311 11345
rect 35253 11305 35265 11339
rect 35299 11336 35311 11339
rect 35342 11336 35348 11348
rect 35299 11308 35348 11336
rect 35299 11305 35311 11308
rect 35253 11299 35311 11305
rect 35342 11296 35348 11308
rect 35400 11296 35406 11348
rect 35526 11296 35532 11348
rect 35584 11336 35590 11348
rect 41322 11336 41328 11348
rect 35584 11308 41328 11336
rect 35584 11296 35590 11308
rect 41322 11296 41328 11308
rect 41380 11296 41386 11348
rect 42610 11336 42616 11348
rect 41432 11308 42616 11336
rect 25004 11240 26924 11268
rect 25004 11228 25010 11240
rect 26970 11228 26976 11280
rect 27028 11268 27034 11280
rect 31297 11271 31355 11277
rect 27028 11240 30236 11268
rect 27028 11228 27034 11240
rect 25314 11200 25320 11212
rect 20732 11172 25320 11200
rect 14921 11135 14979 11141
rect 14921 11132 14933 11135
rect 13096 11104 14933 11132
rect 12989 11095 13047 11101
rect 14921 11101 14933 11104
rect 14967 11132 14979 11135
rect 14967 11104 15792 11132
rect 14967 11101 14979 11104
rect 14921 11095 14979 11101
rect 8996 11036 12434 11064
rect 8996 11024 9002 11036
rect 15654 11024 15660 11076
rect 15712 11024 15718 11076
rect 15764 11064 15792 11104
rect 16298 11092 16304 11144
rect 16356 11092 16362 11144
rect 16666 11092 16672 11144
rect 16724 11092 16730 11144
rect 16850 11092 16856 11144
rect 16908 11092 16914 11144
rect 17032 11104 17632 11132
rect 17032 11064 17060 11104
rect 15764 11036 17060 11064
rect 17494 11024 17500 11076
rect 17552 11024 17558 11076
rect 17604 11064 17632 11104
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 18601 11135 18659 11141
rect 18601 11132 18613 11135
rect 18288 11104 18613 11132
rect 18288 11092 18294 11104
rect 18601 11101 18613 11104
rect 18647 11101 18659 11135
rect 18601 11095 18659 11101
rect 19426 11092 19432 11144
rect 19484 11132 19490 11144
rect 21468 11141 21496 11172
rect 25314 11160 25320 11172
rect 25372 11160 25378 11212
rect 26786 11160 26792 11212
rect 26844 11200 26850 11212
rect 27801 11203 27859 11209
rect 27801 11200 27813 11203
rect 26844 11172 27813 11200
rect 26844 11160 26850 11172
rect 27801 11169 27813 11172
rect 27847 11169 27859 11203
rect 27801 11163 27859 11169
rect 29546 11160 29552 11212
rect 29604 11200 29610 11212
rect 30101 11203 30159 11209
rect 30101 11200 30113 11203
rect 29604 11172 30113 11200
rect 29604 11160 29610 11172
rect 30101 11169 30113 11172
rect 30147 11169 30159 11203
rect 30208 11200 30236 11240
rect 31297 11237 31309 11271
rect 31343 11268 31355 11271
rect 32398 11268 32404 11280
rect 31343 11240 32404 11268
rect 31343 11237 31355 11240
rect 31297 11231 31355 11237
rect 32398 11228 32404 11240
rect 32456 11228 32462 11280
rect 32490 11228 32496 11280
rect 32548 11268 32554 11280
rect 33134 11268 33140 11280
rect 32548 11240 33140 11268
rect 32548 11228 32554 11240
rect 33134 11228 33140 11240
rect 33192 11268 33198 11280
rect 39206 11268 39212 11280
rect 33192 11240 33456 11268
rect 33192 11228 33198 11240
rect 33428 11209 33456 11240
rect 37384 11240 39212 11268
rect 33413 11203 33471 11209
rect 30208 11172 32996 11200
rect 30101 11163 30159 11169
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 19484 11104 19625 11132
rect 19484 11092 19490 11104
rect 19613 11101 19625 11104
rect 19659 11132 19671 11135
rect 21453 11135 21511 11141
rect 19659 11104 20300 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 19886 11073 19892 11076
rect 19869 11067 19892 11073
rect 17604 11036 19840 11064
rect 12802 10956 12808 11008
rect 12860 10996 12866 11008
rect 13078 10996 13084 11008
rect 12860 10968 13084 10996
rect 12860 10956 12866 10968
rect 13078 10956 13084 10968
rect 13136 10956 13142 11008
rect 17402 10956 17408 11008
rect 17460 10996 17466 11008
rect 17589 10999 17647 11005
rect 17589 10996 17601 10999
rect 17460 10968 17601 10996
rect 17460 10956 17466 10968
rect 17589 10965 17601 10968
rect 17635 10965 17647 10999
rect 17589 10959 17647 10965
rect 17678 10956 17684 11008
rect 17736 10996 17742 11008
rect 19610 10996 19616 11008
rect 17736 10968 19616 10996
rect 17736 10956 17742 10968
rect 19610 10956 19616 10968
rect 19668 10956 19674 11008
rect 19812 10996 19840 11036
rect 19869 11033 19881 11067
rect 19869 11027 19892 11033
rect 19886 11024 19892 11027
rect 19944 11024 19950 11076
rect 20272 11064 20300 11104
rect 21453 11101 21465 11135
rect 21499 11101 21511 11135
rect 21453 11095 21511 11101
rect 21634 11092 21640 11144
rect 21692 11132 21698 11144
rect 22002 11132 22008 11144
rect 21692 11104 22008 11132
rect 21692 11092 21698 11104
rect 22002 11092 22008 11104
rect 22060 11132 22066 11144
rect 24765 11135 24823 11141
rect 24765 11132 24777 11135
rect 22060 11104 24777 11132
rect 22060 11092 22066 11104
rect 24765 11101 24777 11104
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 25130 11092 25136 11144
rect 25188 11132 25194 11144
rect 26237 11135 26295 11141
rect 26237 11132 26249 11135
rect 25188 11104 26249 11132
rect 25188 11092 25194 11104
rect 26237 11101 26249 11104
rect 26283 11132 26295 11135
rect 27154 11132 27160 11144
rect 26283 11104 27160 11132
rect 26283 11101 26295 11104
rect 26237 11095 26295 11101
rect 27154 11092 27160 11104
rect 27212 11092 27218 11144
rect 27338 11092 27344 11144
rect 27396 11092 27402 11144
rect 27430 11092 27436 11144
rect 27488 11132 27494 11144
rect 29733 11135 29791 11141
rect 29733 11132 29745 11135
rect 27488 11104 29745 11132
rect 27488 11092 27494 11104
rect 29733 11101 29745 11104
rect 29779 11101 29791 11135
rect 30650 11132 30656 11144
rect 29733 11095 29791 11101
rect 29840 11104 30656 11132
rect 24394 11064 24400 11076
rect 20272 11036 24400 11064
rect 24394 11024 24400 11036
rect 24452 11024 24458 11076
rect 24670 11024 24676 11076
rect 24728 11064 24734 11076
rect 25593 11067 25651 11073
rect 25593 11064 25605 11067
rect 24728 11036 25605 11064
rect 24728 11024 24734 11036
rect 25593 11033 25605 11036
rect 25639 11064 25651 11067
rect 27522 11064 27528 11076
rect 25639 11036 27528 11064
rect 25639 11033 25651 11036
rect 25593 11027 25651 11033
rect 27522 11024 27528 11036
rect 27580 11064 27586 11076
rect 28074 11064 28080 11076
rect 27580 11036 28080 11064
rect 27580 11024 27586 11036
rect 28074 11024 28080 11036
rect 28132 11024 28138 11076
rect 28258 11024 28264 11076
rect 28316 11064 28322 11076
rect 29840 11064 29868 11104
rect 30650 11092 30656 11104
rect 30708 11132 30714 11144
rect 31573 11135 31631 11141
rect 31573 11132 31585 11135
rect 30708 11104 31585 11132
rect 30708 11092 30714 11104
rect 31573 11101 31585 11104
rect 31619 11132 31631 11135
rect 31662 11132 31668 11144
rect 31619 11104 31668 11132
rect 31619 11101 31631 11104
rect 31573 11095 31631 11101
rect 31662 11092 31668 11104
rect 31720 11092 31726 11144
rect 31846 11092 31852 11144
rect 31904 11132 31910 11144
rect 32033 11135 32091 11141
rect 32033 11132 32045 11135
rect 31904 11104 32045 11132
rect 31904 11092 31910 11104
rect 32033 11101 32045 11104
rect 32079 11101 32091 11135
rect 32033 11095 32091 11101
rect 32125 11135 32183 11141
rect 32125 11101 32137 11135
rect 32171 11132 32183 11135
rect 32490 11132 32496 11144
rect 32171 11104 32496 11132
rect 32171 11101 32183 11104
rect 32125 11095 32183 11101
rect 32490 11092 32496 11104
rect 32548 11092 32554 11144
rect 32968 11141 32996 11172
rect 33413 11169 33425 11203
rect 33459 11169 33471 11203
rect 33413 11163 33471 11169
rect 35802 11160 35808 11212
rect 35860 11160 35866 11212
rect 35894 11160 35900 11212
rect 35952 11200 35958 11212
rect 36814 11200 36820 11212
rect 35952 11172 36820 11200
rect 35952 11160 35958 11172
rect 36814 11160 36820 11172
rect 36872 11160 36878 11212
rect 32953 11135 33011 11141
rect 32953 11101 32965 11135
rect 32999 11101 33011 11135
rect 32953 11095 33011 11101
rect 33042 11092 33048 11144
rect 33100 11132 33106 11144
rect 33502 11132 33508 11144
rect 33100 11104 33508 11132
rect 33100 11092 33106 11104
rect 33502 11092 33508 11104
rect 33560 11092 33566 11144
rect 35621 11135 35679 11141
rect 35621 11101 35633 11135
rect 35667 11132 35679 11135
rect 37384 11132 37412 11240
rect 39206 11228 39212 11240
rect 39264 11228 39270 11280
rect 38102 11160 38108 11212
rect 38160 11200 38166 11212
rect 38838 11200 38844 11212
rect 38160 11172 38844 11200
rect 38160 11160 38166 11172
rect 38838 11160 38844 11172
rect 38896 11160 38902 11212
rect 41432 11209 41460 11308
rect 42610 11296 42616 11308
rect 42668 11296 42674 11348
rect 46198 11296 46204 11348
rect 46256 11336 46262 11348
rect 57238 11336 57244 11348
rect 46256 11308 57244 11336
rect 46256 11296 46262 11308
rect 57238 11296 57244 11308
rect 57296 11296 57302 11348
rect 46750 11228 46756 11280
rect 46808 11268 46814 11280
rect 46937 11271 46995 11277
rect 46937 11268 46949 11271
rect 46808 11240 46949 11268
rect 46808 11228 46814 11240
rect 46937 11237 46949 11240
rect 46983 11237 46995 11271
rect 46937 11231 46995 11237
rect 53558 11228 53564 11280
rect 53616 11268 53622 11280
rect 53653 11271 53711 11277
rect 53653 11268 53665 11271
rect 53616 11240 53665 11268
rect 53616 11228 53622 11240
rect 53653 11237 53665 11240
rect 53699 11237 53711 11271
rect 53653 11231 53711 11237
rect 56137 11271 56195 11277
rect 56137 11237 56149 11271
rect 56183 11237 56195 11271
rect 56137 11231 56195 11237
rect 41417 11203 41475 11209
rect 41417 11169 41429 11203
rect 41463 11169 41475 11203
rect 41782 11200 41788 11212
rect 41417 11163 41475 11169
rect 41524 11172 41788 11200
rect 35667 11104 37412 11132
rect 35667 11101 35679 11104
rect 35621 11095 35679 11101
rect 38470 11092 38476 11144
rect 38528 11092 38534 11144
rect 41524 11141 41552 11172
rect 41782 11160 41788 11172
rect 41840 11160 41846 11212
rect 42242 11160 42248 11212
rect 42300 11200 42306 11212
rect 42300 11172 43208 11200
rect 42300 11160 42306 11172
rect 41509 11135 41567 11141
rect 38626 11104 41092 11132
rect 28316 11036 29868 11064
rect 28316 11024 28322 11036
rect 30190 11024 30196 11076
rect 30248 11064 30254 11076
rect 30248 11036 31248 11064
rect 30248 11024 30254 11036
rect 20714 10996 20720 11008
rect 19812 10968 20720 10996
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 25498 10956 25504 11008
rect 25556 10996 25562 11008
rect 26050 10996 26056 11008
rect 25556 10968 26056 10996
rect 25556 10956 25562 10968
rect 26050 10956 26056 10968
rect 26108 10996 26114 11008
rect 30650 10996 30656 11008
rect 26108 10968 30656 10996
rect 26108 10956 26114 10968
rect 30650 10956 30656 10968
rect 30708 10956 30714 11008
rect 31220 10996 31248 11036
rect 31294 11024 31300 11076
rect 31352 11064 31358 11076
rect 32858 11064 32864 11076
rect 31352 11036 32864 11064
rect 31352 11024 31358 11036
rect 32858 11024 32864 11036
rect 32916 11024 32922 11076
rect 33318 11024 33324 11076
rect 33376 11064 33382 11076
rect 33778 11064 33784 11076
rect 33376 11036 33784 11064
rect 33376 11024 33382 11036
rect 33778 11024 33784 11036
rect 33836 11024 33842 11076
rect 34422 11024 34428 11076
rect 34480 11064 34486 11076
rect 35713 11067 35771 11073
rect 35713 11064 35725 11067
rect 34480 11036 35725 11064
rect 34480 11024 34486 11036
rect 35713 11033 35725 11036
rect 35759 11064 35771 11067
rect 35986 11064 35992 11076
rect 35759 11036 35992 11064
rect 35759 11033 35771 11036
rect 35713 11027 35771 11033
rect 35986 11024 35992 11036
rect 36044 11024 36050 11076
rect 37366 11024 37372 11076
rect 37424 11064 37430 11076
rect 38289 11067 38347 11073
rect 38289 11064 38301 11067
rect 37424 11036 38301 11064
rect 37424 11024 37430 11036
rect 38289 11033 38301 11036
rect 38335 11033 38347 11067
rect 38289 11027 38347 11033
rect 38378 11024 38384 11076
rect 38436 11064 38442 11076
rect 38626 11064 38654 11104
rect 41064 11076 41092 11104
rect 41509 11101 41521 11135
rect 41555 11101 41567 11135
rect 41509 11095 41567 11101
rect 41877 11135 41935 11141
rect 41877 11101 41889 11135
rect 41923 11132 41935 11135
rect 41966 11132 41972 11144
rect 41923 11104 41972 11132
rect 41923 11101 41935 11104
rect 41877 11095 41935 11101
rect 41966 11092 41972 11104
rect 42024 11092 42030 11144
rect 42061 11135 42119 11141
rect 42061 11101 42073 11135
rect 42107 11132 42119 11135
rect 42978 11132 42984 11144
rect 42107 11104 42984 11132
rect 42107 11101 42119 11104
rect 42061 11095 42119 11101
rect 42978 11092 42984 11104
rect 43036 11132 43042 11144
rect 43180 11141 43208 11172
rect 43254 11160 43260 11212
rect 43312 11160 43318 11212
rect 45462 11200 45468 11212
rect 43548 11172 45468 11200
rect 43548 11141 43576 11172
rect 45462 11160 45468 11172
rect 45520 11160 45526 11212
rect 54202 11200 54208 11212
rect 53116 11172 54208 11200
rect 43165 11135 43223 11141
rect 43036 11104 43116 11132
rect 43036 11092 43042 11104
rect 38436 11036 38654 11064
rect 38841 11067 38899 11073
rect 38436 11024 38442 11036
rect 38841 11033 38853 11067
rect 38887 11064 38899 11067
rect 39022 11064 39028 11076
rect 38887 11036 39028 11064
rect 38887 11033 38899 11036
rect 38841 11027 38899 11033
rect 39022 11024 39028 11036
rect 39080 11024 39086 11076
rect 39390 11024 39396 11076
rect 39448 11064 39454 11076
rect 40218 11064 40224 11076
rect 39448 11036 40224 11064
rect 39448 11024 39454 11036
rect 40218 11024 40224 11036
rect 40276 11024 40282 11076
rect 40494 11024 40500 11076
rect 40552 11064 40558 11076
rect 40865 11067 40923 11073
rect 40865 11064 40877 11067
rect 40552 11036 40877 11064
rect 40552 11024 40558 11036
rect 40865 11033 40877 11036
rect 40911 11064 40923 11067
rect 40954 11064 40960 11076
rect 40911 11036 40960 11064
rect 40911 11033 40923 11036
rect 40865 11027 40923 11033
rect 40954 11024 40960 11036
rect 41012 11024 41018 11076
rect 41046 11024 41052 11076
rect 41104 11064 41110 11076
rect 42334 11064 42340 11076
rect 41104 11036 42340 11064
rect 41104 11024 41110 11036
rect 42334 11024 42340 11036
rect 42392 11024 42398 11076
rect 42518 11024 42524 11076
rect 42576 11024 42582 11076
rect 43088 11064 43116 11104
rect 43165 11101 43177 11135
rect 43211 11101 43223 11135
rect 43165 11095 43223 11101
rect 43533 11135 43591 11141
rect 43533 11101 43545 11135
rect 43579 11101 43591 11135
rect 43533 11095 43591 11101
rect 43625 11135 43683 11141
rect 43625 11101 43637 11135
rect 43671 11101 43683 11135
rect 43625 11095 43683 11101
rect 44177 11135 44235 11141
rect 44177 11101 44189 11135
rect 44223 11132 44235 11135
rect 45557 11135 45615 11141
rect 44223 11104 45508 11132
rect 44223 11101 44235 11104
rect 44177 11095 44235 11101
rect 43640 11064 43668 11095
rect 43088 11036 43668 11064
rect 44450 11024 44456 11076
rect 44508 11024 44514 11076
rect 45480 11064 45508 11104
rect 45557 11101 45569 11135
rect 45603 11132 45615 11135
rect 46934 11132 46940 11144
rect 45603 11104 46940 11132
rect 45603 11101 45615 11104
rect 45557 11095 45615 11101
rect 46934 11092 46940 11104
rect 46992 11132 46998 11144
rect 47762 11132 47768 11144
rect 46992 11104 47768 11132
rect 46992 11092 46998 11104
rect 47762 11092 47768 11104
rect 47820 11092 47826 11144
rect 53116 11141 53144 11172
rect 54202 11160 54208 11172
rect 54260 11160 54266 11212
rect 56152 11200 56180 11231
rect 57882 11228 57888 11280
rect 57940 11268 57946 11280
rect 58253 11271 58311 11277
rect 58253 11268 58265 11271
rect 57940 11240 58265 11268
rect 57940 11228 57946 11240
rect 58253 11237 58265 11240
rect 58299 11237 58311 11271
rect 58253 11231 58311 11237
rect 56152 11172 57008 11200
rect 53101 11135 53159 11141
rect 53101 11101 53113 11135
rect 53147 11101 53159 11135
rect 53101 11095 53159 11101
rect 53190 11092 53196 11144
rect 53248 11132 53254 11144
rect 53285 11135 53343 11141
rect 53285 11132 53297 11135
rect 53248 11104 53297 11132
rect 53248 11092 53254 11104
rect 53285 11101 53297 11104
rect 53331 11101 53343 11135
rect 53285 11095 53343 11101
rect 53466 11092 53472 11144
rect 53524 11092 53530 11144
rect 56134 11092 56140 11144
rect 56192 11092 56198 11144
rect 56410 11092 56416 11144
rect 56468 11092 56474 11144
rect 56870 11092 56876 11144
rect 56928 11092 56934 11144
rect 56980 11132 57008 11172
rect 57129 11135 57187 11141
rect 57129 11132 57141 11135
rect 56980 11104 57141 11132
rect 57129 11101 57141 11104
rect 57175 11101 57187 11135
rect 57129 11095 57187 11101
rect 45824 11067 45882 11073
rect 45480 11036 45784 11064
rect 31481 10999 31539 11005
rect 31481 10996 31493 10999
rect 31220 10968 31493 10996
rect 31481 10965 31493 10968
rect 31527 10965 31539 10999
rect 31481 10959 31539 10965
rect 35894 10956 35900 11008
rect 35952 10996 35958 11008
rect 39942 10996 39948 11008
rect 35952 10968 39948 10996
rect 35952 10956 35958 10968
rect 39942 10956 39948 10968
rect 40000 10956 40006 11008
rect 45756 10996 45784 11036
rect 45824 11033 45836 11067
rect 45870 11064 45882 11067
rect 46290 11064 46296 11076
rect 45870 11036 46296 11064
rect 45870 11033 45882 11036
rect 45824 11027 45882 11033
rect 46290 11024 46296 11036
rect 46348 11024 46354 11076
rect 46658 11064 46664 11076
rect 46400 11036 46664 11064
rect 46400 10996 46428 11036
rect 46658 11024 46664 11036
rect 46716 11024 46722 11076
rect 53377 11067 53435 11073
rect 53377 11033 53389 11067
rect 53423 11064 53435 11067
rect 56042 11064 56048 11076
rect 53423 11036 56048 11064
rect 53423 11033 53435 11036
rect 53377 11027 53435 11033
rect 56042 11024 56048 11036
rect 56100 11024 56106 11076
rect 56321 11067 56379 11073
rect 56321 11033 56333 11067
rect 56367 11064 56379 11067
rect 56962 11064 56968 11076
rect 56367 11036 56968 11064
rect 56367 11033 56379 11036
rect 56321 11027 56379 11033
rect 56962 11024 56968 11036
rect 57020 11024 57026 11076
rect 45756 10968 46428 10996
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 3510 10752 3516 10804
rect 3568 10792 3574 10804
rect 9309 10795 9367 10801
rect 9309 10792 9321 10795
rect 3568 10764 9321 10792
rect 3568 10752 3574 10764
rect 9309 10761 9321 10764
rect 9355 10761 9367 10795
rect 9309 10755 9367 10761
rect 9416 10764 9904 10792
rect 934 10684 940 10736
rect 992 10724 998 10736
rect 1857 10727 1915 10733
rect 1857 10724 1869 10727
rect 992 10696 1869 10724
rect 992 10684 998 10696
rect 1857 10693 1869 10696
rect 1903 10693 1915 10727
rect 9416 10724 9444 10764
rect 1857 10687 1915 10693
rect 9324 10696 9444 10724
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10656 1639 10659
rect 9324 10656 9352 10696
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 9876 10724 9904 10764
rect 12158 10752 12164 10804
rect 12216 10752 12222 10804
rect 17678 10792 17684 10804
rect 12406 10764 17684 10792
rect 12406 10724 12434 10764
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 18509 10795 18567 10801
rect 18509 10761 18521 10795
rect 18555 10761 18567 10795
rect 18509 10755 18567 10761
rect 18877 10795 18935 10801
rect 18877 10761 18889 10795
rect 18923 10792 18935 10795
rect 19334 10792 19340 10804
rect 18923 10764 19340 10792
rect 18923 10761 18935 10764
rect 18877 10755 18935 10761
rect 17037 10727 17095 10733
rect 9732 10696 9812 10724
rect 9876 10696 12434 10724
rect 12912 10696 14136 10724
rect 9732 10684 9738 10696
rect 1627 10628 9352 10656
rect 1627 10625 1639 10628
rect 1581 10619 1639 10625
rect 9490 10616 9496 10668
rect 9548 10616 9554 10668
rect 9582 10616 9588 10668
rect 9640 10616 9646 10668
rect 9784 10665 9812 10696
rect 9769 10659 9827 10665
rect 9769 10625 9781 10659
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 11330 10616 11336 10668
rect 11388 10656 11394 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11388 10628 11713 10656
rect 11388 10616 11394 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 12802 10616 12808 10668
rect 12860 10656 12866 10668
rect 12912 10665 12940 10696
rect 12897 10659 12955 10665
rect 12897 10656 12909 10659
rect 12860 10628 12909 10656
rect 12860 10616 12866 10628
rect 12897 10625 12909 10628
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10656 13231 10659
rect 13998 10656 14004 10668
rect 13219 10628 14004 10656
rect 13219 10625 13231 10628
rect 13173 10619 13231 10625
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 9677 10591 9735 10597
rect 1728 10560 9628 10588
rect 1728 10548 1734 10560
rect 9600 10520 9628 10560
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 11348 10588 11376 10616
rect 13357 10591 13415 10597
rect 13357 10588 13369 10591
rect 9723 10560 11376 10588
rect 11808 10560 13369 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 11808 10520 11836 10560
rect 13357 10557 13369 10560
rect 13403 10557 13415 10591
rect 13357 10551 13415 10557
rect 9600 10492 11836 10520
rect 11977 10523 12035 10529
rect 11977 10489 11989 10523
rect 12023 10489 12035 10523
rect 11977 10483 12035 10489
rect 12989 10523 13047 10529
rect 12989 10489 13001 10523
rect 13035 10520 13047 10523
rect 13170 10520 13176 10532
rect 13035 10492 13176 10520
rect 13035 10489 13047 10492
rect 12989 10483 13047 10489
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 10962 10452 10968 10464
rect 9640 10424 10968 10452
rect 9640 10412 9646 10424
rect 10962 10412 10968 10424
rect 11020 10412 11026 10464
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 11992 10452 12020 10483
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 14108 10520 14136 10696
rect 17037 10693 17049 10727
rect 17083 10724 17095 10727
rect 18524 10724 18552 10755
rect 19334 10752 19340 10764
rect 19392 10792 19398 10804
rect 21085 10795 21143 10801
rect 21085 10792 21097 10795
rect 19392 10764 21097 10792
rect 19392 10752 19398 10764
rect 21085 10761 21097 10764
rect 21131 10761 21143 10795
rect 22005 10795 22063 10801
rect 22005 10792 22017 10795
rect 21085 10755 21143 10761
rect 21192 10764 22017 10792
rect 19950 10727 20008 10733
rect 19950 10724 19962 10727
rect 17083 10696 18460 10724
rect 18524 10696 19962 10724
rect 17083 10693 17095 10696
rect 17037 10687 17095 10693
rect 14734 10616 14740 10668
rect 14792 10616 14798 10668
rect 14918 10616 14924 10668
rect 14976 10616 14982 10668
rect 15657 10659 15715 10665
rect 15657 10625 15669 10659
rect 15703 10656 15715 10659
rect 17218 10656 17224 10668
rect 15703 10628 17224 10656
rect 15703 10625 15715 10628
rect 15657 10619 15715 10625
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 17402 10616 17408 10668
rect 17460 10616 17466 10668
rect 17494 10616 17500 10668
rect 17552 10616 17558 10668
rect 18432 10656 18460 10696
rect 19950 10693 19962 10696
rect 19996 10693 20008 10727
rect 19950 10687 20008 10693
rect 20530 10684 20536 10736
rect 20588 10724 20594 10736
rect 21192 10724 21220 10764
rect 22005 10761 22017 10764
rect 22051 10761 22063 10795
rect 22005 10755 22063 10761
rect 22278 10752 22284 10804
rect 22336 10792 22342 10804
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 22336 10764 22385 10792
rect 22336 10752 22342 10764
rect 22373 10761 22385 10764
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 23569 10795 23627 10801
rect 23569 10761 23581 10795
rect 23615 10792 23627 10795
rect 31205 10795 31263 10801
rect 31205 10792 31217 10795
rect 23615 10764 31217 10792
rect 23615 10761 23627 10764
rect 23569 10755 23627 10761
rect 31205 10761 31217 10764
rect 31251 10761 31263 10795
rect 31205 10755 31263 10761
rect 32950 10752 32956 10804
rect 33008 10792 33014 10804
rect 33781 10795 33839 10801
rect 33781 10792 33793 10795
rect 33008 10764 33793 10792
rect 33008 10752 33014 10764
rect 33781 10761 33793 10764
rect 33827 10761 33839 10795
rect 33781 10755 33839 10761
rect 34330 10752 34336 10804
rect 34388 10792 34394 10804
rect 34388 10764 34468 10792
rect 34388 10752 34394 10764
rect 20588 10696 21220 10724
rect 20588 10684 20594 10696
rect 21450 10684 21456 10736
rect 21508 10724 21514 10736
rect 26329 10727 26387 10733
rect 26329 10724 26341 10727
rect 21508 10696 26341 10724
rect 21508 10684 21514 10696
rect 18432 10628 19104 10656
rect 15470 10548 15476 10600
rect 15528 10588 15534 10600
rect 15930 10588 15936 10600
rect 15528 10560 15936 10588
rect 15528 10548 15534 10560
rect 15930 10548 15936 10560
rect 15988 10548 15994 10600
rect 16942 10548 16948 10600
rect 17000 10548 17006 10600
rect 17957 10591 18015 10597
rect 17957 10588 17969 10591
rect 17052 10560 17969 10588
rect 15105 10523 15163 10529
rect 15105 10520 15117 10523
rect 14108 10492 15117 10520
rect 15105 10489 15117 10492
rect 15151 10489 15163 10523
rect 15105 10483 15163 10489
rect 16114 10480 16120 10532
rect 16172 10520 16178 10532
rect 17052 10520 17080 10560
rect 17957 10557 17969 10560
rect 18003 10588 18015 10591
rect 18414 10588 18420 10600
rect 18003 10560 18420 10588
rect 18003 10557 18015 10560
rect 17957 10551 18015 10557
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 18598 10548 18604 10600
rect 18656 10588 18662 10600
rect 18969 10591 19027 10597
rect 18969 10588 18981 10591
rect 18656 10560 18981 10588
rect 18656 10548 18662 10560
rect 18969 10557 18981 10560
rect 19015 10557 19027 10591
rect 18969 10551 19027 10557
rect 16172 10492 17080 10520
rect 16172 10480 16178 10492
rect 17218 10480 17224 10532
rect 17276 10520 17282 10532
rect 18506 10520 18512 10532
rect 17276 10492 18512 10520
rect 17276 10480 17282 10492
rect 18506 10480 18512 10492
rect 18564 10480 18570 10532
rect 19076 10520 19104 10628
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19705 10659 19763 10665
rect 19705 10656 19717 10659
rect 19484 10628 19717 10656
rect 19484 10616 19490 10628
rect 19705 10625 19717 10628
rect 19751 10625 19763 10659
rect 20898 10656 20904 10668
rect 19705 10619 19763 10625
rect 19812 10628 20904 10656
rect 19153 10591 19211 10597
rect 19153 10557 19165 10591
rect 19199 10588 19211 10591
rect 19812 10588 19840 10628
rect 20898 10616 20904 10628
rect 20956 10616 20962 10668
rect 23385 10659 23443 10665
rect 23385 10625 23397 10659
rect 23431 10625 23443 10659
rect 23385 10619 23443 10625
rect 23569 10659 23627 10665
rect 23569 10625 23581 10659
rect 23615 10656 23627 10659
rect 23750 10656 23756 10668
rect 23615 10628 23756 10656
rect 23615 10625 23627 10628
rect 23569 10619 23627 10625
rect 19199 10560 19840 10588
rect 19199 10557 19211 10560
rect 19153 10551 19211 10557
rect 21082 10548 21088 10600
rect 21140 10588 21146 10600
rect 22465 10591 22523 10597
rect 22465 10588 22477 10591
rect 21140 10560 22477 10588
rect 21140 10548 21146 10560
rect 22465 10557 22477 10560
rect 22511 10557 22523 10591
rect 22465 10551 22523 10557
rect 22557 10591 22615 10597
rect 22557 10557 22569 10591
rect 22603 10557 22615 10591
rect 23400 10588 23428 10619
rect 23750 10616 23756 10628
rect 23808 10616 23814 10668
rect 24504 10665 24532 10696
rect 26329 10693 26341 10696
rect 26375 10724 26387 10727
rect 27798 10724 27804 10736
rect 26375 10696 27804 10724
rect 26375 10693 26387 10696
rect 26329 10687 26387 10693
rect 27798 10684 27804 10696
rect 27856 10684 27862 10736
rect 31754 10724 31760 10736
rect 29472 10696 31760 10724
rect 24489 10659 24547 10665
rect 24489 10625 24501 10659
rect 24535 10625 24547 10659
rect 24489 10619 24547 10625
rect 24857 10659 24915 10665
rect 24857 10625 24869 10659
rect 24903 10656 24915 10659
rect 25685 10659 25743 10665
rect 24903 10628 25452 10656
rect 24903 10625 24915 10628
rect 24857 10619 24915 10625
rect 23842 10588 23848 10600
rect 23400 10560 23848 10588
rect 22557 10551 22615 10557
rect 19702 10520 19708 10532
rect 19076 10492 19708 10520
rect 19702 10480 19708 10492
rect 19760 10480 19766 10532
rect 21818 10480 21824 10532
rect 21876 10520 21882 10532
rect 22572 10520 22600 10551
rect 23842 10548 23848 10560
rect 23900 10588 23906 10600
rect 24118 10588 24124 10600
rect 23900 10560 24124 10588
rect 23900 10548 23906 10560
rect 24118 10548 24124 10560
rect 24176 10548 24182 10600
rect 24946 10548 24952 10600
rect 25004 10548 25010 10600
rect 25424 10588 25452 10628
rect 25685 10625 25697 10659
rect 25731 10656 25743 10659
rect 25731 10628 25912 10656
rect 25731 10625 25743 10628
rect 25685 10619 25743 10625
rect 25774 10588 25780 10600
rect 25424 10560 25780 10588
rect 25774 10548 25780 10560
rect 25832 10548 25838 10600
rect 21876 10492 22600 10520
rect 21876 10480 21882 10492
rect 24302 10480 24308 10532
rect 24360 10480 24366 10532
rect 24486 10480 24492 10532
rect 24544 10520 24550 10532
rect 25884 10520 25912 10628
rect 27062 10616 27068 10668
rect 27120 10656 27126 10668
rect 27614 10656 27620 10668
rect 27120 10628 27620 10656
rect 27120 10616 27126 10628
rect 27614 10616 27620 10628
rect 27672 10656 27678 10668
rect 27709 10659 27767 10665
rect 27709 10656 27721 10659
rect 27672 10628 27721 10656
rect 27672 10616 27678 10628
rect 27709 10625 27721 10628
rect 27755 10625 27767 10659
rect 27709 10619 27767 10625
rect 27890 10616 27896 10668
rect 27948 10616 27954 10668
rect 28077 10659 28135 10665
rect 28077 10625 28089 10659
rect 28123 10656 28135 10659
rect 28258 10656 28264 10668
rect 28123 10628 28264 10656
rect 28123 10625 28135 10628
rect 28077 10619 28135 10625
rect 28258 10616 28264 10628
rect 28316 10616 28322 10668
rect 28534 10616 28540 10668
rect 28592 10665 28598 10668
rect 28592 10619 28602 10665
rect 28592 10616 28598 10619
rect 28810 10616 28816 10668
rect 28868 10616 28874 10668
rect 29472 10656 29500 10696
rect 31754 10684 31760 10696
rect 31812 10724 31818 10736
rect 34440 10733 34468 10764
rect 34606 10752 34612 10804
rect 34664 10752 34670 10804
rect 34793 10795 34851 10801
rect 34793 10761 34805 10795
rect 34839 10792 34851 10795
rect 34839 10764 35296 10792
rect 34839 10761 34851 10764
rect 34793 10755 34851 10761
rect 34425 10727 34483 10733
rect 31812 10696 34376 10724
rect 31812 10684 31818 10696
rect 28966 10628 29500 10656
rect 27798 10548 27804 10600
rect 27856 10588 27862 10600
rect 28966 10588 28994 10628
rect 31018 10616 31024 10668
rect 31076 10656 31082 10668
rect 31146 10659 31204 10665
rect 31146 10656 31158 10659
rect 31076 10628 31158 10656
rect 31076 10616 31082 10628
rect 31146 10625 31158 10628
rect 31192 10625 31204 10659
rect 31146 10619 31204 10625
rect 33134 10616 33140 10668
rect 33192 10616 33198 10668
rect 33318 10665 33324 10668
rect 33285 10659 33324 10665
rect 33285 10625 33297 10659
rect 33285 10619 33324 10625
rect 33318 10616 33324 10619
rect 33376 10616 33382 10668
rect 33410 10616 33416 10668
rect 33468 10616 33474 10668
rect 33502 10616 33508 10668
rect 33560 10616 33566 10668
rect 33643 10659 33701 10665
rect 33643 10625 33655 10659
rect 33689 10656 33701 10659
rect 33870 10656 33876 10668
rect 33689 10628 33876 10656
rect 33689 10625 33701 10628
rect 33643 10619 33701 10625
rect 33870 10616 33876 10628
rect 33928 10616 33934 10668
rect 34238 10616 34244 10668
rect 34296 10616 34302 10668
rect 34348 10656 34376 10696
rect 34425 10693 34437 10727
rect 34471 10693 34483 10727
rect 34425 10687 34483 10693
rect 34517 10727 34575 10733
rect 34517 10693 34529 10727
rect 34563 10724 34575 10727
rect 34624 10724 34652 10752
rect 35268 10733 35296 10764
rect 35342 10752 35348 10804
rect 35400 10792 35406 10804
rect 36170 10792 36176 10804
rect 35400 10764 36176 10792
rect 35400 10752 35406 10764
rect 36170 10752 36176 10764
rect 36228 10752 36234 10804
rect 40678 10752 40684 10804
rect 40736 10792 40742 10804
rect 45186 10792 45192 10804
rect 40736 10764 45192 10792
rect 40736 10752 40742 10764
rect 45186 10752 45192 10764
rect 45244 10792 45250 10804
rect 45465 10795 45523 10801
rect 45465 10792 45477 10795
rect 45244 10764 45477 10792
rect 45244 10752 45250 10764
rect 45465 10761 45477 10764
rect 45511 10761 45523 10795
rect 45465 10755 45523 10761
rect 56962 10752 56968 10804
rect 57020 10792 57026 10804
rect 57241 10795 57299 10801
rect 57241 10792 57253 10795
rect 57020 10764 57253 10792
rect 57020 10752 57026 10764
rect 57241 10761 57253 10764
rect 57287 10761 57299 10795
rect 57241 10755 57299 10761
rect 34563 10696 34652 10724
rect 35253 10727 35311 10733
rect 34563 10693 34575 10696
rect 34517 10687 34575 10693
rect 35253 10693 35265 10727
rect 35299 10693 35311 10727
rect 37550 10724 37556 10736
rect 35253 10687 35311 10693
rect 35360 10696 37556 10724
rect 34609 10659 34667 10665
rect 34609 10656 34621 10659
rect 34348 10628 34621 10656
rect 34609 10625 34621 10628
rect 34655 10625 34667 10659
rect 34609 10619 34667 10625
rect 35158 10616 35164 10668
rect 35216 10656 35222 10668
rect 35360 10656 35388 10696
rect 37550 10684 37556 10696
rect 37608 10724 37614 10736
rect 38197 10727 38255 10733
rect 38197 10724 38209 10727
rect 37608 10696 38209 10724
rect 37608 10684 37614 10696
rect 38197 10693 38209 10696
rect 38243 10693 38255 10727
rect 38197 10687 38255 10693
rect 38289 10727 38347 10733
rect 38289 10693 38301 10727
rect 38335 10724 38347 10727
rect 55766 10724 55772 10736
rect 38335 10696 55772 10724
rect 38335 10693 38347 10696
rect 38289 10687 38347 10693
rect 55766 10684 55772 10696
rect 55824 10684 55830 10736
rect 35216 10628 35388 10656
rect 35216 10616 35222 10628
rect 35434 10616 35440 10668
rect 35492 10616 35498 10668
rect 35529 10659 35587 10665
rect 35529 10625 35541 10659
rect 35575 10625 35587 10659
rect 35529 10619 35587 10625
rect 38013 10659 38071 10665
rect 38013 10625 38025 10659
rect 38059 10625 38071 10659
rect 38013 10619 38071 10625
rect 27856 10560 28304 10588
rect 27856 10548 27862 10560
rect 24544 10492 25912 10520
rect 24544 10480 24550 10492
rect 27154 10480 27160 10532
rect 27212 10520 27218 10532
rect 28276 10520 28304 10560
rect 28552 10560 28994 10588
rect 28552 10520 28580 10560
rect 29270 10548 29276 10600
rect 29328 10588 29334 10600
rect 31573 10591 31631 10597
rect 31573 10588 31585 10591
rect 29328 10560 31585 10588
rect 29328 10548 29334 10560
rect 31573 10557 31585 10560
rect 31619 10557 31631 10591
rect 31573 10551 31631 10557
rect 31665 10591 31723 10597
rect 31665 10557 31677 10591
rect 31711 10588 31723 10591
rect 32582 10588 32588 10600
rect 31711 10560 32588 10588
rect 31711 10557 31723 10560
rect 31665 10551 31723 10557
rect 32582 10548 32588 10560
rect 32640 10548 32646 10600
rect 32674 10548 32680 10600
rect 32732 10588 32738 10600
rect 35544 10588 35572 10619
rect 32732 10560 35572 10588
rect 38028 10588 38056 10619
rect 38378 10616 38384 10668
rect 38436 10616 38442 10668
rect 40948 10659 41006 10665
rect 40948 10625 40960 10659
rect 40994 10656 41006 10659
rect 41322 10656 41328 10668
rect 40994 10628 41328 10656
rect 40994 10625 41006 10628
rect 40948 10619 41006 10625
rect 41322 10616 41328 10628
rect 41380 10616 41386 10668
rect 44174 10616 44180 10668
rect 44232 10656 44238 10668
rect 44818 10656 44824 10668
rect 44232 10628 44824 10656
rect 44232 10616 44238 10628
rect 44818 10616 44824 10628
rect 44876 10616 44882 10668
rect 56778 10616 56784 10668
rect 56836 10656 56842 10668
rect 57149 10659 57207 10665
rect 57149 10656 57161 10659
rect 56836 10628 57161 10656
rect 56836 10616 56842 10628
rect 57149 10625 57161 10628
rect 57195 10625 57207 10659
rect 57149 10619 57207 10625
rect 57333 10659 57391 10665
rect 57333 10625 57345 10659
rect 57379 10656 57391 10659
rect 57882 10656 57888 10668
rect 57379 10628 57888 10656
rect 57379 10625 57391 10628
rect 57333 10619 57391 10625
rect 57882 10616 57888 10628
rect 57940 10616 57946 10668
rect 38028 10560 38700 10588
rect 32732 10548 32738 10560
rect 27212 10492 28120 10520
rect 28276 10492 28580 10520
rect 31021 10523 31079 10529
rect 27212 10480 27218 10492
rect 11204 10424 12020 10452
rect 11204 10412 11210 10424
rect 14826 10412 14832 10464
rect 14884 10412 14890 10464
rect 16850 10412 16856 10464
rect 16908 10452 16914 10464
rect 17310 10452 17316 10464
rect 16908 10424 17316 10452
rect 16908 10412 16914 10424
rect 17310 10412 17316 10424
rect 17368 10412 17374 10464
rect 24118 10412 24124 10464
rect 24176 10452 24182 10464
rect 24578 10452 24584 10464
rect 24176 10424 24584 10452
rect 24176 10412 24182 10424
rect 24578 10412 24584 10424
rect 24636 10452 24642 10464
rect 25130 10452 25136 10464
rect 24636 10424 25136 10452
rect 24636 10412 24642 10424
rect 25130 10412 25136 10424
rect 25188 10412 25194 10464
rect 25406 10412 25412 10464
rect 25464 10452 25470 10464
rect 27982 10452 27988 10464
rect 25464 10424 27988 10452
rect 25464 10412 25470 10424
rect 27982 10412 27988 10424
rect 28040 10412 28046 10464
rect 28092 10452 28120 10492
rect 31021 10489 31033 10523
rect 31067 10520 31079 10523
rect 36538 10520 36544 10532
rect 31067 10492 36544 10520
rect 31067 10489 31079 10492
rect 31021 10483 31079 10489
rect 36538 10480 36544 10492
rect 36596 10480 36602 10532
rect 29546 10452 29552 10464
rect 28092 10424 29552 10452
rect 29546 10412 29552 10424
rect 29604 10452 29610 10464
rect 29917 10455 29975 10461
rect 29917 10452 29929 10455
rect 29604 10424 29929 10452
rect 29604 10412 29610 10424
rect 29917 10421 29929 10424
rect 29963 10421 29975 10455
rect 29917 10415 29975 10421
rect 31754 10412 31760 10464
rect 31812 10452 31818 10464
rect 32306 10452 32312 10464
rect 31812 10424 32312 10452
rect 31812 10412 31818 10424
rect 32306 10412 32312 10424
rect 32364 10452 32370 10464
rect 35158 10452 35164 10464
rect 32364 10424 35164 10452
rect 32364 10412 32370 10424
rect 35158 10412 35164 10424
rect 35216 10412 35222 10464
rect 35526 10412 35532 10464
rect 35584 10412 35590 10464
rect 35710 10412 35716 10464
rect 35768 10412 35774 10464
rect 38010 10412 38016 10464
rect 38068 10452 38074 10464
rect 38565 10455 38623 10461
rect 38565 10452 38577 10455
rect 38068 10424 38577 10452
rect 38068 10412 38074 10424
rect 38565 10421 38577 10424
rect 38611 10421 38623 10455
rect 38672 10452 38700 10560
rect 40034 10548 40040 10600
rect 40092 10588 40098 10600
rect 40678 10588 40684 10600
rect 40092 10560 40684 10588
rect 40092 10548 40098 10560
rect 40678 10548 40684 10560
rect 40736 10548 40742 10600
rect 41598 10452 41604 10464
rect 38672 10424 41604 10452
rect 38565 10415 38623 10421
rect 41598 10412 41604 10424
rect 41656 10412 41662 10464
rect 41782 10412 41788 10464
rect 41840 10452 41846 10464
rect 42061 10455 42119 10461
rect 42061 10452 42073 10455
rect 41840 10424 42073 10452
rect 41840 10412 41846 10424
rect 42061 10421 42073 10424
rect 42107 10421 42119 10455
rect 42061 10415 42119 10421
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 11422 10208 11428 10260
rect 11480 10248 11486 10260
rect 11517 10251 11575 10257
rect 11517 10248 11529 10251
rect 11480 10220 11529 10248
rect 11480 10208 11486 10220
rect 11517 10217 11529 10220
rect 11563 10217 11575 10251
rect 11517 10211 11575 10217
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 15378 10248 15384 10260
rect 14056 10220 15384 10248
rect 14056 10208 14062 10220
rect 15378 10208 15384 10220
rect 15436 10248 15442 10260
rect 16390 10248 16396 10260
rect 15436 10220 16396 10248
rect 15436 10208 15442 10220
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 16482 10208 16488 10260
rect 16540 10248 16546 10260
rect 16540 10220 17172 10248
rect 16540 10208 16546 10220
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 11333 10183 11391 10189
rect 11333 10180 11345 10183
rect 8536 10152 11345 10180
rect 8536 10140 8542 10152
rect 11333 10149 11345 10152
rect 11379 10149 11391 10183
rect 11333 10143 11391 10149
rect 12897 10183 12955 10189
rect 12897 10149 12909 10183
rect 12943 10180 12955 10183
rect 13170 10180 13176 10192
rect 12943 10152 13176 10180
rect 12943 10149 12955 10152
rect 12897 10143 12955 10149
rect 13170 10140 13176 10152
rect 13228 10140 13234 10192
rect 14734 10140 14740 10192
rect 14792 10180 14798 10192
rect 16666 10180 16672 10192
rect 14792 10152 16672 10180
rect 14792 10140 14798 10152
rect 16666 10140 16672 10152
rect 16724 10140 16730 10192
rect 16945 10183 17003 10189
rect 16945 10149 16957 10183
rect 16991 10180 17003 10183
rect 17034 10180 17040 10192
rect 16991 10152 17040 10180
rect 16991 10149 17003 10152
rect 16945 10143 17003 10149
rect 17034 10140 17040 10152
rect 17092 10140 17098 10192
rect 17144 10180 17172 10220
rect 18782 10208 18788 10260
rect 18840 10248 18846 10260
rect 19150 10248 19156 10260
rect 18840 10220 19156 10248
rect 18840 10208 18846 10220
rect 19150 10208 19156 10220
rect 19208 10248 19214 10260
rect 24486 10248 24492 10260
rect 19208 10220 24492 10248
rect 19208 10208 19214 10220
rect 24486 10208 24492 10220
rect 24544 10208 24550 10260
rect 31846 10248 31852 10260
rect 27908 10220 31852 10248
rect 19058 10180 19064 10192
rect 17144 10152 19064 10180
rect 19058 10140 19064 10152
rect 19116 10140 19122 10192
rect 21082 10180 21088 10192
rect 20824 10152 21088 10180
rect 934 10072 940 10124
rect 992 10112 998 10124
rect 1765 10115 1823 10121
rect 1765 10112 1777 10115
rect 992 10084 1777 10112
rect 992 10072 998 10084
rect 1765 10081 1777 10084
rect 1811 10081 1823 10115
rect 17218 10112 17224 10124
rect 1765 10075 1823 10081
rect 2746 10084 17224 10112
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 2746 10044 2774 10084
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 18325 10115 18383 10121
rect 18325 10081 18337 10115
rect 18371 10112 18383 10115
rect 18506 10112 18512 10124
rect 18371 10084 18512 10112
rect 18371 10081 18383 10084
rect 18325 10075 18383 10081
rect 18506 10072 18512 10084
rect 18564 10072 18570 10124
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19797 10115 19855 10121
rect 19797 10112 19809 10115
rect 19484 10084 19809 10112
rect 19484 10072 19490 10084
rect 19797 10081 19809 10084
rect 19843 10081 19855 10115
rect 19797 10075 19855 10081
rect 1627 10016 2774 10044
rect 11057 10047 11115 10053
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 11057 10013 11069 10047
rect 11103 10044 11115 10047
rect 11330 10044 11336 10056
rect 11103 10016 11336 10044
rect 11103 10013 11115 10016
rect 11057 10007 11115 10013
rect 11330 10004 11336 10016
rect 11388 10044 11394 10056
rect 11698 10044 11704 10056
rect 11388 10016 11704 10044
rect 11388 10004 11394 10016
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 12802 10004 12808 10056
rect 12860 10004 12866 10056
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10044 13139 10047
rect 13446 10044 13452 10056
rect 13127 10016 13452 10044
rect 13127 10013 13139 10016
rect 13081 10007 13139 10013
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 14369 10047 14427 10053
rect 14369 10013 14381 10047
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 1946 9868 1952 9920
rect 2004 9908 2010 9920
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 2004 9880 13277 9908
rect 2004 9868 2010 9880
rect 13265 9877 13277 9880
rect 13311 9877 13323 9911
rect 14384 9908 14412 10007
rect 14826 10004 14832 10056
rect 14884 10044 14890 10056
rect 15841 10047 15899 10053
rect 14884 10016 15516 10044
rect 14884 10004 14890 10016
rect 15488 9988 15516 10016
rect 15841 10013 15853 10047
rect 15887 10044 15899 10047
rect 16114 10044 16120 10056
rect 15887 10016 16120 10044
rect 15887 10013 15899 10016
rect 15841 10007 15899 10013
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 14458 9936 14464 9988
rect 14516 9976 14522 9988
rect 14921 9979 14979 9985
rect 14921 9976 14933 9979
rect 14516 9948 14933 9976
rect 14516 9936 14522 9948
rect 14921 9945 14933 9948
rect 14967 9976 14979 9979
rect 14967 9948 15424 9976
rect 14967 9945 14979 9948
rect 14921 9939 14979 9945
rect 15194 9908 15200 9920
rect 14384 9880 15200 9908
rect 13265 9871 13323 9877
rect 15194 9868 15200 9880
rect 15252 9868 15258 9920
rect 15396 9908 15424 9948
rect 15470 9936 15476 9988
rect 15528 9976 15534 9988
rect 16316 9976 16344 10007
rect 16390 10004 16396 10056
rect 16448 10004 16454 10056
rect 16666 10004 16672 10056
rect 16724 10044 16730 10056
rect 16761 10047 16819 10053
rect 16761 10044 16773 10047
rect 16724 10016 16773 10044
rect 16724 10004 16730 10016
rect 16761 10013 16773 10016
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 17678 10004 17684 10056
rect 17736 10004 17742 10056
rect 20064 10047 20122 10053
rect 20064 10013 20076 10047
rect 20110 10044 20122 10047
rect 20530 10044 20536 10056
rect 20110 10016 20536 10044
rect 20110 10013 20122 10016
rect 20064 10007 20122 10013
rect 20530 10004 20536 10016
rect 20588 10004 20594 10056
rect 17402 9976 17408 9988
rect 15528 9948 17408 9976
rect 15528 9936 15534 9948
rect 17402 9936 17408 9948
rect 17460 9936 17466 9988
rect 18966 9936 18972 9988
rect 19024 9976 19030 9988
rect 20824 9976 20852 10152
rect 21082 10140 21088 10152
rect 21140 10180 21146 10192
rect 21177 10183 21235 10189
rect 21177 10180 21189 10183
rect 21140 10152 21189 10180
rect 21140 10140 21146 10152
rect 21177 10149 21189 10152
rect 21223 10149 21235 10183
rect 21177 10143 21235 10149
rect 21266 10140 21272 10192
rect 21324 10180 21330 10192
rect 21818 10180 21824 10192
rect 21324 10152 21824 10180
rect 21324 10140 21330 10152
rect 21818 10140 21824 10152
rect 21876 10180 21882 10192
rect 24762 10189 24768 10192
rect 24746 10183 24768 10189
rect 21876 10152 22094 10180
rect 21876 10140 21882 10152
rect 22066 10112 22094 10152
rect 24746 10149 24758 10183
rect 24746 10143 24768 10149
rect 24762 10140 24768 10143
rect 24820 10140 24826 10192
rect 24854 10140 24860 10192
rect 24912 10140 24918 10192
rect 27706 10140 27712 10192
rect 27764 10140 27770 10192
rect 22189 10115 22247 10121
rect 22189 10112 22201 10115
rect 22066 10084 22201 10112
rect 22189 10081 22201 10084
rect 22235 10081 22247 10115
rect 22189 10075 22247 10081
rect 23566 10072 23572 10124
rect 23624 10112 23630 10124
rect 23661 10115 23719 10121
rect 23661 10112 23673 10115
rect 23624 10084 23673 10112
rect 23624 10072 23630 10084
rect 23661 10081 23673 10084
rect 23707 10081 23719 10115
rect 23661 10075 23719 10081
rect 24949 10115 25007 10121
rect 24949 10081 24961 10115
rect 24995 10112 25007 10115
rect 25038 10112 25044 10124
rect 24995 10084 25044 10112
rect 24995 10081 25007 10084
rect 24949 10075 25007 10081
rect 25038 10072 25044 10084
rect 25096 10072 25102 10124
rect 25130 10072 25136 10124
rect 25188 10112 25194 10124
rect 25777 10115 25835 10121
rect 25777 10112 25789 10115
rect 25188 10084 25789 10112
rect 25188 10072 25194 10084
rect 25777 10081 25789 10084
rect 25823 10081 25835 10115
rect 25777 10075 25835 10081
rect 26160 10084 27660 10112
rect 26160 10056 26188 10084
rect 21082 10004 21088 10056
rect 21140 10044 21146 10056
rect 22097 10047 22155 10053
rect 22097 10044 22109 10047
rect 21140 10016 22109 10044
rect 21140 10004 21146 10016
rect 22097 10013 22109 10016
rect 22143 10013 22155 10047
rect 22097 10007 22155 10013
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10044 23903 10047
rect 23891 10016 24532 10044
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 19024 9948 20852 9976
rect 19024 9936 19030 9948
rect 20898 9936 20904 9988
rect 20956 9976 20962 9988
rect 24029 9979 24087 9985
rect 24029 9976 24041 9979
rect 20956 9948 24041 9976
rect 20956 9936 20962 9948
rect 24029 9945 24041 9948
rect 24075 9945 24087 9979
rect 24029 9939 24087 9945
rect 16482 9908 16488 9920
rect 15396 9880 16488 9908
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 16850 9908 16856 9920
rect 16632 9880 16856 9908
rect 16632 9868 16638 9880
rect 16850 9868 16856 9880
rect 16908 9868 16914 9920
rect 19058 9868 19064 9920
rect 19116 9908 19122 9920
rect 21450 9908 21456 9920
rect 19116 9880 21456 9908
rect 19116 9868 19122 9880
rect 21450 9868 21456 9880
rect 21508 9868 21514 9920
rect 21634 9868 21640 9920
rect 21692 9868 21698 9920
rect 22005 9911 22063 9917
rect 22005 9877 22017 9911
rect 22051 9908 22063 9911
rect 22462 9908 22468 9920
rect 22051 9880 22468 9908
rect 22051 9877 22063 9880
rect 22005 9871 22063 9877
rect 22462 9868 22468 9880
rect 22520 9868 22526 9920
rect 24504 9908 24532 10016
rect 24854 10004 24860 10056
rect 24912 10044 24918 10056
rect 25317 10047 25375 10053
rect 25317 10044 25329 10047
rect 24912 10016 25329 10044
rect 24912 10004 24918 10016
rect 25317 10013 25329 10016
rect 25363 10044 25375 10047
rect 25406 10044 25412 10056
rect 25363 10016 25412 10044
rect 25363 10013 25375 10016
rect 25317 10007 25375 10013
rect 25406 10004 25412 10016
rect 25464 10004 25470 10056
rect 25700 10016 26004 10044
rect 24581 9979 24639 9985
rect 24581 9945 24593 9979
rect 24627 9976 24639 9979
rect 25700 9976 25728 10016
rect 24627 9948 25728 9976
rect 25976 9976 26004 10016
rect 26050 10004 26056 10056
rect 26108 10004 26114 10056
rect 26142 10004 26148 10056
rect 26200 10004 26206 10056
rect 26329 10047 26387 10053
rect 26329 10013 26341 10047
rect 26375 10013 26387 10047
rect 26329 10007 26387 10013
rect 26344 9976 26372 10007
rect 26510 10004 26516 10056
rect 26568 10004 26574 10056
rect 26789 10047 26847 10053
rect 26789 10013 26801 10047
rect 26835 10044 26847 10047
rect 27338 10044 27344 10056
rect 26835 10016 27344 10044
rect 26835 10013 26847 10016
rect 26789 10007 26847 10013
rect 27338 10004 27344 10016
rect 27396 10004 27402 10056
rect 27522 9976 27528 9988
rect 25976 9948 27528 9976
rect 24627 9945 24639 9948
rect 24581 9939 24639 9945
rect 27522 9936 27528 9948
rect 27580 9936 27586 9988
rect 27632 9976 27660 10084
rect 27908 10053 27936 10220
rect 31846 10208 31852 10220
rect 31904 10208 31910 10260
rect 31941 10251 31999 10257
rect 31941 10217 31953 10251
rect 31987 10248 31999 10251
rect 33594 10248 33600 10260
rect 31987 10220 33600 10248
rect 31987 10217 31999 10220
rect 31941 10211 31999 10217
rect 33594 10208 33600 10220
rect 33652 10208 33658 10260
rect 34238 10208 34244 10260
rect 34296 10248 34302 10260
rect 36078 10248 36084 10260
rect 34296 10220 36084 10248
rect 34296 10208 34302 10220
rect 36078 10208 36084 10220
rect 36136 10208 36142 10260
rect 36188 10220 39896 10248
rect 34422 10180 34428 10192
rect 28000 10152 34428 10180
rect 28000 10053 28028 10152
rect 34422 10140 34428 10152
rect 34480 10140 34486 10192
rect 28258 10072 28264 10124
rect 28316 10072 28322 10124
rect 29730 10072 29736 10124
rect 29788 10072 29794 10124
rect 30742 10112 30748 10124
rect 29932 10084 30748 10112
rect 27893 10047 27951 10053
rect 27893 10013 27905 10047
rect 27939 10013 27951 10047
rect 28000 10047 28063 10053
rect 28000 10016 28017 10047
rect 27893 10007 27951 10013
rect 28005 10013 28017 10016
rect 28051 10013 28063 10047
rect 28005 10007 28063 10013
rect 28117 10047 28175 10053
rect 28117 10013 28129 10047
rect 28163 10044 28175 10047
rect 28276 10044 28304 10072
rect 28163 10016 28304 10044
rect 28721 10047 28779 10053
rect 28163 10013 28175 10016
rect 28117 10007 28175 10013
rect 28721 10013 28733 10047
rect 28767 10044 28779 10047
rect 29454 10044 29460 10056
rect 28767 10016 29460 10044
rect 28767 10013 28779 10016
rect 28721 10007 28779 10013
rect 29454 10004 29460 10016
rect 29512 10004 29518 10056
rect 29932 9988 29960 10084
rect 30742 10072 30748 10084
rect 30800 10072 30806 10124
rect 36188 10112 36216 10220
rect 38194 10180 38200 10192
rect 37660 10152 38200 10180
rect 37660 10121 37688 10152
rect 38194 10140 38200 10152
rect 38252 10140 38258 10192
rect 32048 10084 36216 10112
rect 37645 10115 37703 10121
rect 32048 10044 32076 10084
rect 37645 10081 37657 10115
rect 37691 10081 37703 10115
rect 39298 10112 39304 10124
rect 37645 10075 37703 10081
rect 38212 10084 39304 10112
rect 30024 10016 32076 10044
rect 28261 9979 28319 9985
rect 28261 9976 28273 9979
rect 27632 9948 28273 9976
rect 28261 9945 28273 9948
rect 28307 9945 28319 9979
rect 28261 9939 28319 9945
rect 28994 9936 29000 9988
rect 29052 9936 29058 9988
rect 29914 9936 29920 9988
rect 29972 9936 29978 9988
rect 25498 9908 25504 9920
rect 24504 9880 25504 9908
rect 25498 9868 25504 9880
rect 25556 9868 25562 9920
rect 26878 9868 26884 9920
rect 26936 9908 26942 9920
rect 27062 9908 27068 9920
rect 26936 9880 27068 9908
rect 26936 9868 26942 9880
rect 27062 9868 27068 9880
rect 27120 9908 27126 9920
rect 27157 9911 27215 9917
rect 27157 9908 27169 9911
rect 27120 9880 27169 9908
rect 27120 9868 27126 9880
rect 27157 9877 27169 9880
rect 27203 9877 27215 9911
rect 27157 9871 27215 9877
rect 28350 9868 28356 9920
rect 28408 9908 28414 9920
rect 28902 9908 28908 9920
rect 28408 9880 28908 9908
rect 28408 9868 28414 9880
rect 28902 9868 28908 9880
rect 28960 9868 28966 9920
rect 30024 9917 30052 10016
rect 32122 10004 32128 10056
rect 32180 10004 32186 10056
rect 32398 10004 32404 10056
rect 32456 10004 32462 10056
rect 33594 10004 33600 10056
rect 33652 10044 33658 10056
rect 33870 10044 33876 10056
rect 33652 10016 33876 10044
rect 33652 10004 33658 10016
rect 33870 10004 33876 10016
rect 33928 10004 33934 10056
rect 35069 10047 35127 10053
rect 35069 10013 35081 10047
rect 35115 10044 35127 10047
rect 35710 10044 35716 10056
rect 35115 10016 35716 10044
rect 35115 10013 35127 10016
rect 35069 10007 35127 10013
rect 35710 10004 35716 10016
rect 35768 10004 35774 10056
rect 35894 10004 35900 10056
rect 35952 10044 35958 10056
rect 37369 10047 37427 10053
rect 37369 10044 37381 10047
rect 35952 10016 37381 10044
rect 35952 10004 35958 10016
rect 37369 10013 37381 10016
rect 37415 10013 37427 10047
rect 37369 10007 37427 10013
rect 30282 9936 30288 9988
rect 30340 9936 30346 9988
rect 31846 9936 31852 9988
rect 31904 9976 31910 9988
rect 32490 9976 32496 9988
rect 31904 9948 32496 9976
rect 31904 9936 31910 9948
rect 32490 9936 32496 9948
rect 32548 9936 32554 9988
rect 30009 9911 30067 9917
rect 30009 9877 30021 9911
rect 30055 9877 30067 9911
rect 30009 9871 30067 9877
rect 30098 9868 30104 9920
rect 30156 9868 30162 9920
rect 30374 9868 30380 9920
rect 30432 9908 30438 9920
rect 30558 9908 30564 9920
rect 30432 9880 30564 9908
rect 30432 9868 30438 9880
rect 30558 9868 30564 9880
rect 30616 9868 30622 9920
rect 32306 9868 32312 9920
rect 32364 9868 32370 9920
rect 33888 9908 33916 10004
rect 35250 9936 35256 9988
rect 35308 9936 35314 9988
rect 35434 9936 35440 9988
rect 35492 9936 35498 9988
rect 37274 9908 37280 9920
rect 33888 9880 37280 9908
rect 37274 9868 37280 9880
rect 37332 9908 37338 9920
rect 38212 9908 38240 10084
rect 38286 10004 38292 10056
rect 38344 10004 38350 10056
rect 38580 10053 38608 10084
rect 39298 10072 39304 10084
rect 39356 10072 39362 10124
rect 39868 10112 39896 10220
rect 41322 10208 41328 10260
rect 41380 10208 41386 10260
rect 39942 10140 39948 10192
rect 40000 10180 40006 10192
rect 46382 10180 46388 10192
rect 40000 10152 46388 10180
rect 40000 10140 40006 10152
rect 41782 10112 41788 10124
rect 39868 10084 41788 10112
rect 41782 10072 41788 10084
rect 41840 10072 41846 10124
rect 41984 10121 42012 10152
rect 46382 10140 46388 10152
rect 46440 10140 46446 10192
rect 41969 10115 42027 10121
rect 41969 10081 41981 10115
rect 42015 10081 42027 10115
rect 41969 10075 42027 10081
rect 42334 10072 42340 10124
rect 42392 10112 42398 10124
rect 42702 10112 42708 10124
rect 42392 10084 42708 10112
rect 42392 10072 42398 10084
rect 42702 10072 42708 10084
rect 42760 10072 42766 10124
rect 45649 10115 45707 10121
rect 45649 10112 45661 10115
rect 44376 10084 45661 10112
rect 38427 10047 38485 10053
rect 38427 10013 38439 10047
rect 38473 10013 38485 10047
rect 38427 10007 38485 10013
rect 38565 10047 38623 10053
rect 38565 10013 38577 10047
rect 38611 10013 38623 10047
rect 38565 10007 38623 10013
rect 38754 10047 38812 10053
rect 38754 10013 38766 10047
rect 38800 10044 38812 10047
rect 38800 10016 38884 10044
rect 38800 10013 38812 10016
rect 38754 10007 38812 10013
rect 38452 9976 38480 10007
rect 38304 9948 38480 9976
rect 38304 9920 38332 9948
rect 38654 9936 38660 9988
rect 38712 9936 38718 9988
rect 38856 9976 38884 10016
rect 39114 9976 39120 9988
rect 38856 9948 39120 9976
rect 39114 9936 39120 9948
rect 39172 9936 39178 9988
rect 41693 9979 41751 9985
rect 41693 9945 41705 9979
rect 41739 9976 41751 9979
rect 41874 9976 41880 9988
rect 41739 9948 41880 9976
rect 41739 9945 41751 9948
rect 41693 9939 41751 9945
rect 41874 9936 41880 9948
rect 41932 9936 41938 9988
rect 42720 9976 42748 10072
rect 44174 10004 44180 10056
rect 44232 10004 44238 10056
rect 44266 10004 44272 10056
rect 44324 10004 44330 10056
rect 44376 10053 44404 10084
rect 45649 10081 45661 10084
rect 45695 10081 45707 10115
rect 46566 10112 46572 10124
rect 45649 10075 45707 10081
rect 45848 10084 46572 10112
rect 45848 10053 45876 10084
rect 46566 10072 46572 10084
rect 46624 10072 46630 10124
rect 58158 10072 58164 10124
rect 58216 10072 58222 10124
rect 44361 10047 44419 10053
rect 44361 10013 44373 10047
rect 44407 10013 44419 10047
rect 44361 10007 44419 10013
rect 44545 10047 44603 10053
rect 44545 10013 44557 10047
rect 44591 10013 44603 10047
rect 44545 10007 44603 10013
rect 45833 10047 45891 10053
rect 45833 10013 45845 10047
rect 45879 10013 45891 10047
rect 45833 10007 45891 10013
rect 44560 9976 44588 10007
rect 46106 10004 46112 10056
rect 46164 10004 46170 10056
rect 52362 10004 52368 10056
rect 52420 10044 52426 10056
rect 57885 10047 57943 10053
rect 57885 10044 57897 10047
rect 52420 10016 57897 10044
rect 52420 10004 52426 10016
rect 57885 10013 57897 10016
rect 57931 10013 57943 10047
rect 57885 10007 57943 10013
rect 42720 9948 44588 9976
rect 44818 9936 44824 9988
rect 44876 9976 44882 9988
rect 46845 9979 46903 9985
rect 46845 9976 46857 9979
rect 44876 9948 46857 9976
rect 44876 9936 44882 9948
rect 46845 9945 46857 9948
rect 46891 9945 46903 9979
rect 46845 9939 46903 9945
rect 55306 9936 55312 9988
rect 55364 9976 55370 9988
rect 57057 9979 57115 9985
rect 55364 9948 57008 9976
rect 55364 9936 55370 9948
rect 37332 9880 38240 9908
rect 37332 9868 37338 9880
rect 38286 9868 38292 9920
rect 38344 9868 38350 9920
rect 38378 9868 38384 9920
rect 38436 9908 38442 9920
rect 38933 9911 38991 9917
rect 38933 9908 38945 9911
rect 38436 9880 38945 9908
rect 38436 9868 38442 9880
rect 38933 9877 38945 9880
rect 38979 9877 38991 9911
rect 38933 9871 38991 9877
rect 43901 9911 43959 9917
rect 43901 9877 43913 9911
rect 43947 9908 43959 9911
rect 45462 9908 45468 9920
rect 43947 9880 45468 9908
rect 43947 9877 43959 9880
rect 43901 9871 43959 9877
rect 45462 9868 45468 9880
rect 45520 9868 45526 9920
rect 46017 9911 46075 9917
rect 46017 9877 46029 9911
rect 46063 9908 46075 9911
rect 46290 9908 46296 9920
rect 46063 9880 46296 9908
rect 46063 9877 46075 9880
rect 46017 9871 46075 9877
rect 46290 9868 46296 9880
rect 46348 9868 46354 9920
rect 46934 9868 46940 9920
rect 46992 9908 46998 9920
rect 48133 9911 48191 9917
rect 48133 9908 48145 9911
rect 46992 9880 48145 9908
rect 46992 9868 46998 9880
rect 48133 9877 48145 9880
rect 48179 9908 48191 9911
rect 56870 9908 56876 9920
rect 48179 9880 56876 9908
rect 48179 9877 48191 9880
rect 48133 9871 48191 9877
rect 56870 9868 56876 9880
rect 56928 9868 56934 9920
rect 56980 9908 57008 9948
rect 57057 9945 57069 9979
rect 57103 9976 57115 9979
rect 58986 9976 58992 9988
rect 57103 9948 58992 9976
rect 57103 9945 57115 9948
rect 57057 9939 57115 9945
rect 58986 9936 58992 9948
rect 59044 9936 59050 9988
rect 57149 9911 57207 9917
rect 57149 9908 57161 9911
rect 56980 9880 57161 9908
rect 57149 9877 57161 9880
rect 57195 9877 57207 9911
rect 57149 9871 57207 9877
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 22002 9704 22008 9716
rect 16592 9676 22008 9704
rect 15930 9636 15936 9648
rect 15580 9608 15936 9636
rect 1581 9571 1639 9577
rect 1581 9537 1593 9571
rect 1627 9568 1639 9571
rect 4062 9568 4068 9580
rect 1627 9540 4068 9568
rect 1627 9537 1639 9540
rect 1581 9531 1639 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 13357 9571 13415 9577
rect 13357 9568 13369 9571
rect 12860 9540 13369 9568
rect 12860 9528 12866 9540
rect 13357 9537 13369 9540
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 13446 9528 13452 9580
rect 13504 9528 13510 9580
rect 13633 9571 13691 9577
rect 13633 9537 13645 9571
rect 13679 9537 13691 9571
rect 13633 9531 13691 9537
rect 13725 9571 13783 9577
rect 13725 9537 13737 9571
rect 13771 9568 13783 9571
rect 14458 9568 14464 9580
rect 13771 9540 14464 9568
rect 13771 9537 13783 9540
rect 13725 9531 13783 9537
rect 934 9460 940 9512
rect 992 9500 998 9512
rect 1765 9503 1823 9509
rect 1765 9500 1777 9503
rect 992 9472 1777 9500
rect 992 9460 998 9472
rect 1765 9469 1777 9472
rect 1811 9469 1823 9503
rect 1765 9463 1823 9469
rect 8754 9460 8760 9512
rect 8812 9460 8818 9512
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9674 9500 9680 9512
rect 9263 9472 9680 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 11054 9460 11060 9512
rect 11112 9500 11118 9512
rect 12342 9500 12348 9512
rect 11112 9472 12348 9500
rect 11112 9460 11118 9472
rect 12342 9460 12348 9472
rect 12400 9500 12406 9512
rect 13648 9500 13676 9531
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 15197 9571 15255 9577
rect 15197 9537 15209 9571
rect 15243 9537 15255 9571
rect 15197 9531 15255 9537
rect 12400 9472 13676 9500
rect 12400 9460 12406 9472
rect 7190 9392 7196 9444
rect 7248 9432 7254 9444
rect 9033 9435 9091 9441
rect 9033 9432 9045 9435
rect 7248 9404 9045 9432
rect 7248 9392 7254 9404
rect 9033 9401 9045 9404
rect 9079 9401 9091 9435
rect 9033 9395 9091 9401
rect 10778 9392 10784 9444
rect 10836 9432 10842 9444
rect 10836 9404 14872 9432
rect 10836 9392 10842 9404
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 13173 9367 13231 9373
rect 13173 9364 13185 9367
rect 11020 9336 13185 9364
rect 11020 9324 11026 9336
rect 13173 9333 13185 9336
rect 13219 9364 13231 9367
rect 14366 9364 14372 9376
rect 13219 9336 14372 9364
rect 13219 9333 13231 9336
rect 13173 9327 13231 9333
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 14844 9373 14872 9404
rect 14918 9392 14924 9444
rect 14976 9432 14982 9444
rect 15212 9432 15240 9531
rect 15470 9528 15476 9580
rect 15528 9528 15534 9580
rect 15580 9577 15608 9608
rect 15930 9596 15936 9608
rect 15988 9636 15994 9648
rect 16592 9636 16620 9676
rect 22002 9664 22008 9676
rect 22060 9664 22066 9716
rect 22830 9664 22836 9716
rect 22888 9704 22894 9716
rect 22888 9676 27476 9704
rect 22888 9664 22894 9676
rect 20064 9639 20122 9645
rect 15988 9608 16620 9636
rect 17052 9608 18828 9636
rect 15988 9596 15994 9608
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 15838 9528 15844 9580
rect 15896 9528 15902 9580
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9537 16175 9571
rect 16117 9531 16175 9537
rect 16132 9500 16160 9531
rect 16206 9528 16212 9580
rect 16264 9568 16270 9580
rect 17052 9577 17080 9608
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 16264 9540 17049 9568
rect 16264 9528 16270 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 18322 9528 18328 9580
rect 18380 9568 18386 9580
rect 18693 9571 18751 9577
rect 18693 9568 18705 9571
rect 18380 9540 18705 9568
rect 18380 9528 18386 9540
rect 18693 9537 18705 9540
rect 18739 9537 18751 9571
rect 18800 9568 18828 9608
rect 20064 9605 20076 9639
rect 20110 9636 20122 9639
rect 21634 9636 21640 9648
rect 20110 9608 21640 9636
rect 20110 9605 20122 9608
rect 20064 9599 20122 9605
rect 21634 9596 21640 9608
rect 21692 9596 21698 9648
rect 21744 9608 23888 9636
rect 20438 9568 20444 9580
rect 18800 9540 20444 9568
rect 18693 9531 18751 9537
rect 20438 9528 20444 9540
rect 20496 9528 20502 9580
rect 17310 9500 17316 9512
rect 16132 9472 17316 9500
rect 17310 9460 17316 9472
rect 17368 9500 17374 9512
rect 17770 9500 17776 9512
rect 17368 9472 17776 9500
rect 17368 9460 17374 9472
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 19426 9460 19432 9512
rect 19484 9500 19490 9512
rect 19797 9503 19855 9509
rect 19797 9500 19809 9503
rect 19484 9472 19809 9500
rect 19484 9460 19490 9472
rect 19797 9469 19809 9472
rect 19843 9469 19855 9503
rect 19797 9463 19855 9469
rect 15562 9432 15568 9444
rect 14976 9404 15568 9432
rect 14976 9392 14982 9404
rect 15562 9392 15568 9404
rect 15620 9432 15626 9444
rect 18785 9435 18843 9441
rect 18785 9432 18797 9435
rect 15620 9404 18797 9432
rect 15620 9392 15626 9404
rect 18785 9401 18797 9404
rect 18831 9401 18843 9435
rect 21744 9432 21772 9608
rect 21818 9528 21824 9580
rect 21876 9568 21882 9580
rect 23382 9568 23388 9580
rect 21876 9540 23388 9568
rect 21876 9528 21882 9540
rect 23382 9528 23388 9540
rect 23440 9528 23446 9580
rect 23860 9500 23888 9608
rect 24210 9596 24216 9648
rect 24268 9636 24274 9648
rect 24673 9639 24731 9645
rect 24673 9636 24685 9639
rect 24268 9608 24685 9636
rect 24268 9596 24274 9608
rect 24673 9605 24685 9608
rect 24719 9605 24731 9639
rect 25498 9636 25504 9648
rect 24673 9599 24731 9605
rect 25332 9608 25504 9636
rect 23937 9571 23995 9577
rect 23937 9537 23949 9571
rect 23983 9568 23995 9571
rect 24578 9568 24584 9580
rect 23983 9540 24584 9568
rect 23983 9537 23995 9540
rect 23937 9531 23995 9537
rect 24578 9528 24584 9540
rect 24636 9528 24642 9580
rect 25332 9577 25360 9608
rect 25498 9596 25504 9608
rect 25556 9636 25562 9648
rect 25958 9636 25964 9648
rect 25556 9608 25964 9636
rect 25556 9596 25562 9608
rect 25958 9596 25964 9608
rect 26016 9596 26022 9648
rect 26050 9596 26056 9648
rect 26108 9636 26114 9648
rect 27448 9636 27476 9676
rect 27522 9664 27528 9716
rect 27580 9664 27586 9716
rect 28166 9704 28172 9716
rect 27632 9676 28172 9704
rect 27632 9636 27660 9676
rect 28166 9664 28172 9676
rect 28224 9664 28230 9716
rect 28813 9707 28871 9713
rect 28813 9673 28825 9707
rect 28859 9704 28871 9707
rect 29825 9707 29883 9713
rect 29825 9704 29837 9707
rect 28859 9676 29837 9704
rect 28859 9673 28871 9676
rect 28813 9667 28871 9673
rect 29825 9673 29837 9676
rect 29871 9704 29883 9707
rect 30098 9704 30104 9716
rect 29871 9676 30104 9704
rect 29871 9673 29883 9676
rect 29825 9667 29883 9673
rect 30098 9664 30104 9676
rect 30156 9664 30162 9716
rect 30374 9664 30380 9716
rect 30432 9704 30438 9716
rect 32030 9704 32036 9716
rect 30432 9676 32036 9704
rect 30432 9664 30438 9676
rect 32030 9664 32036 9676
rect 32088 9664 32094 9716
rect 32122 9664 32128 9716
rect 32180 9704 32186 9716
rect 32493 9707 32551 9713
rect 32493 9704 32505 9707
rect 32180 9676 32505 9704
rect 32180 9664 32186 9676
rect 32493 9673 32505 9676
rect 32539 9673 32551 9707
rect 32493 9667 32551 9673
rect 33134 9664 33140 9716
rect 33192 9704 33198 9716
rect 33192 9676 33272 9704
rect 33192 9664 33198 9676
rect 26108 9608 27200 9636
rect 27448 9608 27660 9636
rect 26108 9596 26114 9608
rect 25225 9571 25283 9577
rect 25225 9537 25237 9571
rect 25271 9537 25283 9571
rect 25225 9531 25283 9537
rect 25317 9571 25375 9577
rect 25317 9537 25329 9571
rect 25363 9537 25375 9571
rect 25317 9531 25375 9537
rect 25593 9571 25651 9577
rect 25593 9537 25605 9571
rect 25639 9568 25651 9571
rect 26694 9568 26700 9580
rect 25639 9540 26700 9568
rect 25639 9537 25651 9540
rect 25593 9531 25651 9537
rect 25240 9500 25268 9531
rect 26694 9528 26700 9540
rect 26752 9528 26758 9580
rect 27172 9577 27200 9608
rect 27706 9596 27712 9648
rect 27764 9636 27770 9648
rect 28442 9636 28448 9648
rect 27764 9608 28448 9636
rect 27764 9596 27770 9608
rect 28442 9596 28448 9608
rect 28500 9596 28506 9648
rect 28731 9639 28789 9645
rect 28731 9605 28743 9639
rect 28777 9636 28789 9639
rect 28777 9608 29132 9636
rect 28777 9605 28789 9608
rect 28731 9599 28789 9605
rect 27157 9571 27215 9577
rect 27157 9537 27169 9571
rect 27203 9568 27215 9571
rect 28166 9568 28172 9580
rect 27203 9540 28172 9568
rect 27203 9537 27215 9540
rect 27157 9531 27215 9537
rect 28166 9528 28172 9540
rect 28224 9568 28230 9580
rect 28629 9571 28687 9577
rect 28224 9540 28580 9568
rect 28224 9528 28230 9540
rect 25406 9500 25412 9512
rect 23860 9472 24348 9500
rect 25240 9472 25412 9500
rect 18785 9395 18843 9401
rect 20732 9404 21772 9432
rect 14829 9367 14887 9373
rect 14829 9333 14841 9367
rect 14875 9364 14887 9367
rect 18506 9364 18512 9376
rect 14875 9336 18512 9364
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 18874 9324 18880 9376
rect 18932 9364 18938 9376
rect 20732 9364 20760 9404
rect 24026 9392 24032 9444
rect 24084 9432 24090 9444
rect 24121 9435 24179 9441
rect 24121 9432 24133 9435
rect 24084 9404 24133 9432
rect 24084 9392 24090 9404
rect 24121 9401 24133 9404
rect 24167 9401 24179 9435
rect 24320 9432 24348 9472
rect 25406 9460 25412 9472
rect 25464 9460 25470 9512
rect 25774 9460 25780 9512
rect 25832 9460 25838 9512
rect 26050 9460 26056 9512
rect 26108 9460 26114 9512
rect 26786 9460 26792 9512
rect 26844 9500 26850 9512
rect 27249 9503 27307 9509
rect 27249 9500 27261 9503
rect 26844 9472 27261 9500
rect 26844 9460 26850 9472
rect 27249 9469 27261 9472
rect 27295 9469 27307 9503
rect 27249 9463 27307 9469
rect 24320 9404 27384 9432
rect 24121 9395 24179 9401
rect 18932 9336 20760 9364
rect 18932 9324 18938 9336
rect 21082 9324 21088 9376
rect 21140 9364 21146 9376
rect 21177 9367 21235 9373
rect 21177 9364 21189 9367
rect 21140 9336 21189 9364
rect 21140 9324 21146 9336
rect 21177 9333 21189 9336
rect 21223 9333 21235 9367
rect 21177 9327 21235 9333
rect 23658 9324 23664 9376
rect 23716 9364 23722 9376
rect 24854 9364 24860 9376
rect 23716 9336 24860 9364
rect 23716 9324 23722 9336
rect 24854 9324 24860 9336
rect 24912 9324 24918 9376
rect 25038 9324 25044 9376
rect 25096 9364 25102 9376
rect 26234 9364 26240 9376
rect 25096 9336 26240 9364
rect 25096 9324 25102 9336
rect 26234 9324 26240 9336
rect 26292 9324 26298 9376
rect 27356 9373 27384 9404
rect 28442 9392 28448 9444
rect 28500 9392 28506 9444
rect 28552 9432 28580 9540
rect 28629 9537 28641 9571
rect 28675 9537 28687 9571
rect 28629 9531 28687 9537
rect 28644 9500 28672 9531
rect 28902 9528 28908 9580
rect 28960 9568 28966 9580
rect 28997 9571 29055 9577
rect 28997 9568 29009 9571
rect 28960 9540 29009 9568
rect 28960 9528 28966 9540
rect 28997 9537 29009 9540
rect 29043 9537 29055 9571
rect 29104 9568 29132 9608
rect 29178 9596 29184 9648
rect 29236 9636 29242 9648
rect 29457 9639 29515 9645
rect 29457 9636 29469 9639
rect 29236 9608 29469 9636
rect 29236 9596 29242 9608
rect 29457 9605 29469 9608
rect 29503 9605 29515 9639
rect 33244 9636 33272 9676
rect 33318 9664 33324 9716
rect 33376 9704 33382 9716
rect 36446 9704 36452 9716
rect 33376 9676 36452 9704
rect 33376 9664 33382 9676
rect 36446 9664 36452 9676
rect 36504 9664 36510 9716
rect 36538 9664 36544 9716
rect 36596 9704 36602 9716
rect 44266 9704 44272 9716
rect 36596 9676 44272 9704
rect 36596 9664 36602 9676
rect 44266 9664 44272 9676
rect 44324 9664 44330 9716
rect 46566 9664 46572 9716
rect 46624 9664 46630 9716
rect 34330 9636 34336 9648
rect 29457 9599 29515 9605
rect 29564 9608 30236 9636
rect 29564 9568 29592 9608
rect 29104 9540 29592 9568
rect 29641 9571 29699 9577
rect 28997 9531 29055 9537
rect 29641 9537 29653 9571
rect 29687 9537 29699 9571
rect 29641 9531 29699 9537
rect 29779 9571 29837 9577
rect 29779 9537 29791 9571
rect 29825 9568 29837 9571
rect 29825 9540 29960 9568
rect 29825 9537 29837 9540
rect 29779 9531 29837 9537
rect 29178 9500 29184 9512
rect 28644 9472 29184 9500
rect 29178 9460 29184 9472
rect 29236 9500 29242 9512
rect 29656 9500 29684 9531
rect 29236 9472 29776 9500
rect 29236 9460 29242 9472
rect 29086 9432 29092 9444
rect 28552 9404 29092 9432
rect 29086 9392 29092 9404
rect 29144 9392 29150 9444
rect 27341 9367 27399 9373
rect 27341 9333 27353 9367
rect 27387 9364 27399 9367
rect 29270 9364 29276 9376
rect 27387 9336 29276 9364
rect 27387 9333 27399 9336
rect 27341 9327 27399 9333
rect 29270 9324 29276 9336
rect 29328 9324 29334 9376
rect 29748 9364 29776 9472
rect 29932 9432 29960 9540
rect 30006 9528 30012 9580
rect 30064 9528 30070 9580
rect 30208 9500 30236 9608
rect 33244 9608 34336 9636
rect 30282 9528 30288 9580
rect 30340 9568 30346 9580
rect 30929 9571 30987 9577
rect 30929 9568 30941 9571
rect 30340 9540 30941 9568
rect 30340 9528 30346 9540
rect 30929 9537 30941 9540
rect 30975 9537 30987 9571
rect 30929 9531 30987 9537
rect 31662 9528 31668 9580
rect 31720 9568 31726 9580
rect 31720 9540 32536 9568
rect 31720 9528 31726 9540
rect 31938 9500 31944 9512
rect 30208 9472 31944 9500
rect 31938 9460 31944 9472
rect 31996 9460 32002 9512
rect 32508 9500 32536 9540
rect 32582 9528 32588 9580
rect 32640 9528 32646 9580
rect 32766 9528 32772 9580
rect 32824 9528 32830 9580
rect 33244 9568 33272 9608
rect 34330 9596 34336 9608
rect 34388 9636 34394 9648
rect 38102 9636 38108 9648
rect 34388 9608 38108 9636
rect 34388 9596 34394 9608
rect 38102 9596 38108 9608
rect 38160 9636 38166 9648
rect 38378 9636 38384 9648
rect 38160 9608 38384 9636
rect 38160 9596 38166 9608
rect 38378 9596 38384 9608
rect 38436 9636 38442 9648
rect 43717 9639 43775 9645
rect 43717 9636 43729 9639
rect 38436 9608 43729 9636
rect 38436 9596 38442 9608
rect 43717 9605 43729 9608
rect 43763 9636 43775 9639
rect 44450 9636 44456 9648
rect 43763 9608 44456 9636
rect 43763 9605 43775 9608
rect 43717 9599 43775 9605
rect 44450 9596 44456 9608
rect 44508 9596 44514 9648
rect 45462 9645 45468 9648
rect 45456 9636 45468 9645
rect 45423 9608 45468 9636
rect 45456 9599 45468 9608
rect 45462 9596 45468 9599
rect 45520 9596 45526 9648
rect 33321 9571 33379 9577
rect 33321 9568 33333 9571
rect 33244 9540 33333 9568
rect 33321 9537 33333 9540
rect 33367 9537 33379 9571
rect 33321 9531 33379 9537
rect 33410 9528 33416 9580
rect 33468 9568 33474 9580
rect 35986 9568 35992 9580
rect 33468 9540 35992 9568
rect 33468 9528 33474 9540
rect 35986 9528 35992 9540
rect 36044 9528 36050 9580
rect 36170 9528 36176 9580
rect 36228 9528 36234 9580
rect 37642 9577 37648 9580
rect 37461 9571 37519 9577
rect 37461 9537 37473 9571
rect 37507 9537 37519 9571
rect 37461 9531 37519 9537
rect 37609 9571 37648 9577
rect 37609 9537 37621 9571
rect 37609 9531 37648 9537
rect 33505 9503 33563 9509
rect 33505 9500 33517 9503
rect 32508 9472 33517 9500
rect 33505 9469 33517 9472
rect 33551 9500 33563 9503
rect 34238 9500 34244 9512
rect 33551 9472 34244 9500
rect 33551 9469 33563 9472
rect 33505 9463 33563 9469
rect 34238 9460 34244 9472
rect 34296 9460 34302 9512
rect 36538 9432 36544 9444
rect 29932 9404 36544 9432
rect 36538 9392 36544 9404
rect 36596 9392 36602 9444
rect 37476 9432 37504 9531
rect 37642 9528 37648 9531
rect 37700 9528 37706 9580
rect 37734 9528 37740 9580
rect 37792 9528 37798 9580
rect 37829 9571 37887 9577
rect 37829 9537 37841 9571
rect 37875 9537 37887 9571
rect 37829 9531 37887 9537
rect 37844 9500 37872 9531
rect 37918 9528 37924 9580
rect 37976 9577 37982 9580
rect 37976 9568 37984 9577
rect 40497 9571 40555 9577
rect 37976 9540 38021 9568
rect 37976 9531 37984 9540
rect 40497 9537 40509 9571
rect 40543 9568 40555 9571
rect 41414 9568 41420 9580
rect 40543 9540 41420 9568
rect 40543 9537 40555 9540
rect 40497 9531 40555 9537
rect 37976 9528 37982 9531
rect 41414 9528 41420 9540
rect 41472 9528 41478 9580
rect 43898 9528 43904 9580
rect 43956 9528 43962 9580
rect 43990 9528 43996 9580
rect 44048 9528 44054 9580
rect 44085 9571 44143 9577
rect 44085 9537 44097 9571
rect 44131 9568 44143 9571
rect 45094 9568 45100 9580
rect 44131 9540 45100 9568
rect 44131 9537 44143 9540
rect 44085 9531 44143 9537
rect 45094 9528 45100 9540
rect 45152 9528 45158 9580
rect 45186 9528 45192 9580
rect 45244 9528 45250 9580
rect 56778 9528 56784 9580
rect 56836 9568 56842 9580
rect 57057 9571 57115 9577
rect 57057 9568 57069 9571
rect 56836 9540 57069 9568
rect 56836 9528 56842 9540
rect 57057 9537 57069 9540
rect 57103 9537 57115 9571
rect 57057 9531 57115 9537
rect 57238 9528 57244 9580
rect 57296 9528 57302 9580
rect 37844 9472 43852 9500
rect 37734 9432 37740 9444
rect 37476 9404 37740 9432
rect 37734 9392 37740 9404
rect 37792 9392 37798 9444
rect 39390 9392 39396 9444
rect 39448 9432 39454 9444
rect 43824 9432 43852 9472
rect 39448 9404 41414 9432
rect 43824 9404 44404 9432
rect 39448 9392 39454 9404
rect 30282 9364 30288 9376
rect 29748 9336 30288 9364
rect 30282 9324 30288 9336
rect 30340 9324 30346 9376
rect 31205 9367 31263 9373
rect 31205 9333 31217 9367
rect 31251 9364 31263 9367
rect 31478 9364 31484 9376
rect 31251 9336 31484 9364
rect 31251 9333 31263 9336
rect 31205 9327 31263 9333
rect 31478 9324 31484 9336
rect 31536 9324 31542 9376
rect 32309 9367 32367 9373
rect 32309 9333 32321 9367
rect 32355 9364 32367 9367
rect 32950 9364 32956 9376
rect 32355 9336 32956 9364
rect 32355 9333 32367 9336
rect 32309 9327 32367 9333
rect 32950 9324 32956 9336
rect 33008 9364 33014 9376
rect 35894 9364 35900 9376
rect 33008 9336 35900 9364
rect 33008 9324 33014 9336
rect 35894 9324 35900 9336
rect 35952 9324 35958 9376
rect 35989 9367 36047 9373
rect 35989 9333 36001 9367
rect 36035 9364 36047 9367
rect 36262 9364 36268 9376
rect 36035 9336 36268 9364
rect 36035 9333 36047 9336
rect 35989 9327 36047 9333
rect 36262 9324 36268 9336
rect 36320 9324 36326 9376
rect 37550 9324 37556 9376
rect 37608 9364 37614 9376
rect 38105 9367 38163 9373
rect 38105 9364 38117 9367
rect 37608 9336 38117 9364
rect 37608 9324 37614 9336
rect 38105 9333 38117 9336
rect 38151 9333 38163 9367
rect 38105 9327 38163 9333
rect 40586 9324 40592 9376
rect 40644 9324 40650 9376
rect 41386 9364 41414 9404
rect 44269 9367 44327 9373
rect 44269 9364 44281 9367
rect 41386 9336 44281 9364
rect 44269 9333 44281 9336
rect 44315 9333 44327 9367
rect 44376 9364 44404 9404
rect 46198 9364 46204 9376
rect 44376 9336 46204 9364
rect 44269 9327 44327 9333
rect 46198 9324 46204 9336
rect 46256 9324 46262 9376
rect 46474 9324 46480 9376
rect 46532 9364 46538 9376
rect 47118 9364 47124 9376
rect 46532 9336 47124 9364
rect 46532 9324 46538 9336
rect 47118 9324 47124 9336
rect 47176 9324 47182 9376
rect 56318 9324 56324 9376
rect 56376 9364 56382 9376
rect 57149 9367 57207 9373
rect 57149 9364 57161 9367
rect 56376 9336 57161 9364
rect 56376 9324 56382 9336
rect 57149 9333 57161 9336
rect 57195 9333 57207 9367
rect 57149 9327 57207 9333
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 25958 9160 25964 9172
rect 2746 9132 25964 9160
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8956 1639 8959
rect 2746 8956 2774 9132
rect 25958 9120 25964 9132
rect 26016 9120 26022 9172
rect 27890 9120 27896 9172
rect 27948 9160 27954 9172
rect 28445 9163 28503 9169
rect 28445 9160 28457 9163
rect 27948 9132 28457 9160
rect 27948 9120 27954 9132
rect 28445 9129 28457 9132
rect 28491 9129 28503 9163
rect 33870 9160 33876 9172
rect 28445 9123 28503 9129
rect 28966 9132 33876 9160
rect 12986 9052 12992 9104
rect 13044 9092 13050 9104
rect 13081 9095 13139 9101
rect 13081 9092 13093 9095
rect 13044 9064 13093 9092
rect 13044 9052 13050 9064
rect 13081 9061 13093 9064
rect 13127 9061 13139 9095
rect 13081 9055 13139 9061
rect 13262 9052 13268 9104
rect 13320 9052 13326 9104
rect 14660 9064 15332 9092
rect 12342 8984 12348 9036
rect 12400 9024 12406 9036
rect 14660 9024 14688 9064
rect 12400 8996 14688 9024
rect 15304 9024 15332 9064
rect 15470 9052 15476 9104
rect 15528 9092 15534 9104
rect 16298 9092 16304 9104
rect 15528 9064 16304 9092
rect 15528 9052 15534 9064
rect 16298 9052 16304 9064
rect 16356 9052 16362 9104
rect 16945 9095 17003 9101
rect 16945 9061 16957 9095
rect 16991 9092 17003 9095
rect 17126 9092 17132 9104
rect 16991 9064 17132 9092
rect 16991 9061 17003 9064
rect 16945 9055 17003 9061
rect 17126 9052 17132 9064
rect 17184 9052 17190 9104
rect 18874 9092 18880 9104
rect 18064 9064 18880 9092
rect 18064 9033 18092 9064
rect 18874 9052 18880 9064
rect 18932 9052 18938 9104
rect 20714 9052 20720 9104
rect 20772 9092 20778 9104
rect 21545 9095 21603 9101
rect 21545 9092 21557 9095
rect 20772 9064 21557 9092
rect 20772 9052 20778 9064
rect 21545 9061 21557 9064
rect 21591 9061 21603 9095
rect 21545 9055 21603 9061
rect 21634 9052 21640 9104
rect 21692 9092 21698 9104
rect 21692 9064 24072 9092
rect 21692 9052 21698 9064
rect 18049 9027 18107 9033
rect 18049 9024 18061 9027
rect 15304 8996 18061 9024
rect 12400 8984 12406 8996
rect 1627 8928 2774 8956
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 13446 8916 13452 8968
rect 13504 8956 13510 8968
rect 13504 8928 15056 8956
rect 13504 8916 13510 8928
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1857 8891 1915 8897
rect 1857 8888 1869 8891
rect 992 8860 1869 8888
rect 992 8848 998 8860
rect 1857 8857 1869 8860
rect 1903 8857 1915 8891
rect 1857 8851 1915 8857
rect 12618 8848 12624 8900
rect 12676 8888 12682 8900
rect 12805 8891 12863 8897
rect 12805 8888 12817 8891
rect 12676 8860 12817 8888
rect 12676 8848 12682 8860
rect 12805 8857 12817 8860
rect 12851 8857 12863 8891
rect 12805 8851 12863 8857
rect 14918 8848 14924 8900
rect 14976 8848 14982 8900
rect 14826 8780 14832 8832
rect 14884 8780 14890 8832
rect 15028 8829 15056 8928
rect 15304 8897 15332 8996
rect 18049 8993 18061 8996
rect 18095 8993 18107 9027
rect 18049 8987 18107 8993
rect 18506 8984 18512 9036
rect 18564 8984 18570 9036
rect 19426 8984 19432 9036
rect 19484 9024 19490 9036
rect 19521 9027 19579 9033
rect 19521 9024 19533 9027
rect 19484 8996 19533 9024
rect 19484 8984 19490 8996
rect 19521 8993 19533 8996
rect 19567 8993 19579 9027
rect 19521 8987 19579 8993
rect 16025 8959 16083 8965
rect 16025 8925 16037 8959
rect 16071 8956 16083 8959
rect 16298 8956 16304 8968
rect 16071 8928 16304 8956
rect 16071 8925 16083 8928
rect 16025 8919 16083 8925
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 16393 8959 16451 8965
rect 16393 8925 16405 8959
rect 16439 8925 16451 8959
rect 16393 8919 16451 8925
rect 15289 8891 15347 8897
rect 15289 8857 15301 8891
rect 15335 8857 15347 8891
rect 16408 8888 16436 8919
rect 16666 8916 16672 8968
rect 16724 8916 16730 8968
rect 17402 8916 17408 8968
rect 17460 8956 17466 8968
rect 17460 8928 18184 8956
rect 17460 8916 17466 8928
rect 16942 8888 16948 8900
rect 16408 8860 16948 8888
rect 15289 8851 15347 8857
rect 16942 8848 16948 8860
rect 17000 8888 17006 8900
rect 17310 8888 17316 8900
rect 17000 8860 17316 8888
rect 17000 8848 17006 8860
rect 17310 8848 17316 8860
rect 17368 8848 17374 8900
rect 17957 8891 18015 8897
rect 17957 8857 17969 8891
rect 18003 8857 18015 8891
rect 18156 8888 18184 8928
rect 18414 8916 18420 8968
rect 18472 8916 18478 8968
rect 18524 8956 18552 8984
rect 21361 8959 21419 8965
rect 18524 8928 20392 8956
rect 18509 8891 18567 8897
rect 18509 8888 18521 8891
rect 18156 8860 18521 8888
rect 17957 8851 18015 8857
rect 18509 8857 18521 8860
rect 18555 8857 18567 8891
rect 18509 8851 18567 8857
rect 18601 8891 18659 8897
rect 18601 8857 18613 8891
rect 18647 8857 18659 8891
rect 18601 8851 18659 8857
rect 19788 8891 19846 8897
rect 19788 8857 19800 8891
rect 19834 8888 19846 8891
rect 20254 8888 20260 8900
rect 19834 8860 20260 8888
rect 19834 8857 19846 8860
rect 19788 8851 19846 8857
rect 15013 8823 15071 8829
rect 15013 8789 15025 8823
rect 15059 8789 15071 8823
rect 15013 8783 15071 8789
rect 15102 8780 15108 8832
rect 15160 8780 15166 8832
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 17972 8820 18000 8851
rect 18322 8820 18328 8832
rect 16724 8792 18328 8820
rect 16724 8780 16730 8792
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 18414 8780 18420 8832
rect 18472 8820 18478 8832
rect 18616 8820 18644 8851
rect 20254 8848 20260 8860
rect 20312 8848 20318 8900
rect 20364 8888 20392 8928
rect 21361 8925 21373 8959
rect 21407 8956 21419 8959
rect 23934 8956 23940 8968
rect 21407 8928 23940 8956
rect 21407 8925 21419 8928
rect 21361 8919 21419 8925
rect 23934 8916 23940 8928
rect 23992 8916 23998 8968
rect 24044 8965 24072 9064
rect 25130 9052 25136 9104
rect 25188 9092 25194 9104
rect 25498 9092 25504 9104
rect 25188 9064 25504 9092
rect 25188 9052 25194 9064
rect 25498 9052 25504 9064
rect 25556 9052 25562 9104
rect 26326 9052 26332 9104
rect 26384 9092 26390 9104
rect 28966 9092 28994 9132
rect 33870 9120 33876 9132
rect 33928 9120 33934 9172
rect 37734 9120 37740 9172
rect 37792 9120 37798 9172
rect 38010 9120 38016 9172
rect 38068 9160 38074 9172
rect 38068 9132 41000 9160
rect 38068 9120 38074 9132
rect 31846 9092 31852 9104
rect 26384 9064 28994 9092
rect 31128 9064 31852 9092
rect 26384 9052 26390 9064
rect 24765 9027 24823 9033
rect 24765 8993 24777 9027
rect 24811 9024 24823 9027
rect 24946 9024 24952 9036
rect 24811 8996 24952 9024
rect 24811 8993 24823 8996
rect 24765 8987 24823 8993
rect 24946 8984 24952 8996
rect 25004 9024 25010 9036
rect 26050 9024 26056 9036
rect 25004 8996 26056 9024
rect 25004 8984 25010 8996
rect 24029 8959 24087 8965
rect 24029 8925 24041 8959
rect 24075 8925 24087 8959
rect 24029 8919 24087 8925
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8956 24639 8959
rect 25038 8956 25044 8968
rect 24627 8928 25044 8956
rect 24627 8925 24639 8928
rect 24581 8919 24639 8925
rect 25038 8916 25044 8928
rect 25096 8916 25102 8968
rect 25130 8916 25136 8968
rect 25188 8916 25194 8968
rect 25240 8928 25544 8956
rect 22646 8888 22652 8900
rect 20364 8860 22652 8888
rect 22646 8848 22652 8860
rect 22704 8848 22710 8900
rect 23474 8848 23480 8900
rect 23532 8848 23538 8900
rect 23658 8848 23664 8900
rect 23716 8848 23722 8900
rect 25240 8888 25268 8928
rect 23768 8860 25268 8888
rect 25317 8891 25375 8897
rect 18472 8792 18644 8820
rect 18472 8780 18478 8792
rect 20898 8780 20904 8832
rect 20956 8780 20962 8832
rect 23768 8829 23796 8860
rect 25317 8857 25329 8891
rect 25363 8888 25375 8891
rect 25406 8888 25412 8900
rect 25363 8860 25412 8888
rect 25363 8857 25375 8860
rect 25317 8851 25375 8857
rect 25406 8848 25412 8860
rect 25464 8848 25470 8900
rect 25516 8888 25544 8928
rect 25774 8916 25780 8968
rect 25832 8956 25838 8968
rect 25976 8965 26004 8996
rect 26050 8984 26056 8996
rect 26108 8984 26114 9036
rect 26421 9027 26479 9033
rect 26421 8993 26433 9027
rect 26467 9024 26479 9027
rect 26970 9024 26976 9036
rect 26467 8996 26976 9024
rect 26467 8993 26479 8996
rect 26421 8987 26479 8993
rect 26970 8984 26976 8996
rect 27028 8984 27034 9036
rect 28810 8984 28816 9036
rect 28868 9024 28874 9036
rect 28994 9024 29000 9036
rect 28868 8996 29000 9024
rect 28868 8984 28874 8996
rect 28994 8984 29000 8996
rect 29052 8984 29058 9036
rect 29086 8984 29092 9036
rect 29144 9024 29150 9036
rect 31128 9024 31156 9064
rect 31846 9052 31852 9064
rect 31904 9052 31910 9104
rect 32950 9052 32956 9104
rect 33008 9092 33014 9104
rect 33045 9095 33103 9101
rect 33045 9092 33057 9095
rect 33008 9064 33057 9092
rect 33008 9052 33014 9064
rect 33045 9061 33057 9064
rect 33091 9061 33103 9095
rect 33045 9055 33103 9061
rect 33134 9052 33140 9104
rect 33192 9092 33198 9104
rect 33965 9095 34023 9101
rect 33965 9092 33977 9095
rect 33192 9064 33977 9092
rect 33192 9052 33198 9064
rect 33965 9061 33977 9064
rect 34011 9061 34023 9095
rect 33965 9055 34023 9061
rect 35802 9052 35808 9104
rect 35860 9052 35866 9104
rect 38286 9052 38292 9104
rect 38344 9092 38350 9104
rect 38654 9092 38660 9104
rect 38344 9064 38660 9092
rect 38344 9052 38350 9064
rect 38654 9052 38660 9064
rect 38712 9052 38718 9104
rect 40972 9092 41000 9132
rect 41414 9120 41420 9172
rect 41472 9160 41478 9172
rect 52362 9160 52368 9172
rect 41472 9132 52368 9160
rect 41472 9120 41478 9132
rect 52362 9120 52368 9132
rect 52420 9120 52426 9172
rect 58342 9160 58348 9172
rect 54680 9132 58348 9160
rect 42702 9092 42708 9104
rect 40972 9064 42708 9092
rect 42702 9052 42708 9064
rect 42760 9052 42766 9104
rect 43898 9052 43904 9104
rect 43956 9092 43962 9104
rect 44910 9092 44916 9104
rect 43956 9064 44916 9092
rect 43956 9052 43962 9064
rect 44910 9052 44916 9064
rect 44968 9092 44974 9104
rect 54680 9092 54708 9132
rect 58342 9120 58348 9132
rect 58400 9120 58406 9172
rect 44968 9064 54708 9092
rect 56137 9095 56195 9101
rect 44968 9052 44974 9064
rect 56137 9061 56149 9095
rect 56183 9092 56195 9095
rect 56183 9064 56824 9092
rect 56183 9061 56195 9064
rect 56137 9055 56195 9061
rect 29144 8996 31156 9024
rect 29144 8984 29150 8996
rect 31386 8984 31392 9036
rect 31444 9024 31450 9036
rect 35820 9024 35848 9052
rect 31444 8996 35848 9024
rect 31444 8984 31450 8996
rect 36262 8984 36268 9036
rect 36320 8984 36326 9036
rect 36722 8984 36728 9036
rect 36780 9024 36786 9036
rect 36780 8996 37596 9024
rect 36780 8984 36786 8996
rect 25869 8959 25927 8965
rect 25869 8956 25881 8959
rect 25832 8928 25881 8956
rect 25832 8916 25838 8928
rect 25869 8925 25881 8928
rect 25915 8925 25927 8959
rect 25869 8919 25927 8925
rect 25961 8959 26019 8965
rect 25961 8925 25973 8959
rect 26007 8925 26019 8959
rect 26602 8956 26608 8968
rect 25961 8919 26019 8925
rect 26068 8928 26608 8956
rect 26068 8888 26096 8928
rect 26602 8916 26608 8928
rect 26660 8916 26666 8968
rect 27801 8959 27859 8965
rect 27801 8925 27813 8959
rect 27847 8956 27859 8959
rect 27890 8956 27896 8968
rect 27847 8928 27896 8956
rect 27847 8925 27859 8928
rect 27801 8919 27859 8925
rect 27890 8916 27896 8928
rect 27948 8916 27954 8968
rect 27985 8959 28043 8965
rect 27985 8925 27997 8959
rect 28031 8956 28043 8959
rect 29178 8956 29184 8968
rect 28031 8928 29184 8956
rect 28031 8925 28043 8928
rect 27985 8919 28043 8925
rect 29178 8916 29184 8928
rect 29236 8916 29242 8968
rect 30834 8916 30840 8968
rect 30892 8956 30898 8968
rect 31113 8959 31171 8965
rect 31113 8956 31125 8959
rect 30892 8928 31125 8956
rect 30892 8916 30898 8928
rect 31113 8925 31125 8928
rect 31159 8925 31171 8959
rect 31113 8919 31171 8925
rect 31297 8959 31355 8965
rect 31297 8925 31309 8959
rect 31343 8956 31355 8959
rect 31478 8956 31484 8968
rect 31343 8928 31484 8956
rect 31343 8925 31355 8928
rect 31297 8919 31355 8925
rect 31478 8916 31484 8928
rect 31536 8956 31542 8968
rect 31846 8956 31852 8968
rect 31536 8928 31852 8956
rect 31536 8916 31542 8928
rect 31846 8916 31852 8928
rect 31904 8916 31910 8968
rect 32122 8916 32128 8968
rect 32180 8916 32186 8968
rect 32582 8916 32588 8968
rect 32640 8956 32646 8968
rect 33321 8959 33379 8965
rect 33321 8956 33333 8959
rect 32640 8928 33333 8956
rect 32640 8916 32646 8928
rect 33321 8925 33333 8928
rect 33367 8956 33379 8959
rect 33410 8956 33416 8968
rect 33367 8928 33416 8956
rect 33367 8925 33379 8928
rect 33321 8919 33379 8925
rect 33410 8916 33416 8928
rect 33468 8916 33474 8968
rect 33505 8959 33563 8965
rect 33505 8925 33517 8959
rect 33551 8925 33563 8959
rect 33505 8919 33563 8925
rect 25516 8860 26096 8888
rect 26234 8848 26240 8900
rect 26292 8888 26298 8900
rect 27706 8888 27712 8900
rect 26292 8860 27712 8888
rect 26292 8848 26298 8860
rect 27706 8848 27712 8860
rect 27764 8848 27770 8900
rect 28905 8891 28963 8897
rect 28905 8888 28917 8891
rect 27816 8860 28917 8888
rect 23753 8823 23811 8829
rect 23753 8789 23765 8823
rect 23799 8789 23811 8823
rect 23753 8783 23811 8789
rect 23845 8823 23903 8829
rect 23845 8789 23857 8823
rect 23891 8820 23903 8823
rect 24026 8820 24032 8832
rect 23891 8792 24032 8820
rect 23891 8789 23903 8792
rect 23845 8783 23903 8789
rect 24026 8780 24032 8792
rect 24084 8780 24090 8832
rect 24946 8780 24952 8832
rect 25004 8820 25010 8832
rect 25225 8823 25283 8829
rect 25225 8820 25237 8823
rect 25004 8792 25237 8820
rect 25004 8780 25010 8792
rect 25225 8789 25237 8792
rect 25271 8820 25283 8823
rect 26694 8820 26700 8832
rect 25271 8792 26700 8820
rect 25271 8789 25283 8792
rect 25225 8783 25283 8789
rect 26694 8780 26700 8792
rect 26752 8780 26758 8832
rect 27522 8780 27528 8832
rect 27580 8820 27586 8832
rect 27816 8820 27844 8860
rect 28905 8857 28917 8860
rect 28951 8857 28963 8891
rect 28905 8851 28963 8857
rect 29730 8848 29736 8900
rect 29788 8848 29794 8900
rect 29822 8848 29828 8900
rect 29880 8888 29886 8900
rect 30469 8891 30527 8897
rect 30469 8888 30481 8891
rect 29880 8860 30481 8888
rect 29880 8848 29886 8860
rect 30469 8857 30481 8860
rect 30515 8857 30527 8891
rect 30469 8851 30527 8857
rect 31662 8848 31668 8900
rect 31720 8848 31726 8900
rect 32398 8848 32404 8900
rect 32456 8888 32462 8900
rect 32674 8888 32680 8900
rect 32456 8860 32680 8888
rect 32456 8848 32462 8860
rect 32674 8848 32680 8860
rect 32732 8848 32738 8900
rect 33520 8888 33548 8919
rect 34146 8916 34152 8968
rect 34204 8916 34210 8968
rect 34238 8916 34244 8968
rect 34296 8916 34302 8968
rect 35802 8916 35808 8968
rect 35860 8916 35866 8968
rect 35894 8916 35900 8968
rect 35952 8956 35958 8968
rect 36354 8956 36360 8968
rect 35952 8928 36360 8956
rect 35952 8916 35958 8928
rect 36354 8916 36360 8928
rect 36412 8916 36418 8968
rect 37182 8916 37188 8968
rect 37240 8916 37246 8968
rect 37458 8916 37464 8968
rect 37516 8916 37522 8968
rect 37568 8965 37596 8996
rect 37826 8984 37832 9036
rect 37884 9024 37890 9036
rect 38102 9024 38108 9036
rect 37884 8996 38108 9024
rect 37884 8984 37890 8996
rect 38102 8984 38108 8996
rect 38160 8984 38166 9036
rect 40034 8984 40040 9036
rect 40092 8984 40098 9036
rect 41386 8996 51074 9024
rect 37553 8959 37611 8965
rect 37553 8925 37565 8959
rect 37599 8925 37611 8959
rect 37553 8919 37611 8925
rect 38562 8916 38568 8968
rect 38620 8956 38626 8968
rect 38841 8959 38899 8965
rect 38841 8956 38853 8959
rect 38620 8928 38853 8956
rect 38620 8916 38626 8928
rect 38841 8925 38853 8928
rect 38887 8956 38899 8959
rect 40126 8956 40132 8968
rect 38887 8928 40132 8956
rect 38887 8925 38899 8928
rect 38841 8919 38899 8925
rect 40126 8916 40132 8928
rect 40184 8916 40190 8968
rect 41386 8956 41414 8996
rect 40236 8928 41414 8956
rect 33152 8860 33548 8888
rect 27580 8792 27844 8820
rect 28813 8823 28871 8829
rect 27580 8780 27586 8792
rect 28813 8789 28825 8823
rect 28859 8820 28871 8823
rect 29546 8820 29552 8832
rect 28859 8792 29552 8820
rect 28859 8789 28871 8792
rect 28813 8783 28871 8789
rect 29546 8780 29552 8792
rect 29604 8820 29610 8832
rect 30650 8820 30656 8832
rect 29604 8792 30656 8820
rect 29604 8780 29610 8792
rect 30650 8780 30656 8792
rect 30708 8780 30714 8832
rect 31386 8780 31392 8832
rect 31444 8780 31450 8832
rect 31478 8780 31484 8832
rect 31536 8820 31542 8832
rect 33152 8820 33180 8860
rect 33962 8848 33968 8900
rect 34020 8848 34026 8900
rect 37369 8891 37427 8897
rect 37369 8857 37381 8891
rect 37415 8888 37427 8891
rect 38194 8888 38200 8900
rect 37415 8860 38200 8888
rect 37415 8857 37427 8860
rect 37369 8851 37427 8857
rect 38194 8848 38200 8860
rect 38252 8848 38258 8900
rect 40236 8888 40264 8928
rect 44450 8916 44456 8968
rect 44508 8916 44514 8968
rect 44542 8916 44548 8968
rect 44600 8956 44606 8968
rect 45189 8959 45247 8965
rect 45189 8956 45201 8959
rect 44600 8928 45201 8956
rect 44600 8916 44606 8928
rect 45189 8925 45201 8928
rect 45235 8925 45247 8959
rect 45189 8919 45247 8925
rect 46106 8916 46112 8968
rect 46164 8916 46170 8968
rect 46290 8916 46296 8968
rect 46348 8916 46354 8968
rect 38672 8860 40264 8888
rect 40304 8891 40362 8897
rect 31536 8792 33180 8820
rect 31536 8780 31542 8792
rect 33226 8780 33232 8832
rect 33284 8780 33290 8832
rect 35989 8823 36047 8829
rect 35989 8789 36001 8823
rect 36035 8820 36047 8823
rect 38672 8820 38700 8860
rect 40304 8857 40316 8891
rect 40350 8857 40362 8891
rect 40304 8851 40362 8857
rect 36035 8792 38700 8820
rect 36035 8789 36047 8792
rect 35989 8783 36047 8789
rect 38930 8780 38936 8832
rect 38988 8820 38994 8832
rect 40328 8820 40356 8851
rect 43714 8848 43720 8900
rect 43772 8848 43778 8900
rect 44174 8848 44180 8900
rect 44232 8888 44238 8900
rect 45465 8891 45523 8897
rect 45465 8888 45477 8891
rect 44232 8860 45477 8888
rect 44232 8848 44238 8860
rect 45465 8857 45477 8860
rect 45511 8857 45523 8891
rect 46308 8888 46336 8916
rect 45465 8851 45523 8857
rect 45572 8860 46336 8888
rect 51046 8888 51074 8996
rect 56134 8916 56140 8968
rect 56192 8916 56198 8968
rect 56318 8916 56324 8968
rect 56376 8916 56382 8968
rect 56413 8959 56471 8965
rect 56413 8925 56425 8959
rect 56459 8925 56471 8959
rect 56796 8956 56824 9064
rect 56870 8984 56876 9036
rect 56928 8984 56934 9036
rect 57129 8959 57187 8965
rect 57129 8956 57141 8959
rect 56796 8928 57141 8956
rect 56413 8919 56471 8925
rect 57129 8925 57141 8928
rect 57175 8925 57187 8959
rect 57129 8919 57187 8925
rect 52270 8888 52276 8900
rect 51046 8860 52276 8888
rect 38988 8792 40356 8820
rect 38988 8780 38994 8792
rect 43898 8780 43904 8832
rect 43956 8820 43962 8832
rect 45572 8820 45600 8860
rect 52270 8848 52276 8860
rect 52328 8848 52334 8900
rect 43956 8792 45600 8820
rect 46293 8823 46351 8829
rect 43956 8780 43962 8792
rect 46293 8789 46305 8823
rect 46339 8820 46351 8823
rect 46658 8820 46664 8832
rect 46339 8792 46664 8820
rect 46339 8789 46351 8792
rect 46293 8783 46351 8789
rect 46658 8780 46664 8792
rect 46716 8780 46722 8832
rect 52362 8780 52368 8832
rect 52420 8820 52426 8832
rect 56428 8820 56456 8919
rect 52420 8792 56456 8820
rect 52420 8780 52426 8792
rect 57238 8780 57244 8832
rect 57296 8820 57302 8832
rect 58253 8823 58311 8829
rect 58253 8820 58265 8823
rect 57296 8792 58265 8820
rect 57296 8780 57302 8792
rect 58253 8789 58265 8792
rect 58299 8789 58311 8823
rect 58253 8783 58311 8789
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 14093 8619 14151 8625
rect 14093 8616 14105 8619
rect 13504 8588 14105 8616
rect 13504 8576 13510 8588
rect 14093 8585 14105 8588
rect 14139 8585 14151 8619
rect 14093 8579 14151 8585
rect 15013 8619 15071 8625
rect 15013 8585 15025 8619
rect 15059 8616 15071 8619
rect 15102 8616 15108 8628
rect 15059 8588 15108 8616
rect 15059 8585 15071 8588
rect 15013 8579 15071 8585
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15286 8576 15292 8628
rect 15344 8616 15350 8628
rect 15344 8588 17264 8616
rect 15344 8576 15350 8588
rect 16298 8548 16304 8560
rect 14936 8520 16304 8548
rect 1581 8483 1639 8489
rect 1581 8449 1593 8483
rect 1627 8480 1639 8483
rect 10594 8480 10600 8492
rect 1627 8452 10600 8480
rect 1627 8449 1639 8452
rect 1581 8443 1639 8449
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 13998 8440 14004 8492
rect 14056 8440 14062 8492
rect 14936 8489 14964 8520
rect 16298 8508 16304 8520
rect 16356 8508 16362 8560
rect 16942 8508 16948 8560
rect 17000 8508 17006 8560
rect 17236 8548 17264 8588
rect 17402 8576 17408 8628
rect 17460 8576 17466 8628
rect 17494 8576 17500 8628
rect 17552 8616 17558 8628
rect 18046 8616 18052 8628
rect 17552 8588 18052 8616
rect 17552 8576 17558 8588
rect 18046 8576 18052 8588
rect 18104 8616 18110 8628
rect 18104 8588 19012 8616
rect 18104 8576 18110 8588
rect 18414 8548 18420 8560
rect 17236 8520 18420 8548
rect 18414 8508 18420 8520
rect 18472 8548 18478 8560
rect 18472 8520 18644 8548
rect 18472 8508 18478 8520
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8480 15715 8483
rect 17681 8483 17739 8489
rect 17681 8480 17693 8483
rect 15703 8452 17693 8480
rect 15703 8449 15715 8452
rect 15657 8443 15715 8449
rect 17681 8449 17693 8452
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 18616 8489 18644 8520
rect 18984 8489 19012 8588
rect 19150 8576 19156 8628
rect 19208 8616 19214 8628
rect 19337 8619 19395 8625
rect 19337 8616 19349 8619
rect 19208 8588 19349 8616
rect 19208 8576 19214 8588
rect 19337 8585 19349 8588
rect 19383 8585 19395 8619
rect 19337 8579 19395 8585
rect 20254 8576 20260 8628
rect 20312 8576 20318 8628
rect 20625 8619 20683 8625
rect 20625 8585 20637 8619
rect 20671 8616 20683 8619
rect 21174 8616 21180 8628
rect 20671 8588 21180 8616
rect 20671 8585 20683 8588
rect 20625 8579 20683 8585
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 23382 8576 23388 8628
rect 23440 8616 23446 8628
rect 23569 8619 23627 8625
rect 23569 8616 23581 8619
rect 23440 8588 23581 8616
rect 23440 8576 23446 8588
rect 23569 8585 23581 8588
rect 23615 8585 23627 8619
rect 23569 8579 23627 8585
rect 23661 8619 23719 8625
rect 23661 8585 23673 8619
rect 23707 8616 23719 8619
rect 23707 8588 23886 8616
rect 23707 8585 23719 8588
rect 23661 8579 23719 8585
rect 19242 8508 19248 8560
rect 19300 8548 19306 8560
rect 20717 8551 20775 8557
rect 20717 8548 20729 8551
rect 19300 8520 20729 8548
rect 19300 8508 19306 8520
rect 20717 8517 20729 8520
rect 20763 8548 20775 8551
rect 20898 8548 20904 8560
rect 20763 8520 20904 8548
rect 20763 8517 20775 8520
rect 20717 8511 20775 8517
rect 20898 8508 20904 8520
rect 20956 8508 20962 8560
rect 23290 8508 23296 8560
rect 23348 8508 23354 8560
rect 23858 8548 23886 8588
rect 25314 8576 25320 8628
rect 25372 8576 25378 8628
rect 25958 8576 25964 8628
rect 26016 8576 26022 8628
rect 26145 8619 26203 8625
rect 26145 8585 26157 8619
rect 26191 8616 26203 8619
rect 26510 8616 26516 8628
rect 26191 8588 26372 8616
rect 26191 8585 26203 8588
rect 26145 8579 26203 8585
rect 24026 8548 24032 8560
rect 23858 8520 24032 8548
rect 24026 8508 24032 8520
rect 24084 8548 24090 8560
rect 26255 8551 26313 8557
rect 26255 8548 26267 8551
rect 24084 8520 26267 8548
rect 24084 8508 24090 8520
rect 26255 8517 26267 8520
rect 26301 8517 26313 8551
rect 26255 8511 26313 8517
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 17920 8452 18245 8480
rect 17920 8440 17926 8452
rect 18233 8449 18245 8452
rect 18279 8449 18291 8483
rect 18233 8443 18291 8449
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8449 18659 8483
rect 18601 8443 18659 8449
rect 18969 8483 19027 8489
rect 18969 8449 18981 8483
rect 19015 8449 19027 8483
rect 19797 8483 19855 8489
rect 19797 8480 19809 8483
rect 18969 8443 19027 8449
rect 19306 8452 19809 8480
rect 934 8372 940 8424
rect 992 8412 998 8424
rect 1765 8415 1823 8421
rect 1765 8412 1777 8415
rect 992 8384 1777 8412
rect 992 8372 998 8384
rect 1765 8381 1777 8384
rect 1811 8381 1823 8415
rect 14016 8412 14044 8440
rect 15286 8412 15292 8424
rect 14016 8384 15292 8412
rect 1765 8375 1823 8381
rect 15286 8372 15292 8384
rect 15344 8372 15350 8424
rect 16206 8372 16212 8424
rect 16264 8372 16270 8424
rect 16298 8372 16304 8424
rect 16356 8412 16362 8424
rect 16356 8384 17080 8412
rect 16356 8372 16362 8384
rect 16945 8347 17003 8353
rect 16945 8313 16957 8347
rect 16991 8344 17003 8347
rect 17052 8344 17080 8384
rect 17402 8344 17408 8356
rect 16991 8316 17408 8344
rect 16991 8313 17003 8316
rect 16945 8307 17003 8313
rect 17402 8304 17408 8316
rect 17460 8344 17466 8356
rect 19306 8344 19334 8452
rect 19797 8449 19809 8452
rect 19843 8480 19855 8483
rect 23477 8483 23535 8489
rect 19843 8452 23428 8480
rect 19843 8449 19855 8452
rect 19797 8443 19855 8449
rect 20901 8415 20959 8421
rect 20901 8381 20913 8415
rect 20947 8412 20959 8415
rect 21266 8412 21272 8424
rect 20947 8384 21272 8412
rect 20947 8381 20959 8384
rect 20901 8375 20959 8381
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 23400 8412 23428 8452
rect 23477 8449 23489 8483
rect 23523 8480 23535 8483
rect 23566 8480 23572 8492
rect 23523 8452 23572 8480
rect 23523 8449 23535 8452
rect 23477 8443 23535 8449
rect 23566 8440 23572 8452
rect 23624 8440 23630 8492
rect 23658 8440 23664 8492
rect 23716 8480 23722 8492
rect 23845 8483 23903 8489
rect 23845 8480 23857 8483
rect 23716 8452 23857 8480
rect 23716 8440 23722 8452
rect 23845 8449 23857 8452
rect 23891 8449 23903 8483
rect 23845 8443 23903 8449
rect 24302 8440 24308 8492
rect 24360 8440 24366 8492
rect 24486 8440 24492 8492
rect 24544 8440 24550 8492
rect 25133 8483 25191 8489
rect 25133 8449 25145 8483
rect 25179 8449 25191 8483
rect 25133 8443 25191 8449
rect 24946 8412 24952 8424
rect 23400 8384 24952 8412
rect 24946 8372 24952 8384
rect 25004 8372 25010 8424
rect 25148 8412 25176 8443
rect 26050 8440 26056 8492
rect 26108 8440 26114 8492
rect 25866 8412 25872 8424
rect 25148 8384 25872 8412
rect 25866 8372 25872 8384
rect 25924 8372 25930 8424
rect 26270 8412 26298 8511
rect 26344 8480 26372 8588
rect 26436 8588 26516 8616
rect 26436 8557 26464 8588
rect 26510 8576 26516 8588
rect 26568 8576 26574 8628
rect 27706 8576 27712 8628
rect 27764 8616 27770 8628
rect 28718 8616 28724 8628
rect 27764 8588 28724 8616
rect 27764 8576 27770 8588
rect 28718 8576 28724 8588
rect 28776 8576 28782 8628
rect 31294 8576 31300 8628
rect 31352 8576 31358 8628
rect 31389 8619 31447 8625
rect 31389 8585 31401 8619
rect 31435 8616 31447 8619
rect 31478 8616 31484 8628
rect 31435 8588 31484 8616
rect 31435 8585 31447 8588
rect 31389 8579 31447 8585
rect 31478 8576 31484 8588
rect 31536 8616 31542 8628
rect 31938 8616 31944 8628
rect 31536 8588 31944 8616
rect 31536 8576 31542 8588
rect 31938 8576 31944 8588
rect 31996 8576 32002 8628
rect 32858 8576 32864 8628
rect 32916 8576 32922 8628
rect 33318 8616 33324 8628
rect 33152 8588 33324 8616
rect 26421 8551 26479 8557
rect 26421 8517 26433 8551
rect 26467 8517 26479 8551
rect 26421 8511 26479 8517
rect 27525 8551 27583 8557
rect 27525 8517 27537 8551
rect 27571 8548 27583 8551
rect 28905 8551 28963 8557
rect 28905 8548 28917 8551
rect 27571 8520 28917 8548
rect 27571 8517 27583 8520
rect 27525 8511 27583 8517
rect 28905 8517 28917 8520
rect 28951 8548 28963 8551
rect 29086 8548 29092 8560
rect 28951 8520 29092 8548
rect 28951 8517 28963 8520
rect 28905 8511 28963 8517
rect 29086 8508 29092 8520
rect 29144 8508 29150 8560
rect 30926 8508 30932 8560
rect 30984 8548 30990 8560
rect 31021 8551 31079 8557
rect 31021 8548 31033 8551
rect 30984 8520 31033 8548
rect 30984 8508 30990 8520
rect 31021 8517 31033 8520
rect 31067 8517 31079 8551
rect 31021 8511 31079 8517
rect 31205 8551 31263 8557
rect 31205 8517 31217 8551
rect 31251 8548 31263 8551
rect 31846 8548 31852 8560
rect 31251 8520 31852 8548
rect 31251 8517 31263 8520
rect 31205 8511 31263 8517
rect 31846 8508 31852 8520
rect 31904 8508 31910 8560
rect 32876 8548 32904 8576
rect 33152 8557 33180 8588
rect 33318 8576 33324 8588
rect 33376 8576 33382 8628
rect 33413 8619 33471 8625
rect 33413 8585 33425 8619
rect 33459 8616 33471 8619
rect 35802 8616 35808 8628
rect 33459 8588 35808 8616
rect 33459 8585 33471 8588
rect 33413 8579 33471 8585
rect 35802 8576 35808 8588
rect 35860 8576 35866 8628
rect 36538 8576 36544 8628
rect 36596 8616 36602 8628
rect 38749 8619 38807 8625
rect 36596 8588 37964 8616
rect 36596 8576 36602 8588
rect 32784 8520 32904 8548
rect 33137 8551 33195 8557
rect 27246 8480 27252 8492
rect 26344 8452 27252 8480
rect 27246 8440 27252 8452
rect 27304 8440 27310 8492
rect 27338 8440 27344 8492
rect 27396 8440 27402 8492
rect 27614 8440 27620 8492
rect 27672 8440 27678 8492
rect 27706 8440 27712 8492
rect 27764 8440 27770 8492
rect 27982 8440 27988 8492
rect 28040 8480 28046 8492
rect 28166 8480 28172 8492
rect 28040 8452 28172 8480
rect 28040 8440 28046 8452
rect 28166 8440 28172 8452
rect 28224 8440 28230 8492
rect 28445 8483 28503 8489
rect 28445 8449 28457 8483
rect 28491 8480 28503 8483
rect 29178 8480 29184 8492
rect 28491 8452 29184 8480
rect 28491 8449 28503 8452
rect 28445 8443 28503 8449
rect 29178 8440 29184 8452
rect 29236 8440 29242 8492
rect 29546 8440 29552 8492
rect 29604 8440 29610 8492
rect 31570 8440 31576 8492
rect 31628 8440 31634 8492
rect 32784 8489 32812 8520
rect 33137 8517 33149 8551
rect 33183 8517 33195 8551
rect 35434 8548 35440 8560
rect 33137 8511 33195 8517
rect 34164 8520 35440 8548
rect 34164 8492 34192 8520
rect 35434 8508 35440 8520
rect 35492 8508 35498 8560
rect 36354 8548 36360 8560
rect 35912 8520 36360 8548
rect 32769 8483 32827 8489
rect 32769 8449 32781 8483
rect 32815 8449 32827 8483
rect 32769 8443 32827 8449
rect 32858 8440 32864 8492
rect 32916 8480 32922 8492
rect 32916 8452 32961 8480
rect 32916 8440 32922 8452
rect 33042 8440 33048 8492
rect 33100 8440 33106 8492
rect 33234 8483 33292 8489
rect 33234 8449 33246 8483
rect 33280 8449 33292 8483
rect 33234 8443 33292 8449
rect 28258 8412 28264 8424
rect 26270 8384 28264 8412
rect 28258 8372 28264 8384
rect 28316 8372 28322 8424
rect 28718 8372 28724 8424
rect 28776 8412 28782 8424
rect 29914 8412 29920 8424
rect 28776 8384 29920 8412
rect 28776 8372 28782 8384
rect 29914 8372 29920 8384
rect 29972 8372 29978 8424
rect 33249 8412 33277 8443
rect 33870 8440 33876 8492
rect 33928 8440 33934 8492
rect 33962 8440 33968 8492
rect 34020 8480 34026 8492
rect 34020 8452 34065 8480
rect 34020 8440 34026 8452
rect 34146 8440 34152 8492
rect 34204 8440 34210 8492
rect 34241 8483 34299 8489
rect 34241 8449 34253 8483
rect 34287 8449 34299 8483
rect 34241 8443 34299 8449
rect 33244 8384 33277 8412
rect 34256 8412 34284 8443
rect 34330 8440 34336 8492
rect 34388 8489 34394 8492
rect 35912 8489 35940 8520
rect 36354 8508 36360 8520
rect 36412 8548 36418 8560
rect 37366 8548 37372 8560
rect 36412 8520 37372 8548
rect 36412 8508 36418 8520
rect 37366 8508 37372 8520
rect 37424 8508 37430 8560
rect 37936 8548 37964 8588
rect 38749 8585 38761 8619
rect 38795 8616 38807 8619
rect 38930 8616 38936 8628
rect 38795 8588 38936 8616
rect 38795 8585 38807 8588
rect 38749 8579 38807 8585
rect 38930 8576 38936 8588
rect 38988 8576 38994 8628
rect 40037 8619 40095 8625
rect 40037 8585 40049 8619
rect 40083 8616 40095 8619
rect 40586 8616 40592 8628
rect 40083 8588 40592 8616
rect 40083 8585 40095 8588
rect 40037 8579 40095 8585
rect 40586 8576 40592 8588
rect 40644 8576 40650 8628
rect 44174 8616 44180 8628
rect 42444 8588 44180 8616
rect 37476 8520 37872 8548
rect 37936 8520 39620 8548
rect 34388 8480 34396 8489
rect 35897 8483 35955 8489
rect 34388 8452 34433 8480
rect 34388 8443 34396 8452
rect 35897 8449 35909 8483
rect 35943 8449 35955 8483
rect 35897 8443 35955 8449
rect 34388 8440 34394 8443
rect 36722 8440 36728 8492
rect 36780 8440 36786 8492
rect 37476 8489 37504 8520
rect 37461 8483 37519 8489
rect 37461 8449 37473 8483
rect 37507 8449 37519 8483
rect 37461 8443 37519 8449
rect 37550 8440 37556 8492
rect 37608 8440 37614 8492
rect 37737 8483 37795 8489
rect 37737 8449 37749 8483
rect 37783 8449 37795 8483
rect 37844 8480 37872 8520
rect 38102 8480 38108 8492
rect 37844 8452 38108 8480
rect 37737 8443 37795 8449
rect 35345 8415 35403 8421
rect 35345 8412 35357 8415
rect 34256 8384 34376 8412
rect 17460 8316 19334 8344
rect 17460 8304 17466 8316
rect 23842 8304 23848 8356
rect 23900 8344 23906 8356
rect 24581 8347 24639 8353
rect 24581 8344 24593 8347
rect 23900 8316 24593 8344
rect 23900 8304 23906 8316
rect 24581 8313 24593 8316
rect 24627 8313 24639 8347
rect 28276 8344 28304 8372
rect 29822 8344 29828 8356
rect 28276 8316 29828 8344
rect 24581 8307 24639 8313
rect 29822 8304 29828 8316
rect 29880 8344 29886 8356
rect 30006 8344 30012 8356
rect 29880 8316 30012 8344
rect 29880 8304 29886 8316
rect 30006 8304 30012 8316
rect 30064 8304 30070 8356
rect 30834 8304 30840 8356
rect 30892 8344 30898 8356
rect 31754 8344 31760 8356
rect 30892 8316 31760 8344
rect 30892 8304 30898 8316
rect 31754 8304 31760 8316
rect 31812 8344 31818 8356
rect 33244 8344 33272 8384
rect 34348 8356 34376 8384
rect 34532 8384 35357 8412
rect 31812 8316 33272 8344
rect 31812 8304 31818 8316
rect 34330 8304 34336 8356
rect 34388 8304 34394 8356
rect 34532 8353 34560 8384
rect 35345 8381 35357 8384
rect 35391 8381 35403 8415
rect 35345 8375 35403 8381
rect 35710 8372 35716 8424
rect 35768 8372 35774 8424
rect 35802 8372 35808 8424
rect 35860 8372 35866 8424
rect 36541 8415 36599 8421
rect 36541 8381 36553 8415
rect 36587 8381 36599 8415
rect 36541 8375 36599 8381
rect 34517 8347 34575 8353
rect 34517 8313 34529 8347
rect 34563 8313 34575 8347
rect 36556 8344 36584 8375
rect 36630 8372 36636 8424
rect 36688 8412 36694 8424
rect 37752 8412 37780 8443
rect 38102 8440 38108 8452
rect 38160 8440 38166 8492
rect 38197 8483 38255 8489
rect 38197 8449 38209 8483
rect 38243 8480 38255 8483
rect 38286 8480 38292 8492
rect 38243 8452 38292 8480
rect 38243 8449 38255 8452
rect 38197 8443 38255 8449
rect 38286 8440 38292 8452
rect 38344 8440 38350 8492
rect 38930 8440 38936 8492
rect 38988 8440 38994 8492
rect 39206 8440 39212 8492
rect 39264 8440 39270 8492
rect 39393 8483 39451 8489
rect 39393 8449 39405 8483
rect 39439 8449 39451 8483
rect 39592 8480 39620 8520
rect 39666 8508 39672 8560
rect 39724 8548 39730 8560
rect 39853 8551 39911 8557
rect 39853 8548 39865 8551
rect 39724 8520 39865 8548
rect 39724 8508 39730 8520
rect 39853 8517 39865 8520
rect 39899 8517 39911 8551
rect 39853 8511 39911 8517
rect 39942 8480 39948 8492
rect 39592 8452 39948 8480
rect 39393 8443 39451 8449
rect 39298 8412 39304 8424
rect 36688 8384 37780 8412
rect 37844 8384 39304 8412
rect 36688 8372 36694 8384
rect 37734 8344 37740 8356
rect 36556 8316 37740 8344
rect 34517 8307 34575 8313
rect 37734 8304 37740 8316
rect 37792 8344 37798 8356
rect 37844 8344 37872 8384
rect 39298 8372 39304 8384
rect 39356 8372 39362 8424
rect 39408 8412 39436 8443
rect 39942 8440 39948 8452
rect 40000 8440 40006 8492
rect 40129 8483 40187 8489
rect 40129 8470 40141 8483
rect 40052 8449 40141 8470
rect 40175 8480 40187 8483
rect 42444 8480 42472 8588
rect 44174 8576 44180 8588
rect 44232 8576 44238 8628
rect 44269 8619 44327 8625
rect 44269 8585 44281 8619
rect 44315 8616 44327 8619
rect 46106 8616 46112 8628
rect 44315 8588 46112 8616
rect 44315 8585 44327 8588
rect 44269 8579 44327 8585
rect 46106 8576 46112 8588
rect 46164 8576 46170 8628
rect 46198 8576 46204 8628
rect 46256 8616 46262 8628
rect 58894 8616 58900 8628
rect 46256 8588 58900 8616
rect 46256 8576 46262 8588
rect 58894 8576 58900 8588
rect 58952 8576 58958 8628
rect 42702 8508 42708 8560
rect 42760 8548 42766 8560
rect 43165 8551 43223 8557
rect 43165 8548 43177 8551
rect 42760 8520 43177 8548
rect 42760 8508 42766 8520
rect 43165 8517 43177 8520
rect 43211 8517 43223 8551
rect 43165 8511 43223 8517
rect 43622 8508 43628 8560
rect 43680 8548 43686 8560
rect 44910 8548 44916 8560
rect 43680 8520 44220 8548
rect 43680 8508 43686 8520
rect 40175 8452 42472 8480
rect 42797 8483 42855 8489
rect 40175 8449 40187 8452
rect 40052 8443 40187 8449
rect 42797 8449 42809 8483
rect 42843 8480 42855 8483
rect 43806 8480 43812 8492
rect 42843 8452 43812 8480
rect 42843 8449 42855 8452
rect 42797 8443 42855 8449
rect 40052 8442 40181 8443
rect 39408 8384 39896 8412
rect 37792 8316 37872 8344
rect 37792 8304 37798 8316
rect 38654 8304 38660 8356
rect 38712 8344 38718 8356
rect 39868 8353 39896 8384
rect 39025 8347 39083 8353
rect 39025 8344 39037 8347
rect 38712 8316 39037 8344
rect 38712 8304 38718 8316
rect 39025 8313 39037 8316
rect 39071 8313 39083 8347
rect 39025 8307 39083 8313
rect 39117 8347 39175 8353
rect 39117 8313 39129 8347
rect 39163 8313 39175 8347
rect 39117 8307 39175 8313
rect 39853 8347 39911 8353
rect 39853 8313 39865 8347
rect 39899 8313 39911 8347
rect 40052 8344 40080 8442
rect 43806 8440 43812 8452
rect 43864 8440 43870 8492
rect 44192 8412 44220 8520
rect 44468 8520 44916 8548
rect 44468 8489 44496 8520
rect 44910 8508 44916 8520
rect 44968 8508 44974 8560
rect 57333 8551 57391 8557
rect 45296 8520 51074 8548
rect 44453 8483 44511 8489
rect 44453 8449 44465 8483
rect 44499 8449 44511 8483
rect 44453 8443 44511 8449
rect 44542 8440 44548 8492
rect 44600 8440 44606 8492
rect 44726 8440 44732 8492
rect 44784 8440 44790 8492
rect 45296 8489 45324 8520
rect 44821 8483 44879 8489
rect 44821 8449 44833 8483
rect 44867 8449 44879 8483
rect 44821 8443 44879 8449
rect 45281 8483 45339 8489
rect 45281 8449 45293 8483
rect 45327 8449 45339 8483
rect 45281 8443 45339 8449
rect 44836 8412 44864 8443
rect 46382 8440 46388 8492
rect 46440 8440 46446 8492
rect 45370 8412 45376 8424
rect 44192 8384 45376 8412
rect 45370 8372 45376 8384
rect 45428 8412 45434 8424
rect 45465 8415 45523 8421
rect 45465 8412 45477 8415
rect 45428 8384 45477 8412
rect 45428 8372 45434 8384
rect 45465 8381 45477 8384
rect 45511 8381 45523 8415
rect 45465 8375 45523 8381
rect 46106 8372 46112 8424
rect 46164 8412 46170 8424
rect 46569 8415 46627 8421
rect 46569 8412 46581 8415
rect 46164 8384 46581 8412
rect 46164 8372 46170 8384
rect 46569 8381 46581 8384
rect 46615 8381 46627 8415
rect 51046 8412 51074 8520
rect 57333 8517 57345 8551
rect 57379 8548 57391 8551
rect 58986 8548 58992 8560
rect 57379 8520 58992 8548
rect 57379 8517 57391 8520
rect 57333 8511 57391 8517
rect 58986 8508 58992 8520
rect 59044 8508 59050 8560
rect 56229 8483 56287 8489
rect 56229 8449 56241 8483
rect 56275 8449 56287 8483
rect 56229 8443 56287 8449
rect 57057 8483 57115 8489
rect 57057 8449 57069 8483
rect 57103 8480 57115 8483
rect 57238 8480 57244 8492
rect 57103 8452 57244 8480
rect 57103 8449 57115 8452
rect 57057 8443 57115 8449
rect 53098 8412 53104 8424
rect 51046 8384 53104 8412
rect 46569 8375 46627 8381
rect 53098 8372 53104 8384
rect 53156 8372 53162 8424
rect 56244 8412 56272 8443
rect 57238 8440 57244 8452
rect 57296 8440 57302 8492
rect 58986 8412 58992 8424
rect 56244 8384 58992 8412
rect 58986 8372 58992 8384
rect 59044 8372 59050 8424
rect 39853 8307 39911 8313
rect 39960 8316 40080 8344
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 22922 8276 22928 8288
rect 12952 8248 22928 8276
rect 12952 8236 12958 8248
rect 22922 8236 22928 8248
rect 22980 8236 22986 8288
rect 27430 8236 27436 8288
rect 27488 8276 27494 8288
rect 27614 8276 27620 8288
rect 27488 8248 27620 8276
rect 27488 8236 27494 8248
rect 27614 8236 27620 8248
rect 27672 8236 27678 8288
rect 27890 8236 27896 8288
rect 27948 8236 27954 8288
rect 28258 8236 28264 8288
rect 28316 8276 28322 8288
rect 32306 8276 32312 8288
rect 28316 8248 32312 8276
rect 28316 8236 28322 8248
rect 32306 8236 32312 8248
rect 32364 8236 32370 8288
rect 36262 8236 36268 8288
rect 36320 8276 36326 8288
rect 36538 8276 36544 8288
rect 36320 8248 36544 8276
rect 36320 8236 36326 8248
rect 36538 8236 36544 8248
rect 36596 8236 36602 8288
rect 36906 8236 36912 8288
rect 36964 8236 36970 8288
rect 37366 8236 37372 8288
rect 37424 8276 37430 8288
rect 39132 8276 39160 8307
rect 39960 8276 39988 8316
rect 40126 8304 40132 8356
rect 40184 8344 40190 8356
rect 43622 8344 43628 8356
rect 40184 8316 43628 8344
rect 40184 8304 40190 8316
rect 43622 8304 43628 8316
rect 43680 8304 43686 8356
rect 56410 8304 56416 8356
rect 56468 8304 56474 8356
rect 37424 8248 39988 8276
rect 37424 8236 37430 8248
rect 40034 8236 40040 8288
rect 40092 8276 40098 8288
rect 46290 8276 46296 8288
rect 40092 8248 46296 8276
rect 40092 8236 40098 8248
rect 46290 8236 46296 8248
rect 46348 8236 46354 8288
rect 54846 8236 54852 8288
rect 54904 8276 54910 8288
rect 58710 8276 58716 8288
rect 54904 8248 58716 8276
rect 54904 8236 54910 8248
rect 58710 8236 58716 8248
rect 58768 8236 58774 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 15933 8075 15991 8081
rect 15933 8041 15945 8075
rect 15979 8072 15991 8075
rect 19334 8072 19340 8084
rect 15979 8044 19340 8072
rect 15979 8041 15991 8044
rect 15933 8035 15991 8041
rect 19334 8032 19340 8044
rect 19392 8032 19398 8084
rect 25038 8032 25044 8084
rect 25096 8032 25102 8084
rect 25148 8044 25636 8072
rect 12802 7964 12808 8016
rect 12860 8004 12866 8016
rect 12897 8007 12955 8013
rect 12897 8004 12909 8007
rect 12860 7976 12909 8004
rect 12860 7964 12866 7976
rect 12897 7973 12909 7976
rect 12943 7973 12955 8007
rect 12897 7967 12955 7973
rect 13081 8007 13139 8013
rect 13081 7973 13093 8007
rect 13127 8004 13139 8007
rect 13814 8004 13820 8016
rect 13127 7976 13820 8004
rect 13127 7973 13139 7976
rect 13081 7967 13139 7973
rect 13814 7964 13820 7976
rect 13872 7964 13878 8016
rect 16850 7964 16856 8016
rect 16908 8004 16914 8016
rect 17681 8007 17739 8013
rect 17681 8004 17693 8007
rect 16908 7976 17693 8004
rect 16908 7964 16914 7976
rect 17681 7973 17693 7976
rect 17727 7973 17739 8007
rect 17681 7967 17739 7973
rect 17954 7964 17960 8016
rect 18012 8004 18018 8016
rect 25148 8004 25176 8044
rect 18012 7976 25176 8004
rect 25608 8004 25636 8044
rect 25682 8032 25688 8084
rect 25740 8072 25746 8084
rect 25777 8075 25835 8081
rect 25777 8072 25789 8075
rect 25740 8044 25789 8072
rect 25740 8032 25746 8044
rect 25777 8041 25789 8044
rect 25823 8041 25835 8075
rect 25777 8035 25835 8041
rect 28721 8075 28779 8081
rect 28721 8041 28733 8075
rect 28767 8072 28779 8075
rect 29362 8072 29368 8084
rect 28767 8044 29368 8072
rect 28767 8041 28779 8044
rect 28721 8035 28779 8041
rect 29362 8032 29368 8044
rect 29420 8032 29426 8084
rect 31662 8072 31668 8084
rect 29472 8044 31668 8072
rect 27798 8004 27804 8016
rect 25608 7976 27804 8004
rect 18012 7964 18018 7976
rect 27798 7964 27804 7976
rect 27856 7964 27862 8016
rect 28350 7964 28356 8016
rect 28408 8004 28414 8016
rect 28610 8007 28668 8013
rect 28610 8004 28622 8007
rect 28408 7976 28622 8004
rect 28408 7964 28414 7976
rect 28610 7973 28622 7976
rect 28656 8004 28668 8007
rect 29472 8004 29500 8044
rect 31662 8032 31668 8044
rect 31720 8032 31726 8084
rect 32858 8032 32864 8084
rect 32916 8072 32922 8084
rect 33962 8072 33968 8084
rect 32916 8044 33968 8072
rect 32916 8032 32922 8044
rect 33962 8032 33968 8044
rect 34020 8032 34026 8084
rect 34149 8075 34207 8081
rect 34149 8041 34161 8075
rect 34195 8072 34207 8075
rect 35802 8072 35808 8084
rect 34195 8044 35808 8072
rect 34195 8041 34207 8044
rect 34149 8035 34207 8041
rect 35802 8032 35808 8044
rect 35860 8032 35866 8084
rect 38657 8075 38715 8081
rect 35912 8044 37044 8072
rect 35912 8004 35940 8044
rect 28656 7976 29500 8004
rect 30116 7976 35940 8004
rect 37016 8004 37044 8044
rect 38657 8041 38669 8075
rect 38703 8072 38715 8075
rect 39206 8072 39212 8084
rect 38703 8044 39212 8072
rect 38703 8041 38715 8044
rect 38657 8035 38715 8041
rect 39206 8032 39212 8044
rect 39264 8032 39270 8084
rect 42705 8075 42763 8081
rect 42705 8041 42717 8075
rect 42751 8072 42763 8075
rect 43714 8072 43720 8084
rect 42751 8044 43720 8072
rect 42751 8041 42763 8044
rect 42705 8035 42763 8041
rect 43714 8032 43720 8044
rect 43772 8032 43778 8084
rect 44269 8075 44327 8081
rect 44269 8072 44281 8075
rect 43824 8044 44281 8072
rect 39942 8004 39948 8016
rect 37016 7976 39948 8004
rect 28656 7973 28668 7976
rect 28610 7967 28668 7973
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7936 8631 7939
rect 8938 7936 8944 7948
rect 8619 7908 8944 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 8938 7896 8944 7908
rect 8996 7896 9002 7948
rect 12618 7896 12624 7948
rect 12676 7896 12682 7948
rect 14734 7896 14740 7948
rect 14792 7936 14798 7948
rect 15102 7936 15108 7948
rect 14792 7908 15108 7936
rect 14792 7896 14798 7908
rect 15102 7896 15108 7908
rect 15160 7936 15166 7948
rect 15565 7939 15623 7945
rect 15565 7936 15577 7939
rect 15160 7908 15577 7936
rect 15160 7896 15166 7908
rect 15565 7905 15577 7908
rect 15611 7905 15623 7939
rect 15565 7899 15623 7905
rect 19058 7896 19064 7948
rect 19116 7936 19122 7948
rect 20438 7936 20444 7948
rect 19116 7908 20444 7936
rect 19116 7896 19122 7908
rect 20438 7896 20444 7908
rect 20496 7936 20502 7948
rect 23293 7939 23351 7945
rect 20496 7908 23152 7936
rect 20496 7896 20502 7908
rect 1578 7828 1584 7880
rect 1636 7828 1642 7880
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7156 7840 7849 7868
rect 7156 7828 7162 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 7926 7828 7932 7880
rect 7984 7828 7990 7880
rect 8113 7871 8171 7877
rect 8113 7837 8125 7871
rect 8159 7868 8171 7871
rect 8754 7868 8760 7880
rect 8159 7840 8760 7868
rect 8159 7837 8171 7840
rect 8113 7831 8171 7837
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7868 10103 7871
rect 10134 7868 10140 7880
rect 10091 7840 10140 7868
rect 10091 7837 10103 7840
rect 10045 7831 10103 7837
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7868 11023 7871
rect 11011 7840 15240 7868
rect 11011 7837 11023 7840
rect 10965 7831 11023 7837
rect 934 7760 940 7812
rect 992 7800 998 7812
rect 1857 7803 1915 7809
rect 1857 7800 1869 7803
rect 992 7772 1869 7800
rect 992 7760 998 7772
rect 1857 7769 1869 7772
rect 1903 7769 1915 7803
rect 1857 7763 1915 7769
rect 2682 7760 2688 7812
rect 2740 7800 2746 7812
rect 2740 7760 2774 7800
rect 9858 7760 9864 7812
rect 9916 7760 9922 7812
rect 10321 7803 10379 7809
rect 10321 7800 10333 7803
rect 9968 7772 10333 7800
rect 2746 7732 2774 7760
rect 9968 7732 9996 7772
rect 10321 7769 10333 7772
rect 10367 7800 10379 7803
rect 11977 7803 12035 7809
rect 11977 7800 11989 7803
rect 10367 7772 11989 7800
rect 10367 7769 10379 7772
rect 10321 7763 10379 7769
rect 11977 7769 11989 7772
rect 12023 7800 12035 7803
rect 12526 7800 12532 7812
rect 12023 7772 12532 7800
rect 12023 7769 12035 7772
rect 11977 7763 12035 7769
rect 12526 7760 12532 7772
rect 12584 7760 12590 7812
rect 2746 7704 9996 7732
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10229 7735 10287 7741
rect 10229 7732 10241 7735
rect 10100 7704 10241 7732
rect 10100 7692 10106 7704
rect 10229 7701 10241 7704
rect 10275 7701 10287 7735
rect 15212 7732 15240 7840
rect 15286 7828 15292 7880
rect 15344 7828 15350 7880
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7868 15715 7871
rect 15838 7868 15844 7880
rect 15703 7840 15844 7868
rect 15703 7837 15715 7840
rect 15657 7831 15715 7837
rect 15838 7828 15844 7840
rect 15896 7868 15902 7880
rect 16114 7868 16120 7880
rect 15896 7840 16120 7868
rect 15896 7828 15902 7840
rect 16114 7828 16120 7840
rect 16172 7868 16178 7880
rect 16577 7871 16635 7877
rect 16577 7868 16589 7871
rect 16172 7840 16589 7868
rect 16172 7828 16178 7840
rect 16577 7837 16589 7840
rect 16623 7837 16635 7871
rect 16577 7831 16635 7837
rect 16942 7828 16948 7880
rect 17000 7868 17006 7880
rect 17129 7871 17187 7877
rect 17129 7868 17141 7871
rect 17000 7840 17141 7868
rect 17000 7828 17006 7840
rect 17129 7837 17141 7840
rect 17175 7837 17187 7871
rect 17129 7831 17187 7837
rect 15562 7760 15568 7812
rect 15620 7800 15626 7812
rect 15749 7803 15807 7809
rect 15749 7800 15761 7803
rect 15620 7772 15761 7800
rect 15620 7760 15626 7772
rect 15749 7769 15761 7772
rect 15795 7800 15807 7803
rect 17144 7800 17172 7831
rect 17494 7828 17500 7880
rect 17552 7828 17558 7880
rect 18046 7828 18052 7880
rect 18104 7828 18110 7880
rect 18506 7828 18512 7880
rect 18564 7868 18570 7880
rect 19521 7871 19579 7877
rect 19521 7868 19533 7871
rect 18564 7840 19533 7868
rect 18564 7828 18570 7840
rect 19521 7837 19533 7840
rect 19567 7868 19579 7871
rect 22922 7868 22928 7880
rect 19567 7840 22928 7868
rect 19567 7837 19579 7840
rect 19521 7831 19579 7837
rect 22922 7828 22928 7840
rect 22980 7828 22986 7880
rect 23124 7868 23152 7908
rect 23293 7905 23305 7939
rect 23339 7936 23351 7939
rect 23474 7936 23480 7948
rect 23339 7908 23480 7936
rect 23339 7905 23351 7908
rect 23293 7899 23351 7905
rect 23474 7896 23480 7908
rect 23532 7896 23538 7948
rect 24302 7896 24308 7948
rect 24360 7936 24366 7948
rect 24949 7939 25007 7945
rect 24949 7936 24961 7939
rect 24360 7908 24961 7936
rect 24360 7896 24366 7908
rect 24949 7905 24961 7908
rect 24995 7905 25007 7939
rect 24949 7899 25007 7905
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 23124 7840 24593 7868
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 17862 7800 17868 7812
rect 15795 7772 17868 7800
rect 15795 7769 15807 7772
rect 15749 7763 15807 7769
rect 17862 7760 17868 7772
rect 17920 7760 17926 7812
rect 18414 7760 18420 7812
rect 18472 7800 18478 7812
rect 19889 7803 19947 7809
rect 19889 7800 19901 7803
rect 18472 7772 19901 7800
rect 18472 7760 18478 7772
rect 19889 7769 19901 7772
rect 19935 7769 19947 7803
rect 24118 7800 24124 7812
rect 19889 7763 19947 7769
rect 22066 7772 24124 7800
rect 16482 7732 16488 7744
rect 15212 7704 16488 7732
rect 10229 7695 10287 7701
rect 16482 7692 16488 7704
rect 16540 7692 16546 7744
rect 17034 7692 17040 7744
rect 17092 7732 17098 7744
rect 22066 7732 22094 7772
rect 24118 7760 24124 7772
rect 24176 7760 24182 7812
rect 24964 7800 24992 7899
rect 25038 7896 25044 7948
rect 25096 7936 25102 7948
rect 27430 7936 27436 7948
rect 25096 7908 27436 7936
rect 25096 7896 25102 7908
rect 27430 7896 27436 7908
rect 27488 7896 27494 7948
rect 27816 7936 27844 7964
rect 28813 7939 28871 7945
rect 27816 7908 28396 7936
rect 25593 7871 25651 7877
rect 25593 7837 25605 7871
rect 25639 7868 25651 7871
rect 26418 7868 26424 7880
rect 25639 7840 26424 7868
rect 25639 7837 25651 7840
rect 25593 7831 25651 7837
rect 26418 7828 26424 7840
rect 26476 7828 26482 7880
rect 26694 7828 26700 7880
rect 26752 7828 26758 7880
rect 28368 7868 28396 7908
rect 28813 7905 28825 7939
rect 28859 7936 28871 7939
rect 29178 7936 29184 7948
rect 28859 7908 29184 7936
rect 28859 7905 28871 7908
rect 28813 7899 28871 7905
rect 29178 7896 29184 7908
rect 29236 7896 29242 7948
rect 29270 7896 29276 7948
rect 29328 7936 29334 7948
rect 29328 7908 29868 7936
rect 29328 7896 29334 7908
rect 28368 7840 29684 7868
rect 26602 7800 26608 7812
rect 24964 7772 26608 7800
rect 26602 7760 26608 7772
rect 26660 7760 26666 7812
rect 27525 7803 27583 7809
rect 27525 7769 27537 7803
rect 27571 7769 27583 7803
rect 27525 7763 27583 7769
rect 17092 7704 22094 7732
rect 17092 7692 17098 7704
rect 22646 7692 22652 7744
rect 22704 7692 22710 7744
rect 22922 7692 22928 7744
rect 22980 7732 22986 7744
rect 23017 7735 23075 7741
rect 23017 7732 23029 7735
rect 22980 7704 23029 7732
rect 22980 7692 22986 7704
rect 23017 7701 23029 7704
rect 23063 7701 23075 7735
rect 23017 7695 23075 7701
rect 23106 7692 23112 7744
rect 23164 7692 23170 7744
rect 24762 7692 24768 7744
rect 24820 7692 24826 7744
rect 27154 7692 27160 7744
rect 27212 7732 27218 7744
rect 27540 7732 27568 7763
rect 27890 7760 27896 7812
rect 27948 7800 27954 7812
rect 28445 7803 28503 7809
rect 28445 7800 28457 7803
rect 27948 7772 28457 7800
rect 27948 7760 27954 7772
rect 28445 7769 28457 7772
rect 28491 7800 28503 7803
rect 29270 7800 29276 7812
rect 28491 7772 29276 7800
rect 28491 7769 28503 7772
rect 28445 7763 28503 7769
rect 29270 7760 29276 7772
rect 29328 7760 29334 7812
rect 27212 7704 27568 7732
rect 27212 7692 27218 7704
rect 29086 7692 29092 7744
rect 29144 7692 29150 7744
rect 29656 7732 29684 7840
rect 29840 7800 29868 7908
rect 30006 7828 30012 7880
rect 30064 7828 30070 7880
rect 30116 7877 30144 7976
rect 39942 7964 39948 7976
rect 40000 7964 40006 8016
rect 40034 7964 40040 8016
rect 40092 8004 40098 8016
rect 43824 8004 43852 8044
rect 44269 8041 44281 8044
rect 44315 8041 44327 8075
rect 44269 8035 44327 8041
rect 45373 8075 45431 8081
rect 45373 8041 45385 8075
rect 45419 8072 45431 8075
rect 46382 8072 46388 8084
rect 45419 8044 46388 8072
rect 45419 8041 45431 8044
rect 45373 8035 45431 8041
rect 46382 8032 46388 8044
rect 46440 8032 46446 8084
rect 56778 8072 56784 8084
rect 55508 8044 56784 8072
rect 40092 7976 43852 8004
rect 40092 7964 40098 7976
rect 30193 7939 30251 7945
rect 30193 7905 30205 7939
rect 30239 7936 30251 7939
rect 30282 7936 30288 7948
rect 30239 7908 30288 7936
rect 30239 7905 30251 7908
rect 30193 7899 30251 7905
rect 30282 7896 30288 7908
rect 30340 7896 30346 7948
rect 30466 7896 30472 7948
rect 30524 7936 30530 7948
rect 30929 7939 30987 7945
rect 30929 7936 30941 7939
rect 30524 7908 30941 7936
rect 30524 7896 30530 7908
rect 30929 7905 30941 7908
rect 30975 7905 30987 7939
rect 31481 7939 31539 7945
rect 31481 7936 31493 7939
rect 30929 7899 30987 7905
rect 31036 7908 31493 7936
rect 30101 7871 30159 7877
rect 30101 7837 30113 7871
rect 30147 7837 30159 7871
rect 31036 7868 31064 7908
rect 31481 7905 31493 7908
rect 31527 7905 31539 7939
rect 31481 7899 31539 7905
rect 32677 7939 32735 7945
rect 32677 7905 32689 7939
rect 32723 7936 32735 7939
rect 39022 7936 39028 7948
rect 32723 7908 36216 7936
rect 32723 7905 32735 7908
rect 32677 7899 32735 7905
rect 30101 7831 30159 7837
rect 30208 7840 31064 7868
rect 31389 7871 31447 7877
rect 30208 7800 30236 7840
rect 31389 7837 31401 7871
rect 31435 7837 31447 7871
rect 31389 7831 31447 7837
rect 29840 7772 30236 7800
rect 30466 7760 30472 7812
rect 30524 7760 30530 7812
rect 31404 7732 31432 7831
rect 31662 7828 31668 7880
rect 31720 7828 31726 7880
rect 32861 7871 32919 7877
rect 32861 7837 32873 7871
rect 32907 7868 32919 7871
rect 33226 7868 33232 7880
rect 32907 7840 33232 7868
rect 32907 7837 32919 7840
rect 32861 7831 32919 7837
rect 33226 7828 33232 7840
rect 33284 7828 33290 7880
rect 33410 7828 33416 7880
rect 33468 7868 33474 7880
rect 34149 7871 34207 7877
rect 34149 7868 34161 7871
rect 33468 7840 34161 7868
rect 33468 7828 33474 7840
rect 34149 7837 34161 7840
rect 34195 7837 34207 7871
rect 34149 7831 34207 7837
rect 34333 7871 34391 7877
rect 34333 7837 34345 7871
rect 34379 7837 34391 7871
rect 34333 7831 34391 7837
rect 34977 7871 35035 7877
rect 34977 7837 34989 7871
rect 35023 7868 35035 7871
rect 35342 7868 35348 7880
rect 35023 7840 35348 7868
rect 35023 7837 35035 7840
rect 34977 7831 35035 7837
rect 33134 7760 33140 7812
rect 33192 7760 33198 7812
rect 34348 7800 34376 7831
rect 35342 7828 35348 7840
rect 35400 7828 35406 7880
rect 36078 7828 36084 7880
rect 36136 7828 36142 7880
rect 36188 7800 36216 7908
rect 38028 7908 39028 7936
rect 36348 7871 36406 7877
rect 36348 7837 36360 7871
rect 36394 7868 36406 7871
rect 36906 7868 36912 7880
rect 36394 7840 36912 7868
rect 36394 7837 36406 7840
rect 36348 7831 36406 7837
rect 36906 7828 36912 7840
rect 36964 7828 36970 7880
rect 38028 7877 38056 7908
rect 39022 7896 39028 7908
rect 39080 7896 39086 7948
rect 43898 7896 43904 7948
rect 43956 7936 43962 7948
rect 43956 7908 44128 7936
rect 43956 7896 43962 7908
rect 38013 7871 38071 7877
rect 38013 7837 38025 7871
rect 38059 7837 38071 7871
rect 38013 7831 38071 7837
rect 38102 7828 38108 7880
rect 38160 7828 38166 7880
rect 38194 7828 38200 7880
rect 38252 7868 38258 7880
rect 38381 7871 38439 7877
rect 38381 7868 38393 7871
rect 38252 7840 38393 7868
rect 38252 7828 38258 7840
rect 38381 7837 38393 7840
rect 38427 7837 38439 7871
rect 38381 7831 38439 7837
rect 38478 7871 38536 7877
rect 38478 7837 38490 7871
rect 38524 7837 38536 7871
rect 38478 7831 38536 7837
rect 42613 7871 42671 7877
rect 42613 7837 42625 7871
rect 42659 7868 42671 7871
rect 42702 7868 42708 7880
rect 42659 7840 42708 7868
rect 42659 7837 42671 7840
rect 42613 7831 42671 7837
rect 36998 7800 37004 7812
rect 34348 7772 35204 7800
rect 36188 7772 37004 7800
rect 29656 7704 31432 7732
rect 31662 7692 31668 7744
rect 31720 7732 31726 7744
rect 31849 7735 31907 7741
rect 31849 7732 31861 7735
rect 31720 7704 31861 7732
rect 31720 7692 31726 7704
rect 31849 7701 31861 7704
rect 31895 7701 31907 7735
rect 31849 7695 31907 7701
rect 33042 7692 33048 7744
rect 33100 7692 33106 7744
rect 34514 7692 34520 7744
rect 34572 7732 34578 7744
rect 35069 7735 35127 7741
rect 35069 7732 35081 7735
rect 34572 7704 35081 7732
rect 34572 7692 34578 7704
rect 35069 7701 35081 7704
rect 35115 7701 35127 7735
rect 35176 7732 35204 7772
rect 36998 7760 37004 7772
rect 37056 7760 37062 7812
rect 37550 7760 37556 7812
rect 37608 7800 37614 7812
rect 38286 7800 38292 7812
rect 37608 7772 38292 7800
rect 37608 7760 37614 7772
rect 38286 7760 38292 7772
rect 38344 7760 38350 7812
rect 38493 7800 38521 7831
rect 42702 7828 42708 7840
rect 42760 7828 42766 7880
rect 43622 7828 43628 7880
rect 43680 7868 43686 7880
rect 43809 7871 43867 7877
rect 43809 7868 43821 7871
rect 43680 7840 43821 7868
rect 43680 7828 43686 7840
rect 43809 7837 43821 7840
rect 43855 7837 43867 7871
rect 43809 7831 43867 7837
rect 43990 7828 43996 7880
rect 44048 7828 44054 7880
rect 44100 7877 44128 7908
rect 46474 7896 46480 7948
rect 46532 7936 46538 7948
rect 46569 7939 46627 7945
rect 46569 7936 46581 7939
rect 46532 7908 46581 7936
rect 46532 7896 46538 7908
rect 46569 7905 46581 7908
rect 46615 7905 46627 7939
rect 46569 7899 46627 7905
rect 44085 7871 44143 7877
rect 44085 7837 44097 7871
rect 44131 7837 44143 7871
rect 44085 7831 44143 7837
rect 44726 7828 44732 7880
rect 44784 7868 44790 7880
rect 45557 7871 45615 7877
rect 45557 7868 45569 7871
rect 44784 7840 45569 7868
rect 44784 7828 44790 7840
rect 45557 7837 45569 7840
rect 45603 7837 45615 7871
rect 45557 7831 45615 7837
rect 46106 7828 46112 7880
rect 46164 7868 46170 7880
rect 55508 7877 55536 8044
rect 56778 8032 56784 8044
rect 56836 8032 56842 8084
rect 56137 8007 56195 8013
rect 56137 7973 56149 8007
rect 56183 8004 56195 8007
rect 56183 7976 56824 8004
rect 56183 7973 56195 7976
rect 56137 7967 56195 7973
rect 55600 7908 56456 7936
rect 46293 7871 46351 7877
rect 46293 7868 46305 7871
rect 46164 7840 46305 7868
rect 46164 7828 46170 7840
rect 46293 7837 46305 7840
rect 46339 7837 46351 7871
rect 46293 7831 46351 7837
rect 55493 7871 55551 7877
rect 55493 7837 55505 7871
rect 55539 7837 55551 7871
rect 55493 7831 55551 7837
rect 38396 7772 38521 7800
rect 38396 7744 38424 7772
rect 45094 7760 45100 7812
rect 45152 7800 45158 7812
rect 45281 7803 45339 7809
rect 45281 7800 45293 7803
rect 45152 7772 45293 7800
rect 45152 7760 45158 7772
rect 45281 7769 45293 7772
rect 45327 7769 45339 7803
rect 45281 7763 45339 7769
rect 45465 7803 45523 7809
rect 45465 7769 45477 7803
rect 45511 7800 45523 7803
rect 46566 7800 46572 7812
rect 45511 7772 46572 7800
rect 45511 7769 45523 7772
rect 45465 7763 45523 7769
rect 46566 7760 46572 7772
rect 46624 7760 46630 7812
rect 52270 7760 52276 7812
rect 52328 7800 52334 7812
rect 55600 7800 55628 7908
rect 56428 7877 56456 7908
rect 55677 7871 55735 7877
rect 55677 7837 55689 7871
rect 55723 7868 55735 7871
rect 56413 7871 56471 7877
rect 55723 7840 56364 7868
rect 55723 7837 55735 7840
rect 55677 7831 55735 7837
rect 52328 7772 55628 7800
rect 52328 7760 52334 7772
rect 55766 7760 55772 7812
rect 55824 7800 55830 7812
rect 56134 7800 56140 7812
rect 55824 7772 56140 7800
rect 55824 7760 55830 7772
rect 56134 7760 56140 7772
rect 56192 7760 56198 7812
rect 56336 7800 56364 7840
rect 56413 7837 56425 7871
rect 56459 7837 56471 7871
rect 56796 7868 56824 7976
rect 56870 7896 56876 7948
rect 56928 7896 56934 7948
rect 57129 7871 57187 7877
rect 57129 7868 57141 7871
rect 56796 7840 57141 7868
rect 56413 7831 56471 7837
rect 57129 7837 57141 7840
rect 57175 7837 57187 7871
rect 57129 7831 57187 7837
rect 57882 7800 57888 7812
rect 56336 7772 57888 7800
rect 57882 7760 57888 7772
rect 57940 7800 57946 7812
rect 57940 7772 58296 7800
rect 57940 7760 57946 7772
rect 36354 7732 36360 7744
rect 35176 7704 36360 7732
rect 35069 7695 35127 7701
rect 36354 7692 36360 7704
rect 36412 7692 36418 7744
rect 36538 7692 36544 7744
rect 36596 7732 36602 7744
rect 37461 7735 37519 7741
rect 37461 7732 37473 7735
rect 36596 7704 37473 7732
rect 36596 7692 36602 7704
rect 37461 7701 37473 7704
rect 37507 7701 37519 7735
rect 37461 7695 37519 7701
rect 38378 7692 38384 7744
rect 38436 7692 38442 7744
rect 40770 7692 40776 7744
rect 40828 7732 40834 7744
rect 49418 7732 49424 7744
rect 40828 7704 49424 7732
rect 40828 7692 40834 7704
rect 49418 7692 49424 7704
rect 49476 7692 49482 7744
rect 58268 7741 58296 7772
rect 55677 7735 55735 7741
rect 55677 7701 55689 7735
rect 55723 7732 55735 7735
rect 56321 7735 56379 7741
rect 56321 7732 56333 7735
rect 55723 7704 56333 7732
rect 55723 7701 55735 7704
rect 55677 7695 55735 7701
rect 56321 7701 56333 7704
rect 56367 7701 56379 7735
rect 56321 7695 56379 7701
rect 58253 7735 58311 7741
rect 58253 7701 58265 7735
rect 58299 7701 58311 7735
rect 58253 7695 58311 7701
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 10594 7488 10600 7540
rect 10652 7488 10658 7540
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 11020 7500 12434 7528
rect 11020 7488 11026 7500
rect 8754 7420 8760 7472
rect 8812 7460 8818 7472
rect 11977 7463 12035 7469
rect 11977 7460 11989 7463
rect 8812 7432 11008 7460
rect 8812 7420 8818 7432
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 10686 7392 10692 7404
rect 1636 7364 10692 7392
rect 1636 7352 1642 7364
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 10778 7352 10784 7404
rect 10836 7352 10842 7404
rect 10980 7401 11008 7432
rect 11348 7432 11989 7460
rect 11348 7404 11376 7432
rect 11977 7429 11989 7432
rect 12023 7429 12035 7463
rect 12406 7460 12434 7500
rect 12526 7488 12532 7540
rect 12584 7528 12590 7540
rect 17034 7528 17040 7540
rect 12584 7500 17040 7528
rect 12584 7488 12590 7500
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 17494 7488 17500 7540
rect 17552 7528 17558 7540
rect 18601 7531 18659 7537
rect 18601 7528 18613 7531
rect 17552 7500 18613 7528
rect 17552 7488 17558 7500
rect 18601 7497 18613 7500
rect 18647 7497 18659 7531
rect 18601 7491 18659 7497
rect 20346 7488 20352 7540
rect 20404 7528 20410 7540
rect 22189 7531 22247 7537
rect 22189 7528 22201 7531
rect 20404 7500 22201 7528
rect 20404 7488 20410 7500
rect 22189 7497 22201 7500
rect 22235 7497 22247 7531
rect 22189 7491 22247 7497
rect 24394 7488 24400 7540
rect 24452 7528 24458 7540
rect 24673 7531 24731 7537
rect 24673 7528 24685 7531
rect 24452 7500 24685 7528
rect 24452 7488 24458 7500
rect 24673 7497 24685 7500
rect 24719 7497 24731 7531
rect 24673 7491 24731 7497
rect 24854 7488 24860 7540
rect 24912 7528 24918 7540
rect 25130 7528 25136 7540
rect 24912 7500 25136 7528
rect 24912 7488 24918 7500
rect 25130 7488 25136 7500
rect 25188 7528 25194 7540
rect 25961 7531 26019 7537
rect 25961 7528 25973 7531
rect 25188 7500 25973 7528
rect 25188 7488 25194 7500
rect 25961 7497 25973 7500
rect 26007 7497 26019 7531
rect 25961 7491 26019 7497
rect 28534 7488 28540 7540
rect 28592 7528 28598 7540
rect 29917 7531 29975 7537
rect 29917 7528 29929 7531
rect 28592 7500 29929 7528
rect 28592 7488 28598 7500
rect 29917 7497 29929 7500
rect 29963 7497 29975 7531
rect 29917 7491 29975 7497
rect 12406 7432 15056 7460
rect 11977 7423 12035 7429
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7392 11023 7395
rect 11330 7392 11336 7404
rect 11011 7364 11336 7392
rect 11011 7361 11023 7364
rect 10965 7355 11023 7361
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7392 11851 7395
rect 12437 7395 12495 7401
rect 12437 7392 12449 7395
rect 11839 7364 12449 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 12437 7361 12449 7364
rect 12483 7392 12495 7395
rect 12618 7392 12624 7404
rect 12483 7364 12624 7392
rect 12483 7361 12495 7364
rect 12437 7355 12495 7361
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 10870 7284 10876 7336
rect 10928 7284 10934 7336
rect 11054 7284 11060 7336
rect 11112 7284 11118 7336
rect 12894 7284 12900 7336
rect 12952 7284 12958 7336
rect 9858 7216 9864 7268
rect 9916 7256 9922 7268
rect 10962 7256 10968 7268
rect 9916 7228 10968 7256
rect 9916 7216 9922 7228
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 12713 7259 12771 7265
rect 12713 7225 12725 7259
rect 12759 7225 12771 7259
rect 12713 7219 12771 7225
rect 7374 7148 7380 7200
rect 7432 7188 7438 7200
rect 12728 7188 12756 7219
rect 7432 7160 12756 7188
rect 15028 7188 15056 7432
rect 15102 7420 15108 7472
rect 15160 7420 15166 7472
rect 15194 7420 15200 7472
rect 15252 7420 15258 7472
rect 15657 7463 15715 7469
rect 15657 7429 15669 7463
rect 15703 7460 15715 7463
rect 15838 7460 15844 7472
rect 15703 7432 15844 7460
rect 15703 7429 15715 7432
rect 15657 7423 15715 7429
rect 15838 7420 15844 7432
rect 15896 7460 15902 7472
rect 15896 7432 16620 7460
rect 15896 7420 15902 7432
rect 15562 7352 15568 7404
rect 15620 7352 15626 7404
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7361 16175 7395
rect 16592 7392 16620 7432
rect 16666 7420 16672 7472
rect 16724 7460 16730 7472
rect 16850 7460 16856 7472
rect 16724 7432 16856 7460
rect 16724 7420 16730 7432
rect 16850 7420 16856 7432
rect 16908 7420 16914 7472
rect 16942 7420 16948 7472
rect 17000 7460 17006 7472
rect 17512 7460 17540 7488
rect 17000 7432 17540 7460
rect 17000 7420 17006 7432
rect 18506 7420 18512 7472
rect 18564 7420 18570 7472
rect 22922 7420 22928 7472
rect 22980 7460 22986 7472
rect 23566 7460 23572 7472
rect 22980 7432 23572 7460
rect 22980 7420 22986 7432
rect 23566 7420 23572 7432
rect 23624 7460 23630 7472
rect 25498 7460 25504 7472
rect 23624 7432 25504 7460
rect 23624 7420 23630 7432
rect 25498 7420 25504 7432
rect 25556 7420 25562 7472
rect 28626 7460 28632 7472
rect 27540 7432 28632 7460
rect 17310 7392 17316 7404
rect 16592 7364 17316 7392
rect 16117 7355 16175 7361
rect 15286 7284 15292 7336
rect 15344 7324 15350 7336
rect 15838 7324 15844 7336
rect 15344 7296 15844 7324
rect 15344 7284 15350 7296
rect 15838 7284 15844 7296
rect 15896 7324 15902 7336
rect 16132 7324 16160 7355
rect 17310 7352 17316 7364
rect 17368 7392 17374 7404
rect 17405 7395 17463 7401
rect 17405 7392 17417 7395
rect 17368 7364 17417 7392
rect 17368 7352 17374 7364
rect 17405 7361 17417 7364
rect 17451 7361 17463 7395
rect 17405 7355 17463 7361
rect 17494 7352 17500 7404
rect 17552 7352 17558 7404
rect 20340 7395 20398 7401
rect 20340 7361 20352 7395
rect 20386 7392 20398 7395
rect 20622 7392 20628 7404
rect 20386 7364 20628 7392
rect 20386 7361 20398 7364
rect 20340 7355 20398 7361
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 22002 7352 22008 7404
rect 22060 7401 22066 7404
rect 22060 7355 22069 7401
rect 23385 7395 23443 7401
rect 23385 7361 23397 7395
rect 23431 7392 23443 7395
rect 27540 7392 27568 7432
rect 28626 7420 28632 7432
rect 28684 7420 28690 7472
rect 29932 7460 29960 7491
rect 30006 7488 30012 7540
rect 30064 7528 30070 7540
rect 35526 7528 35532 7540
rect 30064 7500 35532 7528
rect 30064 7488 30070 7500
rect 35526 7488 35532 7500
rect 35584 7488 35590 7540
rect 36173 7531 36231 7537
rect 36173 7497 36185 7531
rect 36219 7528 36231 7531
rect 36722 7528 36728 7540
rect 36219 7500 36728 7528
rect 36219 7497 36231 7500
rect 36173 7491 36231 7497
rect 36722 7488 36728 7500
rect 36780 7488 36786 7540
rect 37553 7531 37611 7537
rect 37553 7497 37565 7531
rect 37599 7528 37611 7531
rect 38102 7528 38108 7540
rect 37599 7500 38108 7528
rect 37599 7497 37611 7500
rect 37553 7491 37611 7497
rect 38102 7488 38108 7500
rect 38160 7488 38166 7540
rect 41386 7500 56088 7528
rect 31294 7460 31300 7472
rect 29932 7432 31300 7460
rect 31294 7420 31300 7432
rect 31352 7460 31358 7472
rect 36078 7460 36084 7472
rect 31352 7432 31754 7460
rect 31352 7420 31358 7432
rect 23431 7364 27568 7392
rect 27617 7395 27675 7401
rect 23431 7361 23443 7364
rect 23385 7355 23443 7361
rect 27617 7361 27629 7395
rect 27663 7392 27675 7395
rect 29086 7392 29092 7404
rect 27663 7364 29092 7392
rect 27663 7361 27675 7364
rect 27617 7355 27675 7361
rect 22060 7352 22066 7355
rect 29086 7352 29092 7364
rect 29144 7352 29150 7404
rect 31018 7352 31024 7404
rect 31076 7392 31082 7404
rect 31205 7395 31263 7401
rect 31205 7392 31217 7395
rect 31076 7364 31217 7392
rect 31076 7352 31082 7364
rect 31205 7361 31217 7364
rect 31251 7361 31263 7395
rect 31205 7355 31263 7361
rect 15896 7296 16160 7324
rect 17037 7327 17095 7333
rect 15896 7284 15902 7296
rect 17037 7293 17049 7327
rect 17083 7324 17095 7327
rect 17586 7324 17592 7336
rect 17083 7296 17592 7324
rect 17083 7293 17095 7296
rect 17037 7287 17095 7293
rect 17586 7284 17592 7296
rect 17644 7284 17650 7336
rect 17862 7284 17868 7336
rect 17920 7324 17926 7336
rect 17957 7327 18015 7333
rect 17957 7324 17969 7327
rect 17920 7296 17969 7324
rect 17920 7284 17926 7296
rect 17957 7293 17969 7296
rect 18003 7293 18015 7327
rect 17957 7287 18015 7293
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 20070 7324 20076 7336
rect 19484 7296 20076 7324
rect 19484 7284 19490 7296
rect 20070 7284 20076 7296
rect 20128 7284 20134 7336
rect 27706 7284 27712 7336
rect 27764 7284 27770 7336
rect 27982 7284 27988 7336
rect 28040 7284 28046 7336
rect 30650 7284 30656 7336
rect 30708 7324 30714 7336
rect 31297 7327 31355 7333
rect 31297 7324 31309 7327
rect 30708 7296 31309 7324
rect 30708 7284 30714 7296
rect 31297 7293 31309 7296
rect 31343 7293 31355 7327
rect 31297 7287 31355 7293
rect 31478 7284 31484 7336
rect 31536 7284 31542 7336
rect 31726 7324 31754 7432
rect 34164 7432 36084 7460
rect 34164 7333 34192 7432
rect 36078 7420 36084 7432
rect 36136 7420 36142 7472
rect 36538 7420 36544 7472
rect 36596 7420 36602 7472
rect 36998 7420 37004 7472
rect 37056 7460 37062 7472
rect 41386 7460 41414 7500
rect 37056 7432 41414 7460
rect 37056 7420 37062 7432
rect 44542 7420 44548 7472
rect 44600 7460 44606 7472
rect 46201 7463 46259 7469
rect 44600 7432 45232 7460
rect 44600 7420 44606 7432
rect 34422 7401 34428 7404
rect 34416 7355 34428 7401
rect 34422 7352 34428 7355
rect 34480 7352 34486 7404
rect 34790 7352 34796 7404
rect 34848 7392 34854 7404
rect 36633 7395 36691 7401
rect 36633 7392 36645 7395
rect 34848 7364 36645 7392
rect 34848 7352 34854 7364
rect 36633 7361 36645 7364
rect 36679 7392 36691 7395
rect 36722 7392 36728 7404
rect 36679 7364 36728 7392
rect 36679 7361 36691 7364
rect 36633 7355 36691 7361
rect 36722 7352 36728 7364
rect 36780 7352 36786 7404
rect 37461 7395 37519 7401
rect 37461 7361 37473 7395
rect 37507 7361 37519 7395
rect 37461 7355 37519 7361
rect 37645 7395 37703 7401
rect 37645 7361 37657 7395
rect 37691 7392 37703 7395
rect 38378 7392 38384 7404
rect 37691 7364 38384 7392
rect 37691 7361 37703 7364
rect 37645 7355 37703 7361
rect 34149 7327 34207 7333
rect 34149 7324 34161 7327
rect 31726 7296 34161 7324
rect 34149 7293 34161 7296
rect 34195 7293 34207 7327
rect 34149 7287 34207 7293
rect 36814 7284 36820 7336
rect 36872 7284 36878 7336
rect 25038 7256 25044 7268
rect 21008 7228 25044 7256
rect 21008 7188 21036 7228
rect 25038 7216 25044 7228
rect 25096 7216 25102 7268
rect 25130 7216 25136 7268
rect 25188 7256 25194 7268
rect 25406 7256 25412 7268
rect 25188 7228 25412 7256
rect 25188 7216 25194 7228
rect 25406 7216 25412 7228
rect 25464 7256 25470 7268
rect 25593 7259 25651 7265
rect 25593 7256 25605 7259
rect 25464 7228 25605 7256
rect 25464 7216 25470 7228
rect 25593 7225 25605 7228
rect 25639 7225 25651 7259
rect 28000 7256 28028 7284
rect 25593 7219 25651 7225
rect 27908 7228 28028 7256
rect 15028 7160 21036 7188
rect 7432 7148 7438 7160
rect 21450 7148 21456 7200
rect 21508 7148 21514 7200
rect 25498 7148 25504 7200
rect 25556 7188 25562 7200
rect 25961 7191 26019 7197
rect 25961 7188 25973 7191
rect 25556 7160 25973 7188
rect 25556 7148 25562 7160
rect 25961 7157 25973 7160
rect 26007 7157 26019 7191
rect 25961 7151 26019 7157
rect 26145 7191 26203 7197
rect 26145 7157 26157 7191
rect 26191 7188 26203 7191
rect 26510 7188 26516 7200
rect 26191 7160 26516 7188
rect 26191 7157 26203 7160
rect 26145 7151 26203 7157
rect 26510 7148 26516 7160
rect 26568 7148 26574 7200
rect 27801 7191 27859 7197
rect 27801 7157 27813 7191
rect 27847 7188 27859 7191
rect 27908 7188 27936 7228
rect 28258 7216 28264 7268
rect 28316 7256 28322 7268
rect 29730 7256 29736 7268
rect 28316 7228 29736 7256
rect 28316 7216 28322 7228
rect 29730 7216 29736 7228
rect 29788 7216 29794 7268
rect 29914 7216 29920 7268
rect 29972 7256 29978 7268
rect 37476 7256 37504 7355
rect 38378 7352 38384 7364
rect 38436 7352 38442 7404
rect 43990 7352 43996 7404
rect 44048 7392 44054 7404
rect 45204 7401 45232 7432
rect 46201 7429 46213 7463
rect 46247 7460 46259 7463
rect 54846 7460 54852 7472
rect 46247 7432 54852 7460
rect 46247 7429 46259 7432
rect 46201 7423 46259 7429
rect 54846 7420 54852 7432
rect 54904 7420 54910 7472
rect 55766 7420 55772 7472
rect 55824 7420 55830 7472
rect 44453 7395 44511 7401
rect 44453 7392 44465 7395
rect 44048 7364 44465 7392
rect 44048 7352 44054 7364
rect 44453 7361 44465 7364
rect 44499 7361 44511 7395
rect 44453 7355 44511 7361
rect 45189 7395 45247 7401
rect 45189 7361 45201 7395
rect 45235 7361 45247 7395
rect 45189 7355 45247 7361
rect 29972 7228 31754 7256
rect 29972 7216 29978 7228
rect 27847 7160 27936 7188
rect 27847 7157 27859 7160
rect 27801 7151 27859 7157
rect 27982 7148 27988 7200
rect 28040 7148 28046 7200
rect 29638 7148 29644 7200
rect 29696 7188 29702 7200
rect 30190 7188 30196 7200
rect 29696 7160 30196 7188
rect 29696 7148 29702 7160
rect 30190 7148 30196 7160
rect 30248 7148 30254 7200
rect 30837 7191 30895 7197
rect 30837 7157 30849 7191
rect 30883 7188 30895 7191
rect 31110 7188 31116 7200
rect 30883 7160 31116 7188
rect 30883 7157 30895 7160
rect 30837 7151 30895 7157
rect 31110 7148 31116 7160
rect 31168 7148 31174 7200
rect 31726 7188 31754 7228
rect 35084 7228 37504 7256
rect 44468 7256 44496 7355
rect 45370 7352 45376 7404
rect 45428 7352 45434 7404
rect 46290 7352 46296 7404
rect 46348 7352 46354 7404
rect 56060 7401 56088 7500
rect 56134 7420 56140 7472
rect 56192 7460 56198 7472
rect 56965 7463 57023 7469
rect 56965 7460 56977 7463
rect 56192 7432 56977 7460
rect 56192 7420 56198 7432
rect 56965 7429 56977 7432
rect 57011 7429 57023 7463
rect 56965 7423 57023 7429
rect 55953 7395 56011 7401
rect 55953 7361 55965 7395
rect 55999 7361 56011 7395
rect 55953 7355 56011 7361
rect 56045 7395 56103 7401
rect 56045 7361 56057 7395
rect 56091 7361 56103 7395
rect 56045 7355 56103 7361
rect 56597 7395 56655 7401
rect 56597 7361 56609 7395
rect 56643 7392 56655 7395
rect 56686 7392 56692 7404
rect 56643 7364 56692 7392
rect 56643 7361 56655 7364
rect 56597 7355 56655 7361
rect 45094 7284 45100 7336
rect 45152 7324 45158 7336
rect 45281 7327 45339 7333
rect 45281 7324 45293 7327
rect 45152 7296 45293 7324
rect 45152 7284 45158 7296
rect 45281 7293 45293 7296
rect 45327 7293 45339 7327
rect 45281 7287 45339 7293
rect 46474 7284 46480 7336
rect 46532 7284 46538 7336
rect 52270 7256 52276 7268
rect 44468 7228 52276 7256
rect 35084 7188 35112 7228
rect 52270 7216 52276 7228
rect 52328 7216 52334 7268
rect 55968 7256 55996 7355
rect 56686 7352 56692 7364
rect 56744 7352 56750 7404
rect 56778 7352 56784 7404
rect 56836 7392 56842 7404
rect 58069 7395 58127 7401
rect 58069 7392 58081 7395
rect 56836 7364 58081 7392
rect 56836 7352 56842 7364
rect 58069 7361 58081 7364
rect 58115 7361 58127 7395
rect 58069 7355 58127 7361
rect 58250 7352 58256 7404
rect 58308 7352 58314 7404
rect 58161 7259 58219 7265
rect 58161 7256 58173 7259
rect 55968 7228 58173 7256
rect 58161 7225 58173 7228
rect 58207 7225 58219 7259
rect 58161 7219 58219 7225
rect 31726 7160 35112 7188
rect 41506 7148 41512 7200
rect 41564 7188 41570 7200
rect 45462 7188 45468 7200
rect 41564 7160 45468 7188
rect 41564 7148 41570 7160
rect 45462 7148 45468 7160
rect 45520 7148 45526 7200
rect 45830 7148 45836 7200
rect 45888 7148 45894 7200
rect 55769 7191 55827 7197
rect 55769 7157 55781 7191
rect 55815 7188 55827 7191
rect 56962 7188 56968 7200
rect 55815 7160 56968 7188
rect 55815 7157 55827 7160
rect 55769 7151 55827 7157
rect 56962 7148 56968 7160
rect 57020 7148 57026 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 12676 6956 13645 6984
rect 12676 6944 12682 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 18966 6984 18972 6996
rect 13633 6947 13691 6953
rect 15028 6956 18972 6984
rect 10870 6876 10876 6928
rect 10928 6916 10934 6928
rect 15028 6916 15056 6956
rect 18966 6944 18972 6956
rect 19024 6944 19030 6996
rect 20070 6944 20076 6996
rect 20128 6984 20134 6996
rect 20128 6956 20208 6984
rect 20128 6944 20134 6956
rect 10928 6888 15056 6916
rect 10928 6876 10934 6888
rect 15102 6876 15108 6928
rect 15160 6916 15166 6928
rect 17494 6916 17500 6928
rect 15160 6888 17500 6916
rect 15160 6876 15166 6888
rect 934 6808 940 6860
rect 992 6848 998 6860
rect 1765 6851 1823 6857
rect 1765 6848 1777 6851
rect 992 6820 1777 6848
rect 992 6808 998 6820
rect 1765 6817 1777 6820
rect 1811 6817 1823 6851
rect 1765 6811 1823 6817
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 8812 6820 9536 6848
rect 8812 6808 8818 6820
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 9122 6780 9128 6792
rect 1627 6752 9128 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 9122 6740 9128 6752
rect 9180 6740 9186 6792
rect 9508 6789 9536 6820
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 10781 6851 10839 6857
rect 10781 6848 10793 6851
rect 10744 6820 10793 6848
rect 10744 6808 10750 6820
rect 10781 6817 10793 6820
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 11057 6851 11115 6857
rect 11057 6817 11069 6851
rect 11103 6848 11115 6851
rect 15746 6848 15752 6860
rect 11103 6820 15752 6848
rect 11103 6817 11115 6820
rect 11057 6811 11115 6817
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 16025 6851 16083 6857
rect 16025 6848 16037 6851
rect 15988 6820 16037 6848
rect 15988 6808 15994 6820
rect 16025 6817 16037 6820
rect 16071 6817 16083 6851
rect 16025 6811 16083 6817
rect 16117 6851 16175 6857
rect 16117 6817 16129 6851
rect 16163 6848 16175 6851
rect 16390 6848 16396 6860
rect 16163 6820 16396 6848
rect 16163 6817 16175 6820
rect 16117 6811 16175 6817
rect 16390 6808 16396 6820
rect 16448 6808 16454 6860
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 10870 6740 10876 6792
rect 10928 6780 10934 6792
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10928 6752 10977 6780
rect 10928 6740 10934 6752
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11149 6783 11207 6789
rect 11149 6749 11161 6783
rect 11195 6749 11207 6783
rect 11149 6743 11207 6749
rect 11164 6712 11192 6743
rect 11238 6740 11244 6792
rect 11296 6740 11302 6792
rect 16500 6789 16528 6888
rect 17494 6876 17500 6888
rect 17552 6876 17558 6928
rect 20180 6916 20208 6956
rect 20622 6944 20628 6996
rect 20680 6984 20686 6996
rect 20717 6987 20775 6993
rect 20717 6984 20729 6987
rect 20680 6956 20729 6984
rect 20680 6944 20686 6956
rect 20717 6953 20729 6956
rect 20763 6953 20775 6987
rect 23382 6984 23388 6996
rect 20717 6947 20775 6953
rect 22480 6956 23388 6984
rect 20254 6916 20260 6928
rect 19536 6888 20116 6916
rect 20180 6888 20260 6916
rect 17310 6808 17316 6860
rect 17368 6848 17374 6860
rect 17681 6851 17739 6857
rect 17681 6848 17693 6851
rect 17368 6820 17693 6848
rect 17368 6808 17374 6820
rect 17681 6817 17693 6820
rect 17727 6817 17739 6851
rect 17681 6811 17739 6817
rect 16592 6789 16712 6790
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6749 16543 6783
rect 16485 6743 16543 6749
rect 16577 6783 16712 6789
rect 16577 6749 16589 6783
rect 16623 6780 16712 6783
rect 16942 6780 16948 6792
rect 16623 6762 16948 6780
rect 16623 6749 16635 6762
rect 16684 6752 16948 6762
rect 16577 6743 16635 6749
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 17402 6740 17408 6792
rect 17460 6740 17466 6792
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 19536 6780 19564 6888
rect 19978 6848 19984 6860
rect 19628 6820 19984 6848
rect 19628 6789 19656 6820
rect 19978 6808 19984 6820
rect 20036 6808 20042 6860
rect 20088 6848 20116 6888
rect 20254 6876 20260 6888
rect 20312 6916 20318 6928
rect 22480 6916 22508 6956
rect 23382 6944 23388 6956
rect 23440 6984 23446 6996
rect 24394 6984 24400 6996
rect 23440 6956 24400 6984
rect 23440 6944 23446 6956
rect 24394 6944 24400 6956
rect 24452 6944 24458 6996
rect 24486 6944 24492 6996
rect 24544 6984 24550 6996
rect 24544 6956 27844 6984
rect 24544 6944 24550 6956
rect 27816 6916 27844 6956
rect 27890 6944 27896 6996
rect 27948 6984 27954 6996
rect 28123 6987 28181 6993
rect 28123 6984 28135 6987
rect 27948 6956 28135 6984
rect 27948 6944 27954 6956
rect 28123 6953 28135 6956
rect 28169 6953 28181 6987
rect 28123 6947 28181 6953
rect 28261 6987 28319 6993
rect 28261 6953 28273 6987
rect 28307 6984 28319 6987
rect 28350 6984 28356 6996
rect 28307 6956 28356 6984
rect 28307 6953 28319 6956
rect 28261 6947 28319 6953
rect 28350 6944 28356 6956
rect 28408 6944 28414 6996
rect 31662 6984 31668 6996
rect 30024 6956 31668 6984
rect 30024 6928 30052 6956
rect 31662 6944 31668 6956
rect 31720 6944 31726 6996
rect 34333 6987 34391 6993
rect 34333 6953 34345 6987
rect 34379 6984 34391 6987
rect 34422 6984 34428 6996
rect 34379 6956 34428 6984
rect 34379 6953 34391 6956
rect 34333 6947 34391 6953
rect 34422 6944 34428 6956
rect 34480 6944 34486 6996
rect 39022 6944 39028 6996
rect 39080 6984 39086 6996
rect 46106 6984 46112 6996
rect 39080 6956 46112 6984
rect 39080 6944 39086 6956
rect 46106 6944 46112 6956
rect 46164 6944 46170 6996
rect 46290 6944 46296 6996
rect 46348 6984 46354 6996
rect 46569 6987 46627 6993
rect 46569 6984 46581 6987
rect 46348 6956 46581 6984
rect 46348 6944 46354 6956
rect 46569 6953 46581 6956
rect 46615 6953 46627 6987
rect 46569 6947 46627 6953
rect 30006 6916 30012 6928
rect 20312 6888 22508 6916
rect 20312 6876 20318 6888
rect 21082 6848 21088 6860
rect 20088 6820 21088 6848
rect 21082 6808 21088 6820
rect 21140 6808 21146 6860
rect 21266 6808 21272 6860
rect 21324 6808 21330 6860
rect 22480 6857 22508 6888
rect 26436 6888 27292 6916
rect 27816 6888 30012 6916
rect 22465 6851 22523 6857
rect 22465 6817 22477 6851
rect 22511 6817 22523 6851
rect 22465 6811 22523 6817
rect 25409 6851 25467 6857
rect 25409 6817 25421 6851
rect 25455 6848 25467 6851
rect 26436 6848 26464 6888
rect 25455 6820 26464 6848
rect 25455 6817 25467 6820
rect 25409 6811 25467 6817
rect 26510 6808 26516 6860
rect 26568 6808 26574 6860
rect 27154 6848 27160 6860
rect 26620 6820 27160 6848
rect 17644 6752 19564 6780
rect 19613 6783 19671 6789
rect 17644 6740 17650 6752
rect 19613 6749 19625 6783
rect 19659 6749 19671 6783
rect 22732 6783 22790 6789
rect 22732 6780 22744 6783
rect 19613 6743 19671 6749
rect 22664 6752 22744 6780
rect 22664 6724 22692 6752
rect 22732 6749 22744 6752
rect 22778 6749 22790 6783
rect 22732 6743 22790 6749
rect 25961 6783 26019 6789
rect 25961 6749 25973 6783
rect 26007 6780 26019 6783
rect 26050 6780 26056 6792
rect 26007 6752 26056 6780
rect 26007 6749 26019 6752
rect 25961 6743 26019 6749
rect 26050 6740 26056 6752
rect 26108 6740 26114 6792
rect 26620 6789 26648 6820
rect 27154 6808 27160 6820
rect 27212 6808 27218 6860
rect 27264 6848 27292 6888
rect 30006 6876 30012 6888
rect 30064 6876 30070 6928
rect 30742 6876 30748 6928
rect 30800 6916 30806 6928
rect 31478 6916 31484 6928
rect 30800 6888 31484 6916
rect 30800 6876 30806 6888
rect 31478 6876 31484 6888
rect 31536 6916 31542 6928
rect 31536 6888 35572 6916
rect 31536 6876 31542 6888
rect 27614 6848 27620 6860
rect 27264 6820 27620 6848
rect 27614 6808 27620 6820
rect 27672 6808 27678 6860
rect 28074 6808 28080 6860
rect 28132 6848 28138 6860
rect 28353 6851 28411 6857
rect 28353 6848 28365 6851
rect 28132 6820 28365 6848
rect 28132 6808 28138 6820
rect 28353 6817 28365 6820
rect 28399 6817 28411 6851
rect 28353 6811 28411 6817
rect 28626 6808 28632 6860
rect 28684 6848 28690 6860
rect 30101 6851 30159 6857
rect 30101 6848 30113 6851
rect 28684 6820 30113 6848
rect 28684 6808 28690 6820
rect 30101 6817 30113 6820
rect 30147 6817 30159 6851
rect 30101 6811 30159 6817
rect 30926 6808 30932 6860
rect 30984 6848 30990 6860
rect 33778 6848 33784 6860
rect 30984 6820 33784 6848
rect 30984 6808 30990 6820
rect 33778 6808 33784 6820
rect 33836 6848 33842 6860
rect 35544 6857 35572 6888
rect 33965 6851 34023 6857
rect 33965 6848 33977 6851
rect 33836 6820 33977 6848
rect 33836 6808 33842 6820
rect 33965 6817 33977 6820
rect 34011 6817 34023 6851
rect 33965 6811 34023 6817
rect 35529 6851 35587 6857
rect 35529 6817 35541 6851
rect 35575 6848 35587 6851
rect 36814 6848 36820 6860
rect 35575 6820 36820 6848
rect 35575 6817 35587 6820
rect 35529 6811 35587 6817
rect 36814 6808 36820 6820
rect 36872 6848 36878 6860
rect 40034 6848 40040 6860
rect 36872 6820 40040 6848
rect 36872 6808 36878 6820
rect 40034 6808 40040 6820
rect 40092 6808 40098 6860
rect 46842 6808 46848 6860
rect 46900 6848 46906 6860
rect 47397 6851 47455 6857
rect 47397 6848 47409 6851
rect 46900 6820 47409 6848
rect 46900 6808 46906 6820
rect 47397 6817 47409 6820
rect 47443 6848 47455 6851
rect 49602 6848 49608 6860
rect 47443 6820 49608 6848
rect 47443 6817 47455 6820
rect 47397 6811 47455 6817
rect 49602 6808 49608 6820
rect 49660 6808 49666 6860
rect 56870 6808 56876 6860
rect 56928 6808 56934 6860
rect 26605 6783 26663 6789
rect 26605 6749 26617 6783
rect 26651 6749 26663 6783
rect 26605 6743 26663 6749
rect 26970 6740 26976 6792
rect 27028 6740 27034 6792
rect 27065 6783 27123 6789
rect 27065 6749 27077 6783
rect 27111 6749 27123 6783
rect 29733 6783 29791 6789
rect 29733 6780 29745 6783
rect 27065 6743 27123 6749
rect 27172 6752 29745 6780
rect 11330 6712 11336 6724
rect 11164 6684 11336 6712
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 13541 6715 13599 6721
rect 13541 6681 13553 6715
rect 13587 6712 13599 6715
rect 14369 6715 14427 6721
rect 13587 6684 13768 6712
rect 13587 6681 13599 6684
rect 13541 6675 13599 6681
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 9677 6647 9735 6653
rect 9677 6644 9689 6647
rect 9548 6616 9689 6644
rect 9548 6604 9554 6616
rect 9677 6613 9689 6616
rect 9723 6613 9735 6647
rect 9677 6607 9735 6613
rect 11698 6604 11704 6656
rect 11756 6644 11762 6656
rect 13556 6644 13584 6675
rect 11756 6616 13584 6644
rect 13740 6644 13768 6684
rect 14369 6681 14381 6715
rect 14415 6712 14427 6715
rect 16114 6712 16120 6724
rect 14415 6684 16120 6712
rect 14415 6681 14427 6684
rect 14369 6675 14427 6681
rect 16114 6672 16120 6684
rect 16172 6672 16178 6724
rect 16669 6715 16727 6721
rect 16669 6712 16681 6715
rect 16224 6684 16681 6712
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 13740 6616 14473 6644
rect 11756 6604 11762 6616
rect 14461 6613 14473 6616
rect 14507 6613 14519 6647
rect 14461 6607 14519 6613
rect 15746 6604 15752 6656
rect 15804 6644 15810 6656
rect 16224 6644 16252 6684
rect 16669 6681 16681 6684
rect 16715 6712 16727 6715
rect 17862 6712 17868 6724
rect 16715 6684 17868 6712
rect 16715 6681 16727 6684
rect 16669 6675 16727 6681
rect 17862 6672 17868 6684
rect 17920 6672 17926 6724
rect 17954 6672 17960 6724
rect 18012 6712 18018 6724
rect 18230 6712 18236 6724
rect 18012 6684 18236 6712
rect 18012 6672 18018 6684
rect 18230 6672 18236 6684
rect 18288 6672 18294 6724
rect 19426 6672 19432 6724
rect 19484 6712 19490 6724
rect 19981 6715 20039 6721
rect 19981 6712 19993 6715
rect 19484 6684 19993 6712
rect 19484 6672 19490 6684
rect 19981 6681 19993 6684
rect 20027 6712 20039 6715
rect 20438 6712 20444 6724
rect 20027 6684 20444 6712
rect 20027 6681 20039 6684
rect 19981 6675 20039 6681
rect 20438 6672 20444 6684
rect 20496 6672 20502 6724
rect 21085 6715 21143 6721
rect 21085 6681 21097 6715
rect 21131 6712 21143 6715
rect 22370 6712 22376 6724
rect 21131 6684 22376 6712
rect 21131 6681 21143 6684
rect 21085 6675 21143 6681
rect 22370 6672 22376 6684
rect 22428 6672 22434 6724
rect 22646 6672 22652 6724
rect 22704 6672 22710 6724
rect 22848 6684 25912 6712
rect 15804 6616 16252 6644
rect 15804 6604 15810 6616
rect 16574 6604 16580 6656
rect 16632 6644 16638 6656
rect 21177 6647 21235 6653
rect 21177 6644 21189 6647
rect 16632 6616 21189 6644
rect 16632 6604 16638 6616
rect 21177 6613 21189 6616
rect 21223 6644 21235 6647
rect 21450 6644 21456 6656
rect 21223 6616 21456 6644
rect 21223 6613 21235 6616
rect 21177 6607 21235 6613
rect 21450 6604 21456 6616
rect 21508 6604 21514 6656
rect 22186 6604 22192 6656
rect 22244 6644 22250 6656
rect 22848 6644 22876 6684
rect 22244 6616 22876 6644
rect 22244 6604 22250 6616
rect 23842 6604 23848 6656
rect 23900 6604 23906 6656
rect 24765 6647 24823 6653
rect 24765 6613 24777 6647
rect 24811 6644 24823 6647
rect 25038 6644 25044 6656
rect 24811 6616 25044 6644
rect 24811 6613 24823 6616
rect 24765 6607 24823 6613
rect 25038 6604 25044 6616
rect 25096 6604 25102 6656
rect 25130 6604 25136 6656
rect 25188 6604 25194 6656
rect 25225 6647 25283 6653
rect 25225 6613 25237 6647
rect 25271 6644 25283 6647
rect 25774 6644 25780 6656
rect 25271 6616 25780 6644
rect 25271 6613 25283 6616
rect 25225 6607 25283 6613
rect 25774 6604 25780 6616
rect 25832 6604 25838 6656
rect 25884 6644 25912 6684
rect 26786 6672 26792 6724
rect 26844 6712 26850 6724
rect 27080 6712 27108 6743
rect 26844 6684 27108 6712
rect 26844 6672 26850 6684
rect 27172 6644 27200 6752
rect 29733 6749 29745 6752
rect 29779 6749 29791 6783
rect 29733 6743 29791 6749
rect 30374 6740 30380 6792
rect 30432 6780 30438 6792
rect 31389 6783 31447 6789
rect 31389 6780 31401 6783
rect 30432 6752 31401 6780
rect 30432 6740 30438 6752
rect 31389 6749 31401 6752
rect 31435 6749 31447 6783
rect 33686 6780 33692 6792
rect 31389 6743 31447 6749
rect 31496 6752 33692 6780
rect 27798 6672 27804 6724
rect 27856 6712 27862 6724
rect 27985 6715 28043 6721
rect 27985 6712 27997 6715
rect 27856 6684 27997 6712
rect 27856 6672 27862 6684
rect 27985 6681 27997 6684
rect 28031 6681 28043 6715
rect 27985 6675 28043 6681
rect 28534 6672 28540 6724
rect 28592 6712 28598 6724
rect 30282 6712 30288 6724
rect 28592 6684 30288 6712
rect 28592 6672 28598 6684
rect 30282 6672 30288 6684
rect 30340 6672 30346 6724
rect 31202 6672 31208 6724
rect 31260 6672 31266 6724
rect 25884 6616 27200 6644
rect 28442 6604 28448 6656
rect 28500 6644 28506 6656
rect 28629 6647 28687 6653
rect 28629 6644 28641 6647
rect 28500 6616 28641 6644
rect 28500 6604 28506 6616
rect 28629 6613 28641 6616
rect 28675 6613 28687 6647
rect 28629 6607 28687 6613
rect 28718 6604 28724 6656
rect 28776 6644 28782 6656
rect 30834 6644 30840 6656
rect 28776 6616 30840 6644
rect 28776 6604 28782 6616
rect 30834 6604 30840 6616
rect 30892 6604 30898 6656
rect 31496 6653 31524 6752
rect 33686 6740 33692 6752
rect 33744 6740 33750 6792
rect 34149 6783 34207 6789
rect 34149 6749 34161 6783
rect 34195 6780 34207 6783
rect 45189 6783 45247 6789
rect 34195 6752 34928 6780
rect 34195 6749 34207 6752
rect 34149 6743 34207 6749
rect 31754 6672 31760 6724
rect 31812 6672 31818 6724
rect 32582 6672 32588 6724
rect 32640 6712 32646 6724
rect 34790 6712 34796 6724
rect 32640 6684 34796 6712
rect 32640 6672 32646 6684
rect 34790 6672 34796 6684
rect 34848 6672 34854 6724
rect 31481 6647 31539 6653
rect 31481 6613 31493 6647
rect 31527 6613 31539 6647
rect 31481 6607 31539 6613
rect 31573 6647 31631 6653
rect 31573 6613 31585 6647
rect 31619 6644 31631 6647
rect 31938 6644 31944 6656
rect 31619 6616 31944 6644
rect 31619 6613 31631 6616
rect 31573 6607 31631 6613
rect 31938 6604 31944 6616
rect 31996 6644 32002 6656
rect 33134 6644 33140 6656
rect 31996 6616 33140 6644
rect 31996 6604 32002 6616
rect 33134 6604 33140 6616
rect 33192 6604 33198 6656
rect 34900 6653 34928 6752
rect 45189 6749 45201 6783
rect 45235 6780 45247 6783
rect 46934 6780 46940 6792
rect 45235 6752 46940 6780
rect 45235 6749 45247 6752
rect 45189 6743 45247 6749
rect 46934 6740 46940 6752
rect 46992 6740 46998 6792
rect 56962 6740 56968 6792
rect 57020 6780 57026 6792
rect 57129 6783 57187 6789
rect 57129 6780 57141 6783
rect 57020 6752 57141 6780
rect 57020 6740 57026 6752
rect 57129 6749 57141 6752
rect 57175 6749 57187 6783
rect 57129 6743 57187 6749
rect 45456 6715 45514 6721
rect 45456 6681 45468 6715
rect 45502 6712 45514 6715
rect 45830 6712 45836 6724
rect 45502 6684 45836 6712
rect 45502 6681 45514 6684
rect 45456 6675 45514 6681
rect 45830 6672 45836 6684
rect 45888 6672 45894 6724
rect 47121 6715 47179 6721
rect 47121 6681 47133 6715
rect 47167 6681 47179 6715
rect 47121 6675 47179 6681
rect 34885 6647 34943 6653
rect 34885 6613 34897 6647
rect 34931 6613 34943 6647
rect 34885 6607 34943 6613
rect 35250 6604 35256 6656
rect 35308 6604 35314 6656
rect 35342 6604 35348 6656
rect 35400 6604 35406 6656
rect 43070 6604 43076 6656
rect 43128 6644 43134 6656
rect 47136 6644 47164 6675
rect 43128 6616 47164 6644
rect 43128 6604 43134 6616
rect 58250 6604 58256 6656
rect 58308 6604 58314 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 9122 6400 9128 6452
rect 9180 6400 9186 6452
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6440 13231 6443
rect 13354 6440 13360 6452
rect 13219 6412 13360 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 13354 6400 13360 6412
rect 13412 6440 13418 6452
rect 19242 6440 19248 6452
rect 13412 6412 13768 6440
rect 13412 6400 13418 6412
rect 13740 6381 13768 6412
rect 15120 6412 19248 6440
rect 13725 6375 13783 6381
rect 13725 6341 13737 6375
rect 13771 6341 13783 6375
rect 13725 6335 13783 6341
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 9122 6304 9128 6316
rect 1627 6276 9128 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6304 9459 6307
rect 9447 6276 12434 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 934 6196 940 6248
rect 992 6236 998 6248
rect 1765 6239 1823 6245
rect 1765 6236 1777 6239
rect 992 6208 1777 6236
rect 992 6196 998 6208
rect 1765 6205 1777 6208
rect 1811 6205 1823 6239
rect 1765 6199 1823 6205
rect 9306 6196 9312 6248
rect 9364 6196 9370 6248
rect 9490 6196 9496 6248
rect 9548 6196 9554 6248
rect 9585 6239 9643 6245
rect 9585 6205 9597 6239
rect 9631 6236 9643 6239
rect 10410 6236 10416 6248
rect 9631 6208 10416 6236
rect 9631 6205 9643 6208
rect 9585 6199 9643 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 12406 6236 12434 6276
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 12989 6307 13047 6313
rect 12989 6304 13001 6307
rect 12676 6276 13001 6304
rect 12676 6264 12682 6276
rect 12989 6273 13001 6276
rect 13035 6273 13047 6307
rect 12989 6267 13047 6273
rect 15120 6236 15148 6412
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 19978 6400 19984 6452
rect 20036 6440 20042 6452
rect 20990 6440 20996 6452
rect 20036 6412 20996 6440
rect 20036 6400 20042 6412
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 23017 6443 23075 6449
rect 23017 6409 23029 6443
rect 23063 6440 23075 6443
rect 23106 6440 23112 6452
rect 23063 6412 23112 6440
rect 23063 6409 23075 6412
rect 23017 6403 23075 6409
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 25130 6440 25136 6452
rect 23584 6412 25136 6440
rect 15194 6332 15200 6384
rect 15252 6372 15258 6384
rect 15289 6375 15347 6381
rect 15289 6372 15301 6375
rect 15252 6344 15301 6372
rect 15252 6332 15258 6344
rect 15289 6341 15301 6344
rect 15335 6341 15347 6375
rect 15289 6335 15347 6341
rect 16853 6375 16911 6381
rect 16853 6341 16865 6375
rect 16899 6372 16911 6375
rect 18046 6372 18052 6384
rect 16899 6344 18052 6372
rect 16899 6341 16911 6344
rect 16853 6335 16911 6341
rect 18046 6332 18052 6344
rect 18104 6372 18110 6384
rect 18509 6375 18567 6381
rect 18509 6372 18521 6375
rect 18104 6344 18521 6372
rect 18104 6332 18110 6344
rect 18509 6341 18521 6344
rect 18555 6341 18567 6375
rect 20254 6372 20260 6384
rect 18509 6335 18567 6341
rect 19444 6344 20260 6372
rect 15378 6264 15384 6316
rect 15436 6264 15442 6316
rect 15746 6264 15752 6316
rect 15804 6264 15810 6316
rect 15838 6264 15844 6316
rect 15896 6264 15902 6316
rect 15930 6264 15936 6316
rect 15988 6304 15994 6316
rect 16301 6307 16359 6313
rect 16301 6304 16313 6307
rect 15988 6276 16313 6304
rect 15988 6264 15994 6276
rect 16301 6273 16313 6276
rect 16347 6273 16359 6307
rect 16301 6267 16359 6273
rect 17494 6264 17500 6316
rect 17552 6304 17558 6316
rect 19444 6313 19472 6344
rect 20254 6332 20260 6344
rect 20312 6332 20318 6384
rect 23198 6332 23204 6384
rect 23256 6372 23262 6384
rect 23477 6375 23535 6381
rect 23477 6372 23489 6375
rect 23256 6344 23489 6372
rect 23256 6332 23262 6344
rect 23477 6341 23489 6344
rect 23523 6341 23535 6375
rect 23477 6335 23535 6341
rect 17589 6307 17647 6313
rect 17589 6304 17601 6307
rect 17552 6276 17601 6304
rect 17552 6264 17558 6276
rect 17589 6273 17601 6276
rect 17635 6273 17647 6307
rect 17589 6267 17647 6273
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6304 18291 6307
rect 19429 6307 19487 6313
rect 18279 6276 19380 6304
rect 18279 6273 18291 6276
rect 18233 6267 18291 6273
rect 12406 6208 15148 6236
rect 14001 6171 14059 6177
rect 14001 6168 14013 6171
rect 13096 6140 14013 6168
rect 7926 6060 7932 6112
rect 7984 6100 7990 6112
rect 13096 6100 13124 6140
rect 14001 6137 14013 6140
rect 14047 6137 14059 6171
rect 14001 6131 14059 6137
rect 14185 6171 14243 6177
rect 14185 6137 14197 6171
rect 14231 6168 14243 6171
rect 17954 6168 17960 6180
rect 14231 6140 17960 6168
rect 14231 6137 14243 6140
rect 14185 6131 14243 6137
rect 17954 6128 17960 6140
rect 18012 6128 18018 6180
rect 7984 6072 13124 6100
rect 19352 6100 19380 6276
rect 19429 6273 19441 6307
rect 19475 6273 19487 6307
rect 19429 6267 19487 6273
rect 19696 6307 19754 6313
rect 19696 6273 19708 6307
rect 19742 6304 19754 6307
rect 19978 6304 19984 6316
rect 19742 6276 19984 6304
rect 19742 6273 19754 6276
rect 19696 6267 19754 6273
rect 19978 6264 19984 6276
rect 20036 6264 20042 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 20824 6276 22017 6304
rect 20824 6177 20852 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 23382 6264 23388 6316
rect 23440 6264 23446 6316
rect 23584 6236 23612 6412
rect 25130 6400 25136 6412
rect 25188 6400 25194 6452
rect 28077 6443 28135 6449
rect 28077 6409 28089 6443
rect 28123 6440 28135 6443
rect 33042 6440 33048 6452
rect 28123 6412 33048 6440
rect 28123 6409 28135 6412
rect 28077 6403 28135 6409
rect 33042 6400 33048 6412
rect 33100 6400 33106 6452
rect 33134 6400 33140 6452
rect 33192 6440 33198 6452
rect 35250 6440 35256 6452
rect 33192 6412 35256 6440
rect 33192 6400 33198 6412
rect 35250 6400 35256 6412
rect 35308 6440 35314 6452
rect 35621 6443 35679 6449
rect 35621 6440 35633 6443
rect 35308 6412 35633 6440
rect 35308 6400 35314 6412
rect 35621 6409 35633 6412
rect 35667 6409 35679 6443
rect 35621 6403 35679 6409
rect 36446 6400 36452 6452
rect 36504 6440 36510 6452
rect 36541 6443 36599 6449
rect 36541 6440 36553 6443
rect 36504 6412 36553 6440
rect 36504 6400 36510 6412
rect 36541 6409 36553 6412
rect 36587 6409 36599 6443
rect 36541 6403 36599 6409
rect 38749 6443 38807 6449
rect 38749 6409 38761 6443
rect 38795 6440 38807 6443
rect 38838 6440 38844 6452
rect 38795 6412 38844 6440
rect 38795 6409 38807 6412
rect 38749 6403 38807 6409
rect 38838 6400 38844 6412
rect 38896 6400 38902 6452
rect 24578 6332 24584 6384
rect 24636 6372 24642 6384
rect 25038 6381 25044 6384
rect 25032 6372 25044 6381
rect 24636 6344 24900 6372
rect 24999 6344 25044 6372
rect 24636 6332 24642 6344
rect 24394 6264 24400 6316
rect 24452 6304 24458 6316
rect 24765 6307 24823 6313
rect 24765 6304 24777 6307
rect 24452 6276 24777 6304
rect 24452 6264 24458 6276
rect 24765 6273 24777 6276
rect 24811 6273 24823 6307
rect 24872 6304 24900 6344
rect 25032 6335 25044 6344
rect 25038 6332 25044 6335
rect 25096 6332 25102 6384
rect 25222 6332 25228 6384
rect 25280 6372 25286 6384
rect 25280 6344 28304 6372
rect 25280 6332 25286 6344
rect 24872 6276 26188 6304
rect 24765 6267 24823 6273
rect 20916 6208 23612 6236
rect 23661 6239 23719 6245
rect 20809 6171 20867 6177
rect 20809 6137 20821 6171
rect 20855 6137 20867 6171
rect 20809 6131 20867 6137
rect 20916 6100 20944 6208
rect 23661 6205 23673 6239
rect 23707 6236 23719 6239
rect 24026 6236 24032 6248
rect 23707 6208 24032 6236
rect 23707 6205 23719 6208
rect 23661 6199 23719 6205
rect 24026 6196 24032 6208
rect 24084 6236 24090 6248
rect 24302 6236 24308 6248
rect 24084 6208 24308 6236
rect 24084 6196 24090 6208
rect 24302 6196 24308 6208
rect 24360 6196 24366 6248
rect 21082 6128 21088 6180
rect 21140 6168 21146 6180
rect 26160 6168 26188 6276
rect 27338 6264 27344 6316
rect 27396 6304 27402 6316
rect 27525 6307 27583 6313
rect 27525 6304 27537 6307
rect 27396 6276 27537 6304
rect 27396 6264 27402 6276
rect 27525 6273 27537 6276
rect 27571 6273 27583 6307
rect 27525 6267 27583 6273
rect 27614 6264 27620 6316
rect 27672 6304 27678 6316
rect 28276 6304 28304 6344
rect 28534 6332 28540 6384
rect 28592 6372 28598 6384
rect 28997 6375 29055 6381
rect 28997 6372 29009 6375
rect 28592 6344 29009 6372
rect 28592 6332 28598 6344
rect 28997 6341 29009 6344
rect 29043 6341 29055 6375
rect 28997 6335 29055 6341
rect 29362 6332 29368 6384
rect 29420 6372 29426 6384
rect 29420 6344 30052 6372
rect 29420 6332 29426 6344
rect 28626 6304 28632 6316
rect 27672 6276 28212 6304
rect 28276 6276 28632 6304
rect 27672 6264 27678 6276
rect 26602 6196 26608 6248
rect 26660 6236 26666 6248
rect 27798 6236 27804 6248
rect 26660 6208 27804 6236
rect 26660 6196 26666 6208
rect 27798 6196 27804 6208
rect 27856 6196 27862 6248
rect 28184 6236 28212 6276
rect 28626 6264 28632 6276
rect 28684 6264 28690 6316
rect 29270 6264 29276 6316
rect 29328 6304 29334 6316
rect 30024 6313 30052 6344
rect 33778 6332 33784 6384
rect 33836 6372 33842 6384
rect 34793 6375 34851 6381
rect 34793 6372 34805 6375
rect 33836 6344 34805 6372
rect 33836 6332 33842 6344
rect 34793 6341 34805 6344
rect 34839 6341 34851 6375
rect 34793 6335 34851 6341
rect 35526 6332 35532 6384
rect 35584 6332 35590 6384
rect 36906 6332 36912 6384
rect 36964 6372 36970 6384
rect 43254 6372 43260 6384
rect 36964 6344 43260 6372
rect 36964 6332 36970 6344
rect 43254 6332 43260 6344
rect 43312 6332 43318 6384
rect 46842 6372 46848 6384
rect 46308 6344 46848 6372
rect 29733 6307 29791 6313
rect 29733 6304 29745 6307
rect 29328 6276 29745 6304
rect 29328 6264 29334 6276
rect 29733 6273 29745 6276
rect 29779 6273 29791 6307
rect 29733 6267 29791 6273
rect 30009 6307 30067 6313
rect 30009 6273 30021 6307
rect 30055 6273 30067 6307
rect 30926 6304 30932 6316
rect 30009 6267 30067 6273
rect 30116 6276 30932 6304
rect 30116 6236 30144 6276
rect 30926 6264 30932 6276
rect 30984 6264 30990 6316
rect 31110 6264 31116 6316
rect 31168 6264 31174 6316
rect 34514 6264 34520 6316
rect 34572 6264 34578 6316
rect 36078 6264 36084 6316
rect 36136 6304 36142 6316
rect 36449 6307 36507 6313
rect 36449 6304 36461 6307
rect 36136 6276 36461 6304
rect 36136 6264 36142 6276
rect 36449 6273 36461 6276
rect 36495 6273 36507 6307
rect 36449 6267 36507 6273
rect 38470 6264 38476 6316
rect 38528 6304 38534 6316
rect 46308 6313 46336 6344
rect 46842 6332 46848 6344
rect 46900 6332 46906 6384
rect 38565 6307 38623 6313
rect 38565 6304 38577 6307
rect 38528 6276 38577 6304
rect 38528 6264 38534 6276
rect 38565 6273 38577 6276
rect 38611 6273 38623 6307
rect 38565 6267 38623 6273
rect 46293 6307 46351 6313
rect 46293 6273 46305 6307
rect 46339 6273 46351 6307
rect 46293 6267 46351 6273
rect 46382 6264 46388 6316
rect 46440 6264 46446 6316
rect 58066 6264 58072 6316
rect 58124 6264 58130 6316
rect 28184 6208 30144 6236
rect 30193 6239 30251 6245
rect 30193 6205 30205 6239
rect 30239 6205 30251 6239
rect 30193 6199 30251 6205
rect 21140 6140 24808 6168
rect 26160 6140 28304 6168
rect 21140 6128 21146 6140
rect 19352 6072 20944 6100
rect 7984 6060 7990 6072
rect 20990 6060 20996 6112
rect 21048 6100 21054 6112
rect 22189 6103 22247 6109
rect 22189 6100 22201 6103
rect 21048 6072 22201 6100
rect 21048 6060 21054 6072
rect 22189 6069 22201 6072
rect 22235 6100 22247 6103
rect 24670 6100 24676 6112
rect 22235 6072 24676 6100
rect 22235 6069 22247 6072
rect 22189 6063 22247 6069
rect 24670 6060 24676 6072
rect 24728 6060 24734 6112
rect 24780 6100 24808 6140
rect 26050 6100 26056 6112
rect 24780 6072 26056 6100
rect 26050 6060 26056 6072
rect 26108 6060 26114 6112
rect 26142 6060 26148 6112
rect 26200 6060 26206 6112
rect 27893 6103 27951 6109
rect 27893 6069 27905 6103
rect 27939 6100 27951 6103
rect 27982 6100 27988 6112
rect 27939 6072 27988 6100
rect 27939 6069 27951 6072
rect 27893 6063 27951 6069
rect 27982 6060 27988 6072
rect 28040 6060 28046 6112
rect 28276 6100 28304 6140
rect 28350 6128 28356 6180
rect 28408 6168 28414 6180
rect 28902 6168 28908 6180
rect 28408 6140 28908 6168
rect 28408 6128 28414 6140
rect 28902 6128 28908 6140
rect 28960 6168 28966 6180
rect 29825 6171 29883 6177
rect 29825 6168 29837 6171
rect 28960 6140 29837 6168
rect 28960 6128 28966 6140
rect 29825 6137 29837 6140
rect 29871 6137 29883 6171
rect 29825 6131 29883 6137
rect 29914 6128 29920 6180
rect 29972 6168 29978 6180
rect 30208 6168 30236 6199
rect 36722 6196 36728 6248
rect 36780 6236 36786 6248
rect 43438 6236 43444 6248
rect 36780 6208 43444 6236
rect 36780 6196 36786 6208
rect 43438 6196 43444 6208
rect 43496 6196 43502 6248
rect 46566 6196 46572 6248
rect 46624 6196 46630 6248
rect 29972 6140 30236 6168
rect 29972 6128 29978 6140
rect 30374 6128 30380 6180
rect 30432 6168 30438 6180
rect 38194 6168 38200 6180
rect 30432 6140 38200 6168
rect 30432 6128 30438 6140
rect 38194 6128 38200 6140
rect 38252 6128 38258 6180
rect 56410 6168 56416 6180
rect 43364 6140 56416 6168
rect 30742 6100 30748 6112
rect 28276 6072 30748 6100
rect 30742 6060 30748 6072
rect 30800 6060 30806 6112
rect 31297 6103 31355 6109
rect 31297 6069 31309 6103
rect 31343 6100 31355 6103
rect 31386 6100 31392 6112
rect 31343 6072 31392 6100
rect 31343 6069 31355 6072
rect 31297 6063 31355 6069
rect 31386 6060 31392 6072
rect 31444 6060 31450 6112
rect 32950 6060 32956 6112
rect 33008 6100 33014 6112
rect 43364 6100 43392 6140
rect 56410 6128 56416 6140
rect 56468 6128 56474 6180
rect 33008 6072 43392 6100
rect 33008 6060 33014 6072
rect 43438 6060 43444 6112
rect 43496 6100 43502 6112
rect 58253 6103 58311 6109
rect 58253 6100 58265 6103
rect 43496 6072 58265 6100
rect 43496 6060 43502 6072
rect 58253 6069 58265 6072
rect 58299 6069 58311 6103
rect 58253 6063 58311 6069
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 9122 5856 9128 5908
rect 9180 5856 9186 5908
rect 10873 5899 10931 5905
rect 10873 5865 10885 5899
rect 10919 5896 10931 5899
rect 11054 5896 11060 5908
rect 10919 5868 11060 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 16684 5868 23520 5896
rect 7834 5788 7840 5840
rect 7892 5828 7898 5840
rect 10689 5831 10747 5837
rect 10689 5828 10701 5831
rect 7892 5800 10701 5828
rect 7892 5788 7898 5800
rect 10689 5797 10701 5800
rect 10735 5797 10747 5831
rect 10689 5791 10747 5797
rect 9401 5763 9459 5769
rect 9401 5729 9413 5763
rect 9447 5760 9459 5763
rect 16574 5760 16580 5772
rect 9447 5732 16580 5760
rect 9447 5729 9459 5732
rect 9401 5723 9459 5729
rect 16574 5720 16580 5732
rect 16632 5720 16638 5772
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5692 1639 5695
rect 1627 5664 2774 5692
rect 1627 5661 1639 5664
rect 1581 5655 1639 5661
rect 934 5584 940 5636
rect 992 5624 998 5636
rect 1857 5627 1915 5633
rect 1857 5624 1869 5627
rect 992 5596 1869 5624
rect 992 5584 998 5596
rect 1857 5593 1869 5596
rect 1903 5593 1915 5627
rect 1857 5587 1915 5593
rect 2746 5556 2774 5664
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 9490 5652 9496 5704
rect 9548 5652 9554 5704
rect 9582 5652 9588 5704
rect 9640 5652 9646 5704
rect 16684 5692 16712 5868
rect 17678 5788 17684 5840
rect 17736 5828 17742 5840
rect 17957 5831 18015 5837
rect 17957 5828 17969 5831
rect 17736 5800 17969 5828
rect 17736 5788 17742 5800
rect 17957 5797 17969 5800
rect 18003 5797 18015 5831
rect 17957 5791 18015 5797
rect 22005 5831 22063 5837
rect 22005 5797 22017 5831
rect 22051 5797 22063 5831
rect 23492 5828 23520 5868
rect 23566 5856 23572 5908
rect 23624 5856 23630 5908
rect 23934 5856 23940 5908
rect 23992 5896 23998 5908
rect 25133 5899 25191 5905
rect 25133 5896 25145 5899
rect 23992 5868 25145 5896
rect 23992 5856 23998 5868
rect 25133 5865 25145 5868
rect 25179 5865 25191 5899
rect 25133 5859 25191 5865
rect 25774 5856 25780 5908
rect 25832 5856 25838 5908
rect 26050 5856 26056 5908
rect 26108 5896 26114 5908
rect 30374 5896 30380 5908
rect 26108 5868 30380 5896
rect 26108 5856 26114 5868
rect 30374 5856 30380 5868
rect 30432 5856 30438 5908
rect 31018 5896 31024 5908
rect 30668 5868 31024 5896
rect 24486 5828 24492 5840
rect 23492 5800 24492 5828
rect 22005 5791 22063 5797
rect 19797 5763 19855 5769
rect 19797 5729 19809 5763
rect 19843 5760 19855 5763
rect 19843 5732 19932 5760
rect 19843 5729 19855 5732
rect 19797 5723 19855 5729
rect 9692 5664 16712 5692
rect 17037 5695 17095 5701
rect 9324 5624 9352 5652
rect 9692 5624 9720 5664
rect 17037 5661 17049 5695
rect 17083 5692 17095 5695
rect 17310 5692 17316 5704
rect 17083 5664 17316 5692
rect 17083 5661 17095 5664
rect 17037 5655 17095 5661
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5661 17463 5695
rect 17405 5655 17463 5661
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5692 17831 5695
rect 18046 5692 18052 5704
rect 17819 5664 18052 5692
rect 17819 5661 17831 5664
rect 17773 5655 17831 5661
rect 9324 5596 9720 5624
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 10413 5627 10471 5633
rect 10413 5624 10425 5627
rect 10100 5596 10425 5624
rect 10100 5584 10106 5596
rect 10413 5593 10425 5596
rect 10459 5624 10471 5627
rect 10594 5624 10600 5636
rect 10459 5596 10600 5624
rect 10459 5593 10471 5596
rect 10413 5587 10471 5593
rect 10594 5584 10600 5596
rect 10652 5584 10658 5636
rect 12710 5584 12716 5636
rect 12768 5624 12774 5636
rect 17420 5624 17448 5655
rect 18046 5652 18052 5664
rect 18104 5652 18110 5704
rect 18414 5652 18420 5704
rect 18472 5652 18478 5704
rect 17862 5624 17868 5636
rect 12768 5596 17356 5624
rect 17420 5596 17868 5624
rect 12768 5584 12774 5596
rect 10226 5556 10232 5568
rect 2746 5528 10232 5556
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 14458 5556 14464 5568
rect 10376 5528 14464 5556
rect 10376 5516 10382 5528
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 17328 5556 17356 5596
rect 17862 5584 17868 5596
rect 17920 5624 17926 5636
rect 19426 5624 19432 5636
rect 17920 5596 19432 5624
rect 17920 5584 17926 5596
rect 19426 5584 19432 5596
rect 19484 5584 19490 5636
rect 19904 5624 19932 5732
rect 20064 5695 20122 5701
rect 20064 5661 20076 5695
rect 20110 5692 20122 5695
rect 22020 5692 22048 5791
rect 24486 5788 24492 5800
rect 24544 5788 24550 5840
rect 27706 5828 27712 5840
rect 25332 5800 27712 5828
rect 22465 5763 22523 5769
rect 22465 5760 22477 5763
rect 20110 5664 22048 5692
rect 22112 5732 22477 5760
rect 20110 5661 20122 5664
rect 20064 5655 20122 5661
rect 20254 5624 20260 5636
rect 19904 5596 20260 5624
rect 20254 5584 20260 5596
rect 20312 5584 20318 5636
rect 21082 5624 21088 5636
rect 20916 5596 21088 5624
rect 20916 5556 20944 5596
rect 21082 5584 21088 5596
rect 21140 5584 21146 5636
rect 22112 5624 22140 5732
rect 22465 5729 22477 5732
rect 22511 5729 22523 5763
rect 22465 5723 22523 5729
rect 22649 5763 22707 5769
rect 22649 5729 22661 5763
rect 22695 5760 22707 5763
rect 23934 5760 23940 5772
rect 22695 5732 23940 5760
rect 22695 5729 22707 5732
rect 22649 5723 22707 5729
rect 22664 5692 22692 5723
rect 23934 5720 23940 5732
rect 23992 5720 23998 5772
rect 25332 5760 25360 5800
rect 27706 5788 27712 5800
rect 27764 5788 27770 5840
rect 28902 5788 28908 5840
rect 28960 5828 28966 5840
rect 29089 5831 29147 5837
rect 29089 5828 29101 5831
rect 28960 5800 29101 5828
rect 28960 5788 28966 5800
rect 29089 5797 29101 5800
rect 29135 5797 29147 5831
rect 29089 5791 29147 5797
rect 29825 5831 29883 5837
rect 29825 5797 29837 5831
rect 29871 5797 29883 5831
rect 29825 5791 29883 5797
rect 24044 5732 25360 5760
rect 21192 5596 22140 5624
rect 22204 5664 22692 5692
rect 23293 5695 23351 5701
rect 17328 5528 20944 5556
rect 20990 5516 20996 5568
rect 21048 5556 21054 5568
rect 21192 5565 21220 5596
rect 21177 5559 21235 5565
rect 21177 5556 21189 5559
rect 21048 5528 21189 5556
rect 21048 5516 21054 5528
rect 21177 5525 21189 5528
rect 21223 5525 21235 5559
rect 21177 5519 21235 5525
rect 21266 5516 21272 5568
rect 21324 5556 21330 5568
rect 22204 5556 22232 5664
rect 23293 5661 23305 5695
rect 23339 5692 23351 5695
rect 23842 5692 23848 5704
rect 23339 5664 23848 5692
rect 23339 5661 23351 5664
rect 23293 5655 23351 5661
rect 23842 5652 23848 5664
rect 23900 5652 23906 5704
rect 21324 5528 22232 5556
rect 22373 5559 22431 5565
rect 21324 5516 21330 5528
rect 22373 5525 22385 5559
rect 22419 5556 22431 5559
rect 24044 5556 24072 5732
rect 26050 5720 26056 5772
rect 26108 5760 26114 5772
rect 26329 5763 26387 5769
rect 26329 5760 26341 5763
rect 26108 5732 26341 5760
rect 26108 5720 26114 5732
rect 26329 5729 26341 5732
rect 26375 5729 26387 5763
rect 26329 5723 26387 5729
rect 26418 5720 26424 5772
rect 26476 5760 26482 5772
rect 29840 5760 29868 5791
rect 26476 5732 29868 5760
rect 26476 5720 26482 5732
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5692 25007 5695
rect 25314 5692 25320 5704
rect 24995 5664 25320 5692
rect 24995 5661 25007 5664
rect 24949 5655 25007 5661
rect 25314 5652 25320 5664
rect 25372 5652 25378 5704
rect 26970 5652 26976 5704
rect 27028 5692 27034 5704
rect 28537 5695 28595 5701
rect 28537 5692 28549 5695
rect 27028 5664 28549 5692
rect 27028 5652 27034 5664
rect 28537 5661 28549 5664
rect 28583 5661 28595 5695
rect 28537 5655 28595 5661
rect 28626 5652 28632 5704
rect 28684 5692 28690 5704
rect 28910 5695 28968 5701
rect 28910 5692 28922 5695
rect 28684 5664 28922 5692
rect 28684 5652 28690 5664
rect 28910 5661 28922 5664
rect 28956 5661 28968 5695
rect 28910 5655 28968 5661
rect 29638 5652 29644 5704
rect 29696 5652 29702 5704
rect 30285 5695 30343 5701
rect 30285 5661 30297 5695
rect 30331 5692 30343 5695
rect 30374 5692 30380 5704
rect 30331 5664 30380 5692
rect 30331 5661 30343 5664
rect 30285 5655 30343 5661
rect 30374 5652 30380 5664
rect 30432 5692 30438 5704
rect 30561 5695 30619 5701
rect 30561 5692 30573 5695
rect 30432 5664 30573 5692
rect 30432 5652 30438 5664
rect 30561 5661 30573 5664
rect 30607 5661 30619 5695
rect 30561 5655 30619 5661
rect 24118 5584 24124 5636
rect 24176 5624 24182 5636
rect 26145 5627 26203 5633
rect 26145 5624 26157 5627
rect 24176 5596 26157 5624
rect 24176 5584 24182 5596
rect 26145 5593 26157 5596
rect 26191 5593 26203 5627
rect 26145 5587 26203 5593
rect 26786 5584 26792 5636
rect 26844 5624 26850 5636
rect 28721 5627 28779 5633
rect 28721 5624 28733 5627
rect 26844 5596 28733 5624
rect 26844 5584 26850 5596
rect 28721 5593 28733 5596
rect 28767 5593 28779 5627
rect 28721 5587 28779 5593
rect 28810 5584 28816 5636
rect 28868 5584 28874 5636
rect 22419 5528 24072 5556
rect 22419 5525 22431 5528
rect 22373 5519 22431 5525
rect 24302 5516 24308 5568
rect 24360 5556 24366 5568
rect 26050 5556 26056 5568
rect 24360 5528 26056 5556
rect 24360 5516 24366 5528
rect 26050 5516 26056 5528
rect 26108 5516 26114 5568
rect 26237 5559 26295 5565
rect 26237 5525 26249 5559
rect 26283 5556 26295 5559
rect 30668 5556 30696 5868
rect 31018 5856 31024 5868
rect 31076 5896 31082 5908
rect 32677 5899 32735 5905
rect 32677 5896 32689 5899
rect 31076 5868 32689 5896
rect 31076 5856 31082 5868
rect 32677 5865 32689 5868
rect 32723 5896 32735 5899
rect 32766 5896 32772 5908
rect 32723 5868 32772 5896
rect 32723 5865 32735 5868
rect 32677 5859 32735 5865
rect 32766 5856 32772 5868
rect 32824 5856 32830 5908
rect 33042 5856 33048 5908
rect 33100 5896 33106 5908
rect 35526 5896 35532 5908
rect 33100 5868 35532 5896
rect 33100 5856 33106 5868
rect 35526 5856 35532 5868
rect 35584 5856 35590 5908
rect 35618 5856 35624 5908
rect 35676 5896 35682 5908
rect 37369 5899 37427 5905
rect 37369 5896 37381 5899
rect 35676 5868 37381 5896
rect 35676 5856 35682 5868
rect 37369 5865 37381 5868
rect 37415 5865 37427 5899
rect 37369 5859 37427 5865
rect 37642 5856 37648 5908
rect 37700 5896 37706 5908
rect 38013 5899 38071 5905
rect 38013 5896 38025 5899
rect 37700 5868 38025 5896
rect 37700 5856 37706 5868
rect 38013 5865 38025 5868
rect 38059 5865 38071 5899
rect 38013 5859 38071 5865
rect 30742 5788 30748 5840
rect 30800 5788 30806 5840
rect 41601 5831 41659 5837
rect 41601 5828 41613 5831
rect 38304 5800 41613 5828
rect 31294 5720 31300 5772
rect 31352 5720 31358 5772
rect 33597 5763 33655 5769
rect 33597 5729 33609 5763
rect 33643 5760 33655 5763
rect 35894 5760 35900 5772
rect 33643 5732 35900 5760
rect 33643 5729 33655 5732
rect 33597 5723 33655 5729
rect 35894 5720 35900 5732
rect 35952 5720 35958 5772
rect 35986 5720 35992 5772
rect 36044 5760 36050 5772
rect 36262 5760 36268 5772
rect 36044 5732 36268 5760
rect 36044 5720 36050 5732
rect 36262 5720 36268 5732
rect 36320 5760 36326 5772
rect 36449 5763 36507 5769
rect 36449 5760 36461 5763
rect 36320 5732 36461 5760
rect 36320 5720 36326 5732
rect 36449 5729 36461 5732
rect 36495 5729 36507 5763
rect 36449 5723 36507 5729
rect 36633 5763 36691 5769
rect 36633 5729 36645 5763
rect 36679 5760 36691 5763
rect 36814 5760 36820 5772
rect 36679 5732 36820 5760
rect 36679 5729 36691 5732
rect 36633 5723 36691 5729
rect 36814 5720 36820 5732
rect 36872 5720 36878 5772
rect 37090 5720 37096 5772
rect 37148 5760 37154 5772
rect 38304 5760 38332 5800
rect 41601 5797 41613 5800
rect 41647 5797 41659 5831
rect 58250 5828 58256 5840
rect 41601 5791 41659 5797
rect 56980 5800 58256 5828
rect 37148 5732 38332 5760
rect 37148 5720 37154 5732
rect 38378 5720 38384 5772
rect 38436 5760 38442 5772
rect 39209 5763 39267 5769
rect 39209 5760 39221 5763
rect 38436 5732 39221 5760
rect 38436 5720 38442 5732
rect 39209 5729 39221 5732
rect 39255 5729 39267 5763
rect 39209 5723 39267 5729
rect 39393 5763 39451 5769
rect 39393 5729 39405 5763
rect 39439 5760 39451 5763
rect 40034 5760 40040 5772
rect 39439 5732 40040 5760
rect 39439 5729 39451 5732
rect 39393 5723 39451 5729
rect 31386 5652 31392 5704
rect 31444 5692 31450 5704
rect 31553 5695 31611 5701
rect 31553 5692 31565 5695
rect 31444 5664 31565 5692
rect 31444 5652 31450 5664
rect 31553 5661 31565 5664
rect 31599 5661 31611 5695
rect 31553 5655 31611 5661
rect 34054 5652 34060 5704
rect 34112 5692 34118 5704
rect 34149 5695 34207 5701
rect 34149 5692 34161 5695
rect 34112 5664 34161 5692
rect 34112 5652 34118 5664
rect 34149 5661 34161 5664
rect 34195 5661 34207 5695
rect 34149 5655 34207 5661
rect 34333 5695 34391 5701
rect 34333 5661 34345 5695
rect 34379 5692 34391 5695
rect 35434 5692 35440 5704
rect 34379 5664 35440 5692
rect 34379 5661 34391 5664
rect 34333 5655 34391 5661
rect 35434 5652 35440 5664
rect 35492 5652 35498 5704
rect 39224 5692 39252 5723
rect 40034 5720 40040 5732
rect 40092 5720 40098 5772
rect 56980 5701 57008 5800
rect 58250 5788 58256 5800
rect 58308 5788 58314 5840
rect 57241 5763 57299 5769
rect 57241 5729 57253 5763
rect 57287 5760 57299 5763
rect 58986 5760 58992 5772
rect 57287 5732 58992 5760
rect 57287 5729 57299 5732
rect 57241 5723 57299 5729
rect 58986 5720 58992 5732
rect 59044 5720 59050 5772
rect 56965 5695 57023 5701
rect 39224 5664 51074 5692
rect 33413 5627 33471 5633
rect 33413 5593 33425 5627
rect 33459 5624 33471 5627
rect 34977 5627 35035 5633
rect 33459 5596 34284 5624
rect 33459 5593 33471 5596
rect 33413 5587 33471 5593
rect 34256 5568 34284 5596
rect 34977 5593 34989 5627
rect 35023 5593 35035 5627
rect 34977 5587 35035 5593
rect 26283 5528 30696 5556
rect 26283 5525 26295 5528
rect 26237 5519 26295 5525
rect 34238 5516 34244 5568
rect 34296 5556 34302 5568
rect 34992 5556 35020 5587
rect 35158 5584 35164 5636
rect 35216 5584 35222 5636
rect 36262 5624 36268 5636
rect 35636 5596 36268 5624
rect 35636 5556 35664 5596
rect 36262 5584 36268 5596
rect 36320 5584 36326 5636
rect 36722 5584 36728 5636
rect 36780 5624 36786 5636
rect 37277 5627 37335 5633
rect 37277 5624 37289 5627
rect 36780 5596 37289 5624
rect 36780 5584 36786 5596
rect 37277 5593 37289 5596
rect 37323 5593 37335 5627
rect 37277 5587 37335 5593
rect 37921 5627 37979 5633
rect 37921 5593 37933 5627
rect 37967 5593 37979 5627
rect 37921 5587 37979 5593
rect 34296 5528 35664 5556
rect 35713 5559 35771 5565
rect 34296 5516 34302 5528
rect 35713 5525 35725 5559
rect 35759 5556 35771 5559
rect 35802 5556 35808 5568
rect 35759 5528 35808 5556
rect 35759 5525 35771 5528
rect 35713 5519 35771 5525
rect 35802 5516 35808 5528
rect 35860 5516 35866 5568
rect 35986 5516 35992 5568
rect 36044 5516 36050 5568
rect 36354 5516 36360 5568
rect 36412 5516 36418 5568
rect 36814 5516 36820 5568
rect 36872 5556 36878 5568
rect 37936 5556 37964 5587
rect 38838 5584 38844 5636
rect 38896 5624 38902 5636
rect 39117 5627 39175 5633
rect 39117 5624 39129 5627
rect 38896 5596 39129 5624
rect 38896 5584 38902 5596
rect 39117 5593 39129 5596
rect 39163 5593 39175 5627
rect 39117 5587 39175 5593
rect 41414 5584 41420 5636
rect 41472 5584 41478 5636
rect 36872 5528 37964 5556
rect 38749 5559 38807 5565
rect 36872 5516 36878 5528
rect 38749 5525 38761 5559
rect 38795 5556 38807 5559
rect 38930 5556 38936 5568
rect 38795 5528 38936 5556
rect 38795 5525 38807 5528
rect 38749 5519 38807 5525
rect 38930 5516 38936 5528
rect 38988 5516 38994 5568
rect 51046 5556 51074 5664
rect 56965 5661 56977 5695
rect 57011 5661 57023 5695
rect 56965 5655 57023 5661
rect 57882 5652 57888 5704
rect 57940 5652 57946 5704
rect 58161 5695 58219 5701
rect 58161 5661 58173 5695
rect 58207 5692 58219 5695
rect 58894 5692 58900 5704
rect 58207 5664 58900 5692
rect 58207 5661 58219 5664
rect 58161 5655 58219 5661
rect 58894 5652 58900 5664
rect 58952 5652 58958 5704
rect 57146 5556 57152 5568
rect 51046 5528 57152 5556
rect 57146 5516 57152 5528
rect 57204 5516 57210 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 9401 5355 9459 5361
rect 9401 5321 9413 5355
rect 9447 5352 9459 5355
rect 9582 5352 9588 5364
rect 9447 5324 9588 5352
rect 9447 5321 9459 5324
rect 9401 5315 9459 5321
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 10226 5312 10232 5364
rect 10284 5312 10290 5364
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 13817 5355 13875 5361
rect 12032 5324 13768 5352
rect 12032 5312 12038 5324
rect 13740 5284 13768 5324
rect 13817 5321 13829 5355
rect 13863 5352 13875 5355
rect 13906 5352 13912 5364
rect 13863 5324 13912 5352
rect 13863 5321 13875 5324
rect 13817 5315 13875 5321
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 15562 5312 15568 5364
rect 15620 5352 15626 5364
rect 16022 5352 16028 5364
rect 15620 5324 16028 5352
rect 15620 5312 15626 5324
rect 16022 5312 16028 5324
rect 16080 5352 16086 5364
rect 19613 5355 19671 5361
rect 16080 5324 19472 5352
rect 16080 5312 16086 5324
rect 13740 5256 19380 5284
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5216 1639 5219
rect 8110 5216 8116 5228
rect 1627 5188 8116 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5216 8263 5219
rect 8251 5188 8984 5216
rect 8251 5185 8263 5188
rect 8205 5179 8263 5185
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 8956 5157 8984 5188
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 10192 5188 10425 5216
rect 10192 5176 10198 5188
rect 10413 5185 10425 5188
rect 10459 5216 10471 5219
rect 10459 5188 11652 5216
rect 10459 5185 10471 5188
rect 10413 5179 10471 5185
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 992 5120 1777 5148
rect 992 5108 998 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 8941 5151 8999 5157
rect 8941 5117 8953 5151
rect 8987 5148 8999 5151
rect 9490 5148 9496 5160
rect 8987 5120 9496 5148
rect 8987 5117 8999 5120
rect 8941 5111 8999 5117
rect 9490 5108 9496 5120
rect 9548 5148 9554 5160
rect 10042 5148 10048 5160
rect 9548 5120 10048 5148
rect 9548 5108 9554 5120
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 10505 5151 10563 5157
rect 10505 5117 10517 5151
rect 10551 5117 10563 5151
rect 10505 5111 10563 5117
rect 6086 5040 6092 5092
rect 6144 5080 6150 5092
rect 9217 5083 9275 5089
rect 9217 5080 9229 5083
rect 6144 5052 9229 5080
rect 6144 5040 6150 5052
rect 9217 5049 9229 5052
rect 9263 5049 9275 5083
rect 10520 5080 10548 5111
rect 10594 5108 10600 5160
rect 10652 5108 10658 5160
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 10870 5148 10876 5160
rect 10735 5120 10876 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 10870 5108 10876 5120
rect 10928 5108 10934 5160
rect 11624 5148 11652 5188
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12437 5219 12495 5225
rect 12437 5216 12449 5219
rect 12308 5188 12449 5216
rect 12308 5176 12314 5188
rect 12437 5185 12449 5188
rect 12483 5185 12495 5219
rect 12437 5179 12495 5185
rect 13354 5176 13360 5228
rect 13412 5176 13418 5228
rect 13906 5176 13912 5228
rect 13964 5216 13970 5228
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 13964 5188 14381 5216
rect 13964 5176 13970 5188
rect 14369 5185 14381 5188
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 18693 5219 18751 5225
rect 18693 5185 18705 5219
rect 18739 5216 18751 5219
rect 19242 5216 19248 5228
rect 18739 5188 19248 5216
rect 18739 5185 18751 5188
rect 18693 5179 18751 5185
rect 19242 5176 19248 5188
rect 19300 5176 19306 5228
rect 11624 5120 18000 5148
rect 11974 5080 11980 5092
rect 10520 5052 11980 5080
rect 9217 5043 9275 5049
rect 11974 5040 11980 5052
rect 12032 5040 12038 5092
rect 12066 5040 12072 5092
rect 12124 5080 12130 5092
rect 13633 5083 13691 5089
rect 13633 5080 13645 5083
rect 12124 5052 13645 5080
rect 12124 5040 12130 5052
rect 13633 5049 13645 5052
rect 13679 5049 13691 5083
rect 13633 5043 13691 5049
rect 16574 5040 16580 5092
rect 16632 5080 16638 5092
rect 17865 5083 17923 5089
rect 17865 5080 17877 5083
rect 16632 5052 17877 5080
rect 16632 5040 16638 5052
rect 17865 5049 17877 5052
rect 17911 5049 17923 5083
rect 17865 5043 17923 5049
rect 8386 4972 8392 5024
rect 8444 4972 8450 5024
rect 12529 5015 12587 5021
rect 12529 4981 12541 5015
rect 12575 5012 12587 5015
rect 13446 5012 13452 5024
rect 12575 4984 13452 5012
rect 12575 4981 12587 4984
rect 12529 4975 12587 4981
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 13538 4972 13544 5024
rect 13596 5012 13602 5024
rect 14461 5015 14519 5021
rect 14461 5012 14473 5015
rect 13596 4984 14473 5012
rect 13596 4972 13602 4984
rect 14461 4981 14473 4984
rect 14507 4981 14519 5015
rect 14461 4975 14519 4981
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 16666 5012 16672 5024
rect 16347 4984 16672 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 17221 5015 17279 5021
rect 17221 5012 17233 5015
rect 17000 4984 17233 5012
rect 17000 4972 17006 4984
rect 17221 4981 17233 4984
rect 17267 4981 17279 5015
rect 17972 5012 18000 5120
rect 18598 5108 18604 5160
rect 18656 5148 18662 5160
rect 18877 5151 18935 5157
rect 18877 5148 18889 5151
rect 18656 5120 18889 5148
rect 18656 5108 18662 5120
rect 18877 5117 18889 5120
rect 18923 5117 18935 5151
rect 18877 5111 18935 5117
rect 19352 5080 19380 5256
rect 19444 5148 19472 5324
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 19886 5352 19892 5364
rect 19659 5324 19892 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 20438 5352 20444 5364
rect 19996 5324 20444 5352
rect 19996 5293 20024 5324
rect 20438 5312 20444 5324
rect 20496 5312 20502 5364
rect 25130 5312 25136 5364
rect 25188 5352 25194 5364
rect 25777 5355 25835 5361
rect 25777 5352 25789 5355
rect 25188 5324 25789 5352
rect 25188 5312 25194 5324
rect 25777 5321 25789 5324
rect 25823 5321 25835 5355
rect 25777 5315 25835 5321
rect 25866 5312 25872 5364
rect 25924 5352 25930 5364
rect 29365 5355 29423 5361
rect 29365 5352 29377 5355
rect 25924 5324 29377 5352
rect 25924 5312 25930 5324
rect 29365 5321 29377 5324
rect 29411 5321 29423 5355
rect 29365 5315 29423 5321
rect 30745 5355 30803 5361
rect 30745 5321 30757 5355
rect 30791 5352 30803 5355
rect 32858 5352 32864 5364
rect 30791 5324 32864 5352
rect 30791 5321 30803 5324
rect 30745 5315 30803 5321
rect 32858 5312 32864 5324
rect 32916 5312 32922 5364
rect 35342 5352 35348 5364
rect 35084 5324 35348 5352
rect 19981 5287 20039 5293
rect 19981 5253 19993 5287
rect 20027 5253 20039 5287
rect 19981 5247 20039 5253
rect 20073 5287 20131 5293
rect 20073 5253 20085 5287
rect 20119 5253 20131 5287
rect 20073 5247 20131 5253
rect 19518 5176 19524 5228
rect 19576 5216 19582 5228
rect 20088 5216 20116 5247
rect 20346 5244 20352 5296
rect 20404 5284 20410 5296
rect 26878 5284 26884 5296
rect 20404 5256 26884 5284
rect 20404 5244 20410 5256
rect 26878 5244 26884 5256
rect 26936 5244 26942 5296
rect 30009 5287 30067 5293
rect 26988 5256 29224 5284
rect 19576 5188 20116 5216
rect 20993 5219 21051 5225
rect 19576 5176 19582 5188
rect 20993 5185 21005 5219
rect 21039 5216 21051 5219
rect 21818 5216 21824 5228
rect 21039 5188 21824 5216
rect 21039 5185 21051 5188
rect 20993 5179 21051 5185
rect 21818 5176 21824 5188
rect 21876 5176 21882 5228
rect 22554 5176 22560 5228
rect 22612 5176 22618 5228
rect 23661 5219 23719 5225
rect 23661 5185 23673 5219
rect 23707 5216 23719 5219
rect 24210 5216 24216 5228
rect 23707 5188 24216 5216
rect 23707 5185 23719 5188
rect 23661 5179 23719 5185
rect 24210 5176 24216 5188
rect 24268 5176 24274 5228
rect 25593 5219 25651 5225
rect 25593 5185 25605 5219
rect 25639 5216 25651 5219
rect 26142 5216 26148 5228
rect 25639 5188 26148 5216
rect 25639 5185 25651 5188
rect 25593 5179 25651 5185
rect 26142 5176 26148 5188
rect 26200 5176 26206 5228
rect 20070 5148 20076 5160
rect 19444 5120 20076 5148
rect 20070 5108 20076 5120
rect 20128 5108 20134 5160
rect 20257 5151 20315 5157
rect 20257 5117 20269 5151
rect 20303 5148 20315 5151
rect 20898 5148 20904 5160
rect 20303 5120 20904 5148
rect 20303 5117 20315 5120
rect 20257 5111 20315 5117
rect 20898 5108 20904 5120
rect 20956 5108 20962 5160
rect 21174 5108 21180 5160
rect 21232 5108 21238 5160
rect 22462 5108 22468 5160
rect 22520 5148 22526 5160
rect 22741 5151 22799 5157
rect 22741 5148 22753 5151
rect 22520 5120 22753 5148
rect 22520 5108 22526 5120
rect 22741 5117 22753 5120
rect 22787 5117 22799 5151
rect 22741 5111 22799 5117
rect 23566 5108 23572 5160
rect 23624 5148 23630 5160
rect 23845 5151 23903 5157
rect 23845 5148 23857 5151
rect 23624 5120 23857 5148
rect 23624 5108 23630 5120
rect 23845 5117 23857 5120
rect 23891 5117 23903 5151
rect 23845 5111 23903 5117
rect 20990 5080 20996 5092
rect 19352 5052 20996 5080
rect 20990 5040 20996 5052
rect 21048 5040 21054 5092
rect 21082 5040 21088 5092
rect 21140 5080 21146 5092
rect 26988 5080 27016 5256
rect 29196 5228 29224 5256
rect 30009 5253 30021 5287
rect 30055 5253 30067 5287
rect 35084 5284 35112 5324
rect 35342 5312 35348 5324
rect 35400 5352 35406 5364
rect 35400 5324 36124 5352
rect 35400 5312 35406 5324
rect 35986 5284 35992 5296
rect 30009 5247 30067 5253
rect 31726 5256 35112 5284
rect 35176 5256 35992 5284
rect 27522 5176 27528 5228
rect 27580 5216 27586 5228
rect 28353 5219 28411 5225
rect 28353 5216 28365 5219
rect 27580 5188 28365 5216
rect 27580 5176 27586 5188
rect 28353 5185 28365 5188
rect 28399 5185 28411 5219
rect 28353 5179 28411 5185
rect 28445 5219 28503 5225
rect 28445 5185 28457 5219
rect 28491 5216 28503 5219
rect 28534 5216 28540 5228
rect 28491 5188 28540 5216
rect 28491 5185 28503 5188
rect 28445 5179 28503 5185
rect 21140 5052 27016 5080
rect 28368 5080 28396 5179
rect 28534 5176 28540 5188
rect 28592 5176 28598 5228
rect 29178 5176 29184 5228
rect 29236 5176 29242 5228
rect 30024 5216 30052 5247
rect 30653 5219 30711 5225
rect 30653 5216 30665 5219
rect 30024 5188 30665 5216
rect 28629 5151 28687 5157
rect 28629 5117 28641 5151
rect 28675 5148 28687 5151
rect 28718 5148 28724 5160
rect 28675 5120 28724 5148
rect 28675 5117 28687 5120
rect 28629 5111 28687 5117
rect 28718 5108 28724 5120
rect 28776 5108 28782 5160
rect 29086 5108 29092 5160
rect 29144 5148 29150 5160
rect 30024 5148 30052 5188
rect 30653 5185 30665 5188
rect 30699 5185 30711 5219
rect 30653 5179 30711 5185
rect 30834 5176 30840 5228
rect 30892 5176 30898 5228
rect 29144 5120 30052 5148
rect 29144 5108 29150 5120
rect 31726 5080 31754 5256
rect 31846 5176 31852 5228
rect 31904 5216 31910 5228
rect 32861 5219 32919 5225
rect 32861 5216 32873 5219
rect 31904 5188 32873 5216
rect 31904 5176 31910 5188
rect 32861 5185 32873 5188
rect 32907 5216 32919 5219
rect 33597 5219 33655 5225
rect 33597 5216 33609 5219
rect 32907 5188 33609 5216
rect 32907 5185 32919 5188
rect 32861 5179 32919 5185
rect 33597 5185 33609 5188
rect 33643 5216 33655 5219
rect 34238 5216 34244 5228
rect 33643 5188 34244 5216
rect 33643 5185 33655 5188
rect 33597 5179 33655 5185
rect 34238 5176 34244 5188
rect 34296 5216 34302 5228
rect 34333 5219 34391 5225
rect 34333 5216 34345 5219
rect 34296 5188 34345 5216
rect 34296 5176 34302 5188
rect 34333 5185 34345 5188
rect 34379 5185 34391 5219
rect 34333 5179 34391 5185
rect 34422 5176 34428 5228
rect 34480 5216 34486 5228
rect 35176 5225 35204 5256
rect 35986 5244 35992 5256
rect 36044 5244 36050 5296
rect 36096 5284 36124 5324
rect 39574 5312 39580 5364
rect 39632 5352 39638 5364
rect 40589 5355 40647 5361
rect 40589 5352 40601 5355
rect 39632 5324 40601 5352
rect 39632 5312 39638 5324
rect 40589 5321 40601 5324
rect 40635 5321 40647 5355
rect 40589 5315 40647 5321
rect 42797 5355 42855 5361
rect 42797 5321 42809 5355
rect 42843 5352 42855 5355
rect 43162 5352 43168 5364
rect 42843 5324 43168 5352
rect 42843 5321 42855 5324
rect 42797 5315 42855 5321
rect 43162 5312 43168 5324
rect 43220 5312 43226 5364
rect 43898 5312 43904 5364
rect 43956 5352 43962 5364
rect 53098 5352 53104 5364
rect 43956 5324 53104 5352
rect 43956 5312 43962 5324
rect 53098 5312 53104 5324
rect 53156 5312 53162 5364
rect 58253 5355 58311 5361
rect 58253 5321 58265 5355
rect 58299 5321 58311 5355
rect 58253 5315 58311 5321
rect 58268 5284 58296 5315
rect 36096 5256 58296 5284
rect 35161 5219 35219 5225
rect 34480 5188 35112 5216
rect 34480 5176 34486 5188
rect 33045 5151 33103 5157
rect 33045 5117 33057 5151
rect 33091 5148 33103 5151
rect 33091 5120 34928 5148
rect 33091 5117 33103 5120
rect 33045 5111 33103 5117
rect 28368 5052 31754 5080
rect 21140 5040 21146 5052
rect 33134 5040 33140 5092
rect 33192 5080 33198 5092
rect 34330 5080 34336 5092
rect 33192 5052 34336 5080
rect 33192 5040 33198 5052
rect 34330 5040 34336 5052
rect 34388 5040 34394 5092
rect 34517 5083 34575 5089
rect 34517 5049 34529 5083
rect 34563 5080 34575 5083
rect 34606 5080 34612 5092
rect 34563 5052 34612 5080
rect 34563 5049 34575 5052
rect 34517 5043 34575 5049
rect 34606 5040 34612 5052
rect 34664 5040 34670 5092
rect 34900 5080 34928 5120
rect 34974 5108 34980 5160
rect 35032 5108 35038 5160
rect 35084 5148 35112 5188
rect 35161 5185 35173 5219
rect 35207 5185 35219 5219
rect 35805 5219 35863 5225
rect 35805 5216 35817 5219
rect 35161 5179 35219 5185
rect 35268 5188 35817 5216
rect 35268 5148 35296 5188
rect 35805 5185 35817 5188
rect 35851 5185 35863 5219
rect 35805 5179 35863 5185
rect 36262 5176 36268 5228
rect 36320 5216 36326 5228
rect 37553 5219 37611 5225
rect 37553 5216 37565 5219
rect 36320 5188 37565 5216
rect 36320 5176 36326 5188
rect 37553 5185 37565 5188
rect 37599 5216 37611 5219
rect 38010 5216 38016 5228
rect 37599 5188 38016 5216
rect 37599 5185 37611 5188
rect 37553 5179 37611 5185
rect 38010 5176 38016 5188
rect 38068 5176 38074 5228
rect 38740 5219 38798 5225
rect 38740 5185 38752 5219
rect 38786 5216 38798 5219
rect 39114 5216 39120 5228
rect 38786 5188 39120 5216
rect 38786 5185 38798 5188
rect 38740 5179 38798 5185
rect 39114 5176 39120 5188
rect 39172 5176 39178 5228
rect 39206 5176 39212 5228
rect 39264 5216 39270 5228
rect 40405 5219 40463 5225
rect 40405 5216 40417 5219
rect 39264 5188 40417 5216
rect 39264 5176 39270 5188
rect 40405 5185 40417 5188
rect 40451 5185 40463 5219
rect 40405 5179 40463 5185
rect 40494 5176 40500 5228
rect 40552 5216 40558 5228
rect 41233 5219 41291 5225
rect 41233 5216 41245 5219
rect 40552 5188 41245 5216
rect 40552 5176 40558 5188
rect 41233 5185 41245 5188
rect 41279 5185 41291 5219
rect 41233 5179 41291 5185
rect 41874 5176 41880 5228
rect 41932 5216 41938 5228
rect 42705 5219 42763 5225
rect 42705 5216 42717 5219
rect 41932 5188 42717 5216
rect 41932 5176 41938 5188
rect 42705 5185 42717 5188
rect 42751 5185 42763 5219
rect 42705 5179 42763 5185
rect 42886 5176 42892 5228
rect 42944 5216 42950 5228
rect 43441 5219 43499 5225
rect 43441 5216 43453 5219
rect 42944 5188 43453 5216
rect 42944 5176 42950 5188
rect 43441 5185 43453 5188
rect 43487 5185 43499 5219
rect 43441 5179 43499 5185
rect 44174 5176 44180 5228
rect 44232 5176 44238 5228
rect 44542 5176 44548 5228
rect 44600 5216 44606 5228
rect 44913 5219 44971 5225
rect 44913 5216 44925 5219
rect 44600 5188 44925 5216
rect 44600 5176 44606 5188
rect 44913 5185 44925 5188
rect 44959 5185 44971 5219
rect 44913 5179 44971 5185
rect 45646 5176 45652 5228
rect 45704 5216 45710 5228
rect 45833 5219 45891 5225
rect 45833 5216 45845 5219
rect 45704 5188 45845 5216
rect 45704 5176 45710 5188
rect 45833 5185 45845 5188
rect 45879 5185 45891 5219
rect 45833 5179 45891 5185
rect 46934 5176 46940 5228
rect 46992 5216 46998 5228
rect 48501 5219 48559 5225
rect 48501 5216 48513 5219
rect 46992 5188 48513 5216
rect 46992 5176 46998 5188
rect 48501 5185 48513 5188
rect 48547 5185 48559 5219
rect 48757 5219 48815 5225
rect 48757 5216 48769 5219
rect 48501 5179 48559 5185
rect 48608 5188 48769 5216
rect 35084 5120 35296 5148
rect 35342 5108 35348 5160
rect 35400 5148 35406 5160
rect 35400 5120 35664 5148
rect 35400 5108 35406 5120
rect 35434 5080 35440 5092
rect 34900 5052 35440 5080
rect 35434 5040 35440 5052
rect 35492 5040 35498 5092
rect 35636 5080 35664 5120
rect 35710 5108 35716 5160
rect 35768 5148 35774 5160
rect 35989 5151 36047 5157
rect 35989 5148 36001 5151
rect 35768 5120 36001 5148
rect 35768 5108 35774 5120
rect 35989 5117 36001 5120
rect 36035 5117 36047 5151
rect 35989 5111 36047 5117
rect 36998 5108 37004 5160
rect 37056 5148 37062 5160
rect 38473 5151 38531 5157
rect 38473 5148 38485 5151
rect 37056 5120 38485 5148
rect 37056 5108 37062 5120
rect 38473 5117 38485 5120
rect 38519 5117 38531 5151
rect 38473 5111 38531 5117
rect 40586 5108 40592 5160
rect 40644 5148 40650 5160
rect 46017 5151 46075 5157
rect 46017 5148 46029 5151
rect 40644 5120 46029 5148
rect 40644 5108 40650 5120
rect 46017 5117 46029 5120
rect 46063 5117 46075 5151
rect 46017 5111 46075 5117
rect 46566 5108 46572 5160
rect 46624 5148 46630 5160
rect 48608 5148 48636 5188
rect 48757 5185 48769 5188
rect 48803 5185 48815 5219
rect 48757 5179 48815 5185
rect 58066 5176 58072 5228
rect 58124 5176 58130 5228
rect 46624 5120 48636 5148
rect 46624 5108 46630 5120
rect 37734 5080 37740 5092
rect 35636 5052 37740 5080
rect 37734 5040 37740 5052
rect 37792 5040 37798 5092
rect 41230 5040 41236 5092
rect 41288 5080 41294 5092
rect 43625 5083 43683 5089
rect 43625 5080 43637 5083
rect 41288 5052 43637 5080
rect 41288 5040 41294 5052
rect 43625 5049 43637 5052
rect 43671 5049 43683 5083
rect 43625 5043 43683 5049
rect 20714 5012 20720 5024
rect 17972 4984 20720 5012
rect 17221 4975 17279 4981
rect 20714 4972 20720 4984
rect 20772 4972 20778 5024
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 23474 5012 23480 5024
rect 20956 4984 23480 5012
rect 20956 4972 20962 4984
rect 23474 4972 23480 4984
rect 23532 5012 23538 5024
rect 23842 5012 23848 5024
rect 23532 4984 23848 5012
rect 23532 4972 23538 4984
rect 23842 4972 23848 4984
rect 23900 4972 23906 5024
rect 26234 4972 26240 5024
rect 26292 5012 26298 5024
rect 26513 5015 26571 5021
rect 26513 5012 26525 5015
rect 26292 4984 26525 5012
rect 26292 4972 26298 4984
rect 26513 4981 26525 4984
rect 26559 4981 26571 5015
rect 26513 4975 26571 4981
rect 27522 4972 27528 5024
rect 27580 5012 27586 5024
rect 27985 5015 28043 5021
rect 27985 5012 27997 5015
rect 27580 4984 27997 5012
rect 27580 4972 27586 4984
rect 27985 4981 27997 4984
rect 28031 4981 28043 5015
rect 27985 4975 28043 4981
rect 28166 4972 28172 5024
rect 28224 5012 28230 5024
rect 30101 5015 30159 5021
rect 30101 5012 30113 5015
rect 28224 4984 30113 5012
rect 28224 4972 28230 4984
rect 30101 4981 30113 4984
rect 30147 4981 30159 5015
rect 30101 4975 30159 4981
rect 33689 5015 33747 5021
rect 33689 4981 33701 5015
rect 33735 5012 33747 5015
rect 34790 5012 34796 5024
rect 33735 4984 34796 5012
rect 33735 4981 33747 4984
rect 33689 4975 33747 4981
rect 34790 4972 34796 4984
rect 34848 4972 34854 5024
rect 35345 5015 35403 5021
rect 35345 4981 35357 5015
rect 35391 5012 35403 5015
rect 35986 5012 35992 5024
rect 35391 4984 35992 5012
rect 35391 4981 35403 4984
rect 35345 4975 35403 4981
rect 35986 4972 35992 4984
rect 36044 4972 36050 5024
rect 37645 5015 37703 5021
rect 37645 4981 37657 5015
rect 37691 5012 37703 5015
rect 38654 5012 38660 5024
rect 37691 4984 38660 5012
rect 37691 4981 37703 4984
rect 37645 4975 37703 4981
rect 38654 4972 38660 4984
rect 38712 4972 38718 5024
rect 38838 4972 38844 5024
rect 38896 5012 38902 5024
rect 39853 5015 39911 5021
rect 39853 5012 39865 5015
rect 38896 4984 39865 5012
rect 38896 4972 38902 4984
rect 39853 4981 39865 4984
rect 39899 4981 39911 5015
rect 39853 4975 39911 4981
rect 41138 4972 41144 5024
rect 41196 5012 41202 5024
rect 41325 5015 41383 5021
rect 41325 5012 41337 5015
rect 41196 4984 41337 5012
rect 41196 4972 41202 4984
rect 41325 4981 41337 4984
rect 41371 4981 41383 5015
rect 41325 4975 41383 4981
rect 43070 4972 43076 5024
rect 43128 5012 43134 5024
rect 44269 5015 44327 5021
rect 44269 5012 44281 5015
rect 43128 4984 44281 5012
rect 43128 4972 43134 4984
rect 44269 4981 44281 4984
rect 44315 4981 44327 5015
rect 44269 4975 44327 4981
rect 45002 4972 45008 5024
rect 45060 4972 45066 5024
rect 49881 5015 49939 5021
rect 49881 4981 49893 5015
rect 49927 5012 49939 5015
rect 51074 5012 51080 5024
rect 49927 4984 51080 5012
rect 49927 4981 49939 4984
rect 49881 4975 49939 4981
rect 51074 4972 51080 4984
rect 51132 4972 51138 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 8110 4768 8116 4820
rect 8168 4808 8174 4820
rect 9677 4811 9735 4817
rect 9677 4808 9689 4811
rect 8168 4780 9689 4808
rect 8168 4768 8174 4780
rect 9677 4777 9689 4780
rect 9723 4777 9735 4811
rect 9677 4771 9735 4777
rect 11149 4811 11207 4817
rect 11149 4777 11161 4811
rect 11195 4808 11207 4811
rect 11238 4808 11244 4820
rect 11195 4780 11244 4808
rect 11195 4777 11207 4780
rect 11149 4771 11207 4777
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 16114 4768 16120 4820
rect 16172 4808 16178 4820
rect 19334 4808 19340 4820
rect 16172 4780 19340 4808
rect 16172 4768 16178 4780
rect 19334 4768 19340 4780
rect 19392 4768 19398 4820
rect 19429 4811 19487 4817
rect 19429 4777 19441 4811
rect 19475 4808 19487 4811
rect 19518 4808 19524 4820
rect 19475 4780 19524 4808
rect 19475 4777 19487 4780
rect 19429 4771 19487 4777
rect 19518 4768 19524 4780
rect 19576 4768 19582 4820
rect 19812 4780 21404 4808
rect 7098 4700 7104 4752
rect 7156 4700 7162 4752
rect 8573 4743 8631 4749
rect 8573 4709 8585 4743
rect 8619 4740 8631 4743
rect 10965 4743 11023 4749
rect 10965 4740 10977 4743
rect 8619 4712 10977 4740
rect 8619 4709 8631 4712
rect 8573 4703 8631 4709
rect 10965 4709 10977 4712
rect 11011 4709 11023 4743
rect 10965 4703 11023 4709
rect 13446 4700 13452 4752
rect 13504 4700 13510 4752
rect 13633 4743 13691 4749
rect 13633 4709 13645 4743
rect 13679 4740 13691 4743
rect 13679 4712 14504 4740
rect 13679 4709 13691 4712
rect 13633 4703 13691 4709
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4672 6331 4675
rect 9766 4672 9772 4684
rect 6319 4644 9772 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 9858 4632 9864 4684
rect 9916 4632 9922 4684
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4672 10011 4675
rect 13173 4675 13231 4681
rect 9999 4644 13124 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 7006 4604 7012 4616
rect 6963 4576 7012 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 9674 4604 9680 4616
rect 8435 4576 9680 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 10042 4564 10048 4616
rect 10100 4564 10106 4616
rect 10137 4607 10195 4613
rect 10137 4573 10149 4607
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 5902 4496 5908 4548
rect 5960 4536 5966 4548
rect 6089 4539 6147 4545
rect 6089 4536 6101 4539
rect 5960 4508 6101 4536
rect 5960 4496 5966 4508
rect 6089 4505 6101 4508
rect 6135 4505 6147 4539
rect 6089 4499 6147 4505
rect 7653 4539 7711 4545
rect 7653 4505 7665 4539
rect 7699 4536 7711 4539
rect 8294 4536 8300 4548
rect 7699 4508 8300 4536
rect 7699 4505 7711 4508
rect 7653 4499 7711 4505
rect 8294 4496 8300 4508
rect 8352 4496 8358 4548
rect 8570 4496 8576 4548
rect 8628 4536 8634 4548
rect 10152 4536 10180 4567
rect 10594 4564 10600 4616
rect 10652 4604 10658 4616
rect 10689 4607 10747 4613
rect 10689 4604 10701 4607
rect 10652 4576 10701 4604
rect 10652 4564 10658 4576
rect 10689 4573 10701 4576
rect 10735 4573 10747 4607
rect 10689 4567 10747 4573
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4604 12035 4607
rect 12710 4604 12716 4616
rect 12023 4576 12716 4604
rect 12023 4573 12035 4576
rect 11977 4567 12035 4573
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 13096 4604 13124 4644
rect 13173 4641 13185 4675
rect 13219 4672 13231 4675
rect 13354 4672 13360 4684
rect 13219 4644 13360 4672
rect 13219 4641 13231 4644
rect 13173 4635 13231 4641
rect 13354 4632 13360 4644
rect 13412 4672 13418 4684
rect 14277 4675 14335 4681
rect 14277 4672 14289 4675
rect 13412 4644 14289 4672
rect 13412 4632 13418 4644
rect 14277 4641 14289 4644
rect 14323 4641 14335 4675
rect 14476 4672 14504 4712
rect 14550 4700 14556 4752
rect 14608 4700 14614 4752
rect 19610 4740 19616 4752
rect 17512 4712 19616 4740
rect 15286 4672 15292 4684
rect 14476 4644 15292 4672
rect 14277 4635 14335 4641
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 15194 4604 15200 4616
rect 13096 4576 15200 4604
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 15378 4564 15384 4616
rect 15436 4604 15442 4616
rect 17037 4607 17095 4613
rect 15436 4576 16528 4604
rect 15436 4564 15442 4576
rect 8628 4508 10180 4536
rect 11793 4539 11851 4545
rect 8628 4496 8634 4508
rect 11793 4505 11805 4539
rect 11839 4536 11851 4539
rect 12529 4539 12587 4545
rect 11839 4508 12020 4536
rect 11839 4505 11851 4508
rect 11793 4499 11851 4505
rect 11992 4480 12020 4508
rect 12529 4505 12541 4539
rect 12575 4536 12587 4539
rect 13078 4536 13084 4548
rect 12575 4508 13084 4536
rect 12575 4505 12587 4508
rect 12529 4499 12587 4505
rect 13078 4496 13084 4508
rect 13136 4496 13142 4548
rect 14182 4536 14188 4548
rect 13556 4508 14188 4536
rect 7558 4428 7564 4480
rect 7616 4468 7622 4480
rect 7745 4471 7803 4477
rect 7745 4468 7757 4471
rect 7616 4440 7757 4468
rect 7616 4428 7622 4440
rect 7745 4437 7757 4440
rect 7791 4437 7803 4471
rect 7745 4431 7803 4437
rect 11974 4428 11980 4480
rect 12032 4428 12038 4480
rect 12621 4471 12679 4477
rect 12621 4437 12633 4471
rect 12667 4468 12679 4471
rect 13556 4468 13584 4508
rect 14182 4496 14188 4508
rect 14240 4496 14246 4548
rect 15286 4496 15292 4548
rect 15344 4536 15350 4548
rect 15657 4539 15715 4545
rect 15657 4536 15669 4539
rect 15344 4508 15669 4536
rect 15344 4496 15350 4508
rect 15657 4505 15669 4508
rect 15703 4505 15715 4539
rect 16500 4536 16528 4576
rect 17037 4573 17049 4607
rect 17083 4604 17095 4607
rect 17218 4604 17224 4616
rect 17083 4576 17224 4604
rect 17083 4573 17095 4576
rect 17037 4567 17095 4573
rect 17218 4564 17224 4576
rect 17276 4564 17282 4616
rect 17512 4613 17540 4712
rect 19610 4700 19616 4712
rect 19668 4700 19674 4752
rect 19812 4672 19840 4780
rect 20070 4700 20076 4752
rect 20128 4740 20134 4752
rect 21082 4740 21088 4752
rect 20128 4712 21088 4740
rect 20128 4700 20134 4712
rect 21082 4700 21088 4712
rect 21140 4700 21146 4752
rect 17604 4644 19840 4672
rect 19981 4675 20039 4681
rect 17497 4607 17555 4613
rect 17497 4573 17509 4607
rect 17543 4573 17555 4607
rect 17497 4567 17555 4573
rect 17604 4536 17632 4644
rect 19981 4641 19993 4675
rect 20027 4641 20039 4675
rect 19981 4635 20039 4641
rect 18417 4607 18475 4613
rect 18417 4573 18429 4607
rect 18463 4604 18475 4607
rect 19058 4604 19064 4616
rect 18463 4576 19064 4604
rect 18463 4573 18475 4576
rect 18417 4567 18475 4573
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19996 4604 20024 4635
rect 21266 4632 21272 4684
rect 21324 4632 21330 4684
rect 21376 4672 21404 4780
rect 33502 4768 33508 4820
rect 33560 4808 33566 4820
rect 36354 4808 36360 4820
rect 33560 4780 36360 4808
rect 33560 4768 33566 4780
rect 36354 4768 36360 4780
rect 36412 4808 36418 4820
rect 37093 4811 37151 4817
rect 37093 4808 37105 4811
rect 36412 4780 37105 4808
rect 36412 4768 36418 4780
rect 37093 4777 37105 4780
rect 37139 4777 37151 4811
rect 37093 4771 37151 4777
rect 37366 4768 37372 4820
rect 37424 4808 37430 4820
rect 38838 4808 38844 4820
rect 37424 4780 38844 4808
rect 37424 4768 37430 4780
rect 38838 4768 38844 4780
rect 38896 4768 38902 4820
rect 39114 4768 39120 4820
rect 39172 4768 39178 4820
rect 40218 4768 40224 4820
rect 40276 4768 40282 4820
rect 40678 4768 40684 4820
rect 40736 4808 40742 4820
rect 41693 4811 41751 4817
rect 41693 4808 41705 4811
rect 40736 4780 41705 4808
rect 40736 4768 40742 4780
rect 41693 4777 41705 4780
rect 41739 4777 41751 4811
rect 41693 4771 41751 4777
rect 42996 4780 51074 4808
rect 29638 4740 29644 4752
rect 23400 4712 29644 4740
rect 23400 4672 23428 4712
rect 29638 4700 29644 4712
rect 29696 4700 29702 4752
rect 32309 4743 32367 4749
rect 32309 4709 32321 4743
rect 32355 4740 32367 4743
rect 32355 4712 33364 4740
rect 32355 4709 32367 4712
rect 32309 4703 32367 4709
rect 21376 4644 23428 4672
rect 23842 4632 23848 4684
rect 23900 4632 23906 4684
rect 24946 4672 24952 4684
rect 23952 4644 24952 4672
rect 20254 4604 20260 4616
rect 19392 4576 20260 4604
rect 19392 4564 19398 4576
rect 20254 4564 20260 4576
rect 20312 4564 20318 4616
rect 22370 4564 22376 4616
rect 22428 4564 22434 4616
rect 23661 4607 23719 4613
rect 23661 4573 23673 4607
rect 23707 4604 23719 4607
rect 23952 4604 23980 4644
rect 24946 4632 24952 4644
rect 25004 4632 25010 4684
rect 27614 4632 27620 4684
rect 27672 4632 27678 4684
rect 28718 4672 28724 4684
rect 28000 4644 28724 4672
rect 23707 4576 23980 4604
rect 23707 4573 23719 4576
rect 23661 4567 23719 4573
rect 24670 4564 24676 4616
rect 24728 4564 24734 4616
rect 26326 4564 26332 4616
rect 26384 4604 26390 4616
rect 26513 4607 26571 4613
rect 26513 4604 26525 4607
rect 26384 4576 26525 4604
rect 26384 4564 26390 4576
rect 26513 4573 26525 4576
rect 26559 4573 26571 4607
rect 26513 4567 26571 4573
rect 27798 4564 27804 4616
rect 27856 4564 27862 4616
rect 16500 4508 17632 4536
rect 17773 4539 17831 4545
rect 15657 4499 15715 4505
rect 17773 4505 17785 4539
rect 17819 4536 17831 4539
rect 18046 4536 18052 4548
rect 17819 4508 18052 4536
rect 17819 4505 17831 4508
rect 17773 4499 17831 4505
rect 18046 4496 18052 4508
rect 18104 4496 18110 4548
rect 18693 4539 18751 4545
rect 18693 4505 18705 4539
rect 18739 4536 18751 4539
rect 19150 4536 19156 4548
rect 18739 4508 19156 4536
rect 18739 4505 18751 4508
rect 18693 4499 18751 4505
rect 19150 4496 19156 4508
rect 19208 4496 19214 4548
rect 19242 4496 19248 4548
rect 19300 4536 19306 4548
rect 20346 4536 20352 4548
rect 19300 4508 20352 4536
rect 19300 4496 19306 4508
rect 20346 4496 20352 4508
rect 20404 4496 20410 4548
rect 20993 4539 21051 4545
rect 20993 4505 21005 4539
rect 21039 4536 21051 4539
rect 22554 4536 22560 4548
rect 21039 4508 22560 4536
rect 21039 4505 21051 4508
rect 20993 4499 21051 4505
rect 22554 4496 22560 4508
rect 22612 4496 22618 4548
rect 22649 4539 22707 4545
rect 22649 4505 22661 4539
rect 22695 4536 22707 4539
rect 22738 4536 22744 4548
rect 22695 4508 22744 4536
rect 22695 4505 22707 4508
rect 22649 4499 22707 4505
rect 22738 4496 22744 4508
rect 22796 4496 22802 4548
rect 23934 4496 23940 4548
rect 23992 4536 23998 4548
rect 28000 4536 28028 4644
rect 28718 4632 28724 4644
rect 28776 4672 28782 4684
rect 28813 4675 28871 4681
rect 28813 4672 28825 4675
rect 28776 4644 28825 4672
rect 28776 4632 28782 4644
rect 28813 4641 28825 4644
rect 28859 4641 28871 4675
rect 28813 4635 28871 4641
rect 29454 4632 29460 4684
rect 29512 4672 29518 4684
rect 32858 4672 32864 4684
rect 29512 4644 32864 4672
rect 29512 4632 29518 4644
rect 32858 4632 32864 4644
rect 32916 4632 32922 4684
rect 33336 4672 33364 4712
rect 36906 4700 36912 4752
rect 36964 4740 36970 4752
rect 37826 4740 37832 4752
rect 36964 4712 37832 4740
rect 36964 4700 36970 4712
rect 37826 4700 37832 4712
rect 37884 4700 37890 4752
rect 38010 4700 38016 4752
rect 38068 4740 38074 4752
rect 38068 4712 39160 4740
rect 38068 4700 38074 4712
rect 39132 4684 39160 4712
rect 38749 4675 38807 4681
rect 38749 4672 38761 4675
rect 33336 4644 33732 4672
rect 28537 4607 28595 4613
rect 28537 4573 28549 4607
rect 28583 4604 28595 4607
rect 28994 4604 29000 4616
rect 28583 4576 29000 4604
rect 28583 4573 28595 4576
rect 28537 4567 28595 4573
rect 28994 4564 29000 4576
rect 29052 4564 29058 4616
rect 29178 4564 29184 4616
rect 29236 4604 29242 4616
rect 32677 4607 32735 4613
rect 32677 4604 32689 4607
rect 29236 4576 32689 4604
rect 29236 4564 29242 4576
rect 32677 4573 32689 4576
rect 32723 4573 32735 4607
rect 32677 4567 32735 4573
rect 32769 4607 32827 4613
rect 32769 4573 32781 4607
rect 32815 4604 32827 4607
rect 32950 4604 32956 4616
rect 32815 4576 32956 4604
rect 32815 4573 32827 4576
rect 32769 4567 32827 4573
rect 23992 4508 28028 4536
rect 23992 4496 23998 4508
rect 30006 4496 30012 4548
rect 30064 4496 30070 4548
rect 30193 4539 30251 4545
rect 30193 4505 30205 4539
rect 30239 4536 30251 4539
rect 30282 4536 30288 4548
rect 30239 4508 30288 4536
rect 30239 4505 30251 4508
rect 30193 4499 30251 4505
rect 30282 4496 30288 4508
rect 30340 4496 30346 4548
rect 32692 4536 32720 4567
rect 32950 4564 32956 4576
rect 33008 4564 33014 4616
rect 33704 4613 33732 4644
rect 37752 4644 38761 4672
rect 37752 4616 37780 4644
rect 38749 4641 38761 4644
rect 38795 4641 38807 4675
rect 38749 4635 38807 4641
rect 39114 4632 39120 4684
rect 39172 4632 39178 4684
rect 41046 4632 41052 4684
rect 41104 4672 41110 4684
rect 41104 4644 42656 4672
rect 41104 4632 41110 4644
rect 33597 4607 33655 4613
rect 33597 4573 33609 4607
rect 33643 4573 33655 4607
rect 33597 4567 33655 4573
rect 33689 4607 33747 4613
rect 33689 4573 33701 4607
rect 33735 4573 33747 4607
rect 33689 4567 33747 4573
rect 33134 4536 33140 4548
rect 31726 4508 32628 4536
rect 32692 4508 33140 4536
rect 12667 4440 13584 4468
rect 12667 4437 12679 4440
rect 12621 4431 12679 4437
rect 14734 4428 14740 4480
rect 14792 4428 14798 4480
rect 14826 4428 14832 4480
rect 14884 4468 14890 4480
rect 19797 4471 19855 4477
rect 19797 4468 19809 4471
rect 14884 4440 19809 4468
rect 14884 4428 14890 4440
rect 19797 4437 19809 4440
rect 19843 4437 19855 4471
rect 19797 4431 19855 4437
rect 19889 4471 19947 4477
rect 19889 4437 19901 4471
rect 19935 4468 19947 4471
rect 20438 4468 20444 4480
rect 19935 4440 20444 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 20438 4428 20444 4440
rect 20496 4428 20502 4480
rect 20622 4428 20628 4480
rect 20680 4428 20686 4480
rect 21085 4471 21143 4477
rect 21085 4437 21097 4471
rect 21131 4468 21143 4471
rect 21174 4468 21180 4480
rect 21131 4440 21180 4468
rect 21131 4437 21143 4440
rect 21085 4431 21143 4437
rect 21174 4428 21180 4440
rect 21232 4428 21238 4480
rect 23293 4471 23351 4477
rect 23293 4437 23305 4471
rect 23339 4468 23351 4471
rect 23474 4468 23480 4480
rect 23339 4440 23480 4468
rect 23339 4437 23351 4440
rect 23293 4431 23351 4437
rect 23474 4428 23480 4440
rect 23532 4428 23538 4480
rect 23750 4428 23756 4480
rect 23808 4428 23814 4480
rect 26878 4428 26884 4480
rect 26936 4468 26942 4480
rect 26973 4471 27031 4477
rect 26973 4468 26985 4471
rect 26936 4440 26985 4468
rect 26936 4428 26942 4440
rect 26973 4437 26985 4440
rect 27019 4437 27031 4471
rect 26973 4431 27031 4437
rect 27985 4471 28043 4477
rect 27985 4437 27997 4471
rect 28031 4468 28043 4471
rect 28534 4468 28540 4480
rect 28031 4440 28540 4468
rect 28031 4437 28043 4440
rect 27985 4431 28043 4437
rect 28534 4428 28540 4440
rect 28592 4428 28598 4480
rect 28718 4428 28724 4480
rect 28776 4468 28782 4480
rect 31726 4468 31754 4508
rect 28776 4440 31754 4468
rect 32600 4468 32628 4508
rect 33134 4496 33140 4508
rect 33192 4496 33198 4548
rect 33612 4536 33640 4567
rect 34514 4564 34520 4616
rect 34572 4604 34578 4616
rect 35713 4607 35771 4613
rect 35713 4604 35725 4607
rect 34572 4576 35725 4604
rect 34572 4564 34578 4576
rect 35713 4573 35725 4576
rect 35759 4604 35771 4607
rect 36998 4604 37004 4616
rect 35759 4576 37004 4604
rect 35759 4573 35771 4576
rect 35713 4567 35771 4573
rect 36998 4564 37004 4576
rect 37056 4564 37062 4616
rect 37734 4564 37740 4616
rect 37792 4564 37798 4616
rect 37826 4564 37832 4616
rect 37884 4564 37890 4616
rect 38930 4564 38936 4616
rect 38988 4564 38994 4616
rect 40034 4564 40040 4616
rect 40092 4564 40098 4616
rect 40218 4564 40224 4616
rect 40276 4604 40282 4616
rect 41509 4607 41567 4613
rect 41509 4604 41521 4607
rect 40276 4576 41521 4604
rect 40276 4564 40282 4576
rect 41509 4573 41521 4576
rect 41555 4573 41567 4607
rect 41509 4567 41567 4573
rect 33778 4536 33784 4548
rect 33612 4508 33784 4536
rect 33778 4496 33784 4508
rect 33836 4496 33842 4548
rect 34054 4496 34060 4548
rect 34112 4536 34118 4548
rect 34422 4536 34428 4548
rect 34112 4508 34428 4536
rect 34112 4496 34118 4508
rect 34422 4496 34428 4508
rect 34480 4536 34486 4548
rect 34977 4539 35035 4545
rect 34977 4536 34989 4539
rect 34480 4508 34989 4536
rect 34480 4496 34486 4508
rect 34977 4505 34989 4508
rect 35023 4505 35035 4539
rect 34977 4499 35035 4505
rect 35161 4539 35219 4545
rect 35161 4505 35173 4539
rect 35207 4536 35219 4539
rect 35342 4536 35348 4548
rect 35207 4508 35348 4536
rect 35207 4505 35219 4508
rect 35161 4499 35219 4505
rect 35342 4496 35348 4508
rect 35400 4496 35406 4548
rect 35986 4545 35992 4548
rect 35980 4536 35992 4545
rect 35947 4508 35992 4536
rect 35980 4499 35992 4508
rect 35986 4496 35992 4499
rect 36044 4496 36050 4548
rect 36354 4496 36360 4548
rect 36412 4536 36418 4548
rect 39022 4536 39028 4548
rect 36412 4508 39028 4536
rect 36412 4496 36418 4508
rect 39022 4496 39028 4508
rect 39080 4496 39086 4548
rect 40862 4496 40868 4548
rect 40920 4496 40926 4548
rect 33502 4468 33508 4480
rect 32600 4440 33508 4468
rect 28776 4428 28782 4440
rect 33502 4428 33508 4440
rect 33560 4428 33566 4480
rect 33594 4428 33600 4480
rect 33652 4468 33658 4480
rect 33873 4471 33931 4477
rect 33873 4468 33885 4471
rect 33652 4440 33885 4468
rect 33652 4428 33658 4440
rect 33873 4437 33885 4440
rect 33919 4437 33931 4471
rect 33873 4431 33931 4437
rect 36262 4428 36268 4480
rect 36320 4468 36326 4480
rect 36722 4468 36728 4480
rect 36320 4440 36728 4468
rect 36320 4428 36326 4440
rect 36722 4428 36728 4440
rect 36780 4428 36786 4480
rect 38010 4428 38016 4480
rect 38068 4428 38074 4480
rect 38838 4428 38844 4480
rect 38896 4468 38902 4480
rect 40957 4471 41015 4477
rect 40957 4468 40969 4471
rect 38896 4440 40969 4468
rect 38896 4428 38902 4440
rect 40957 4437 40969 4440
rect 41003 4437 41015 4471
rect 42628 4468 42656 4644
rect 42702 4564 42708 4616
rect 42760 4564 42766 4616
rect 42853 4607 42911 4613
rect 42853 4573 42865 4607
rect 42899 4604 42911 4607
rect 42996 4604 43024 4780
rect 43254 4700 43260 4752
rect 43312 4740 43318 4752
rect 44453 4743 44511 4749
rect 44453 4740 44465 4743
rect 43312 4712 44465 4740
rect 43312 4700 43318 4712
rect 44453 4709 44465 4712
rect 44499 4709 44511 4743
rect 44453 4703 44511 4709
rect 45462 4700 45468 4752
rect 45520 4700 45526 4752
rect 51046 4740 51074 4780
rect 56686 4768 56692 4820
rect 56744 4808 56750 4820
rect 58253 4811 58311 4817
rect 58253 4808 58265 4811
rect 56744 4780 58265 4808
rect 56744 4768 56750 4780
rect 58253 4777 58265 4780
rect 58299 4777 58311 4811
rect 58253 4771 58311 4777
rect 51350 4740 51356 4752
rect 51046 4712 51356 4740
rect 51350 4700 51356 4712
rect 51408 4700 51414 4752
rect 46201 4675 46259 4681
rect 46201 4641 46213 4675
rect 46247 4641 46259 4675
rect 46201 4635 46259 4641
rect 42899 4576 43024 4604
rect 42899 4573 42911 4576
rect 42853 4567 42911 4573
rect 43070 4564 43076 4616
rect 43128 4564 43134 4616
rect 43211 4607 43269 4613
rect 43211 4573 43223 4607
rect 43257 4604 43269 4607
rect 43438 4604 43444 4616
rect 43257 4576 43444 4604
rect 43257 4573 43269 4576
rect 43211 4567 43269 4573
rect 43438 4564 43444 4576
rect 43496 4564 43502 4616
rect 43898 4564 43904 4616
rect 43956 4564 43962 4616
rect 43990 4564 43996 4616
rect 44048 4604 44054 4616
rect 44274 4607 44332 4613
rect 44274 4604 44286 4607
rect 44048 4576 44286 4604
rect 44048 4564 44054 4576
rect 44274 4573 44286 4576
rect 44320 4573 44332 4607
rect 46216 4604 46244 4635
rect 49602 4632 49608 4684
rect 49660 4672 49666 4684
rect 50893 4675 50951 4681
rect 50893 4672 50905 4675
rect 49660 4644 50905 4672
rect 49660 4632 49666 4644
rect 50893 4641 50905 4644
rect 50939 4641 50951 4675
rect 50893 4635 50951 4641
rect 44274 4567 44332 4573
rect 44376 4576 46244 4604
rect 42978 4496 42984 4548
rect 43036 4496 43042 4548
rect 44085 4539 44143 4545
rect 43088 4508 43484 4536
rect 43088 4468 43116 4508
rect 42628 4440 43116 4468
rect 40957 4431 41015 4437
rect 43346 4428 43352 4480
rect 43404 4428 43410 4480
rect 43456 4468 43484 4508
rect 44085 4505 44097 4539
rect 44131 4505 44143 4539
rect 44085 4499 44143 4505
rect 44177 4539 44235 4545
rect 44177 4505 44189 4539
rect 44223 4536 44235 4539
rect 44376 4536 44404 4576
rect 51074 4564 51080 4616
rect 51132 4564 51138 4616
rect 58069 4607 58127 4613
rect 58069 4573 58081 4607
rect 58115 4604 58127 4607
rect 58802 4604 58808 4616
rect 58115 4576 58808 4604
rect 58115 4573 58127 4576
rect 58069 4567 58127 4573
rect 58802 4564 58808 4576
rect 58860 4564 58866 4616
rect 44223 4508 44404 4536
rect 44223 4505 44235 4508
rect 44177 4499 44235 4505
rect 44100 4468 44128 4499
rect 44450 4496 44456 4548
rect 44508 4536 44514 4548
rect 45281 4539 45339 4545
rect 45281 4536 45293 4539
rect 44508 4508 45293 4536
rect 44508 4496 44514 4508
rect 45281 4505 45293 4508
rect 45327 4505 45339 4539
rect 45281 4499 45339 4505
rect 46014 4496 46020 4548
rect 46072 4496 46078 4548
rect 43456 4440 44128 4468
rect 51261 4471 51319 4477
rect 51261 4437 51273 4471
rect 51307 4468 51319 4471
rect 53742 4468 53748 4480
rect 51307 4440 53748 4468
rect 51307 4437 51319 4440
rect 51261 4431 51319 4437
rect 53742 4428 53748 4440
rect 53800 4428 53806 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 8846 4264 8852 4276
rect 7576 4236 8852 4264
rect 5813 4199 5871 4205
rect 5813 4165 5825 4199
rect 5859 4196 5871 4199
rect 6454 4196 6460 4208
rect 5859 4168 6460 4196
rect 5859 4165 5871 4168
rect 5813 4159 5871 4165
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 6641 4199 6699 4205
rect 6641 4165 6653 4199
rect 6687 4196 6699 4199
rect 6687 4168 7328 4196
rect 6687 4165 6699 4168
rect 6641 4159 6699 4165
rect 1581 4131 1639 4137
rect 1581 4097 1593 4131
rect 1627 4128 1639 4131
rect 5718 4128 5724 4140
rect 1627 4100 5724 4128
rect 1627 4097 1639 4100
rect 1581 4091 1639 4097
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 934 4020 940 4072
rect 992 4060 998 4072
rect 1765 4063 1823 4069
rect 1765 4060 1777 4063
rect 992 4032 1777 4060
rect 992 4020 998 4032
rect 1765 4029 1777 4032
rect 1811 4029 1823 4063
rect 7300 4060 7328 4168
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 7576 4128 7604 4236
rect 8846 4224 8852 4236
rect 8904 4224 8910 4276
rect 11057 4267 11115 4273
rect 11057 4233 11069 4267
rect 11103 4264 11115 4267
rect 11146 4264 11152 4276
rect 11103 4236 11152 4264
rect 11103 4233 11115 4236
rect 11057 4227 11115 4233
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 11885 4267 11943 4273
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 14550 4264 14556 4276
rect 11931 4236 14556 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 14550 4224 14556 4236
rect 14608 4224 14614 4276
rect 15194 4224 15200 4276
rect 15252 4264 15258 4276
rect 21174 4264 21180 4276
rect 15252 4236 21180 4264
rect 15252 4224 15258 4236
rect 21174 4224 21180 4236
rect 21232 4224 21238 4276
rect 24670 4224 24676 4276
rect 24728 4264 24734 4276
rect 24765 4267 24823 4273
rect 24765 4264 24777 4267
rect 24728 4236 24777 4264
rect 24728 4224 24734 4236
rect 24765 4233 24777 4236
rect 24811 4233 24823 4267
rect 28350 4264 28356 4276
rect 24765 4227 24823 4233
rect 26344 4236 28356 4264
rect 9306 4196 9312 4208
rect 8404 4168 9312 4196
rect 8404 4140 8432 4168
rect 9306 4156 9312 4168
rect 9364 4196 9370 4208
rect 9953 4199 10011 4205
rect 9953 4196 9965 4199
rect 9364 4168 9965 4196
rect 9364 4156 9370 4168
rect 9953 4165 9965 4168
rect 9999 4165 10011 4199
rect 9953 4159 10011 4165
rect 10965 4199 11023 4205
rect 10965 4165 10977 4199
rect 11011 4196 11023 4199
rect 11698 4196 11704 4208
rect 11011 4168 11704 4196
rect 11011 4165 11023 4168
rect 10965 4159 11023 4165
rect 11698 4156 11704 4168
rect 11756 4156 11762 4208
rect 11793 4199 11851 4205
rect 11793 4165 11805 4199
rect 11839 4196 11851 4199
rect 12342 4196 12348 4208
rect 11839 4168 12348 4196
rect 11839 4165 11851 4168
rect 11793 4159 11851 4165
rect 12342 4156 12348 4168
rect 12400 4156 12406 4208
rect 12437 4199 12495 4205
rect 12437 4165 12449 4199
rect 12483 4196 12495 4199
rect 13354 4196 13360 4208
rect 12483 4168 13360 4196
rect 12483 4165 12495 4168
rect 12437 4159 12495 4165
rect 13354 4156 13360 4168
rect 13412 4196 13418 4208
rect 14277 4199 14335 4205
rect 14277 4196 14289 4199
rect 13412 4168 14289 4196
rect 13412 4156 13418 4168
rect 14277 4165 14289 4168
rect 14323 4165 14335 4199
rect 19886 4196 19892 4208
rect 14277 4159 14335 4165
rect 18064 4168 19892 4196
rect 7423 4100 7604 4128
rect 8021 4131 8079 4137
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8202 4128 8208 4140
rect 8067 4100 8208 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 8202 4088 8208 4100
rect 8260 4128 8266 4140
rect 8386 4128 8392 4140
rect 8260 4100 8392 4128
rect 8260 4088 8266 4100
rect 8386 4088 8392 4100
rect 8444 4088 8450 4140
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4128 9275 4131
rect 9263 4100 11192 4128
rect 9263 4097 9275 4100
rect 9217 4091 9275 4097
rect 8110 4060 8116 4072
rect 7300 4032 8116 4060
rect 1765 4023 1823 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 8938 4020 8944 4072
rect 8996 4020 9002 4072
rect 9122 4020 9128 4072
rect 9180 4020 9186 4072
rect 9306 4020 9312 4072
rect 9364 4020 9370 4072
rect 9401 4063 9459 4069
rect 9401 4029 9413 4063
rect 9447 4060 9459 4063
rect 9490 4060 9496 4072
rect 9447 4032 9496 4060
rect 9447 4029 9459 4032
rect 9401 4023 9459 4029
rect 9490 4020 9496 4032
rect 9548 4020 9554 4072
rect 10410 4020 10416 4072
rect 10468 4020 10474 4072
rect 5994 3952 6000 4004
rect 6052 3952 6058 4004
rect 6825 3995 6883 4001
rect 6825 3961 6837 3995
rect 6871 3992 6883 3995
rect 6871 3964 8340 3992
rect 6871 3961 6883 3964
rect 6825 3955 6883 3961
rect 7466 3884 7472 3936
rect 7524 3884 7530 3936
rect 8312 3924 8340 3964
rect 8386 3952 8392 4004
rect 8444 3952 8450 4004
rect 8481 3995 8539 4001
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 9766 3992 9772 4004
rect 8527 3964 9772 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 9766 3952 9772 3964
rect 9824 3952 9830 4004
rect 10229 3995 10287 4001
rect 10229 3961 10241 3995
rect 10275 3961 10287 3995
rect 10229 3955 10287 3961
rect 8662 3924 8668 3936
rect 8312 3896 8668 3924
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 10244 3924 10272 3955
rect 9456 3896 10272 3924
rect 11164 3924 11192 4100
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 17037 4131 17095 4137
rect 11296 4100 13676 4128
rect 11296 4088 11302 4100
rect 12894 4020 12900 4072
rect 12952 4020 12958 4072
rect 12710 3952 12716 4004
rect 12768 3952 12774 4004
rect 13648 4001 13676 4100
rect 13832 4100 16988 4128
rect 13832 4069 13860 4100
rect 13817 4063 13875 4069
rect 13817 4029 13829 4063
rect 13863 4029 13875 4063
rect 13817 4023 13875 4029
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4060 14795 4063
rect 14918 4060 14924 4072
rect 14783 4032 14924 4060
rect 14783 4029 14795 4032
rect 14737 4023 14795 4029
rect 14918 4020 14924 4032
rect 14976 4020 14982 4072
rect 15473 4063 15531 4069
rect 15473 4029 15485 4063
rect 15519 4060 15531 4063
rect 15838 4060 15844 4072
rect 15519 4032 15844 4060
rect 15519 4029 15531 4032
rect 15473 4023 15531 4029
rect 15838 4020 15844 4032
rect 15896 4060 15902 4072
rect 16114 4060 16120 4072
rect 15896 4032 16120 4060
rect 15896 4020 15902 4032
rect 16114 4020 16120 4032
rect 16172 4020 16178 4072
rect 16960 4060 16988 4100
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17126 4128 17132 4140
rect 17083 4100 17132 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 17957 4131 18015 4137
rect 17957 4097 17969 4131
rect 18003 4128 18015 4131
rect 18064 4128 18092 4168
rect 19886 4156 19892 4168
rect 19944 4156 19950 4208
rect 20064 4199 20122 4205
rect 20064 4165 20076 4199
rect 20110 4196 20122 4199
rect 20622 4196 20628 4208
rect 20110 4168 20628 4196
rect 20110 4165 20122 4168
rect 20064 4159 20122 4165
rect 20622 4156 20628 4168
rect 20680 4156 20686 4208
rect 20714 4156 20720 4208
rect 20772 4196 20778 4208
rect 26344 4196 26372 4236
rect 28350 4224 28356 4236
rect 28408 4224 28414 4276
rect 29546 4224 29552 4276
rect 29604 4264 29610 4276
rect 32677 4267 32735 4273
rect 29604 4236 31754 4264
rect 29604 4224 29610 4236
rect 20772 4168 26372 4196
rect 26421 4199 26479 4205
rect 20772 4156 20778 4168
rect 26421 4165 26433 4199
rect 26467 4196 26479 4199
rect 27154 4196 27160 4208
rect 26467 4168 27160 4196
rect 26467 4165 26479 4168
rect 26421 4159 26479 4165
rect 27154 4156 27160 4168
rect 27212 4156 27218 4208
rect 27430 4156 27436 4208
rect 27488 4196 27494 4208
rect 27488 4168 29224 4196
rect 27488 4156 27494 4168
rect 18003 4100 18092 4128
rect 18003 4097 18015 4100
rect 17957 4091 18015 4097
rect 18138 4088 18144 4140
rect 18196 4128 18202 4140
rect 18877 4131 18935 4137
rect 18877 4128 18889 4131
rect 18196 4100 18889 4128
rect 18196 4088 18202 4100
rect 18877 4097 18889 4100
rect 18923 4097 18935 4131
rect 18877 4091 18935 4097
rect 18966 4088 18972 4140
rect 19024 4128 19030 4140
rect 19024 4100 19380 4128
rect 19024 4088 19030 4100
rect 16960 4032 17264 4060
rect 13633 3995 13691 4001
rect 13633 3961 13645 3995
rect 13679 3961 13691 3995
rect 13633 3955 13691 3961
rect 13722 3952 13728 4004
rect 13780 3992 13786 4004
rect 14553 3995 14611 4001
rect 14553 3992 14565 3995
rect 13780 3964 14565 3992
rect 13780 3952 13786 3964
rect 14553 3961 14565 3964
rect 14599 3961 14611 3995
rect 14553 3955 14611 3961
rect 14826 3952 14832 4004
rect 14884 3992 14890 4004
rect 15749 3995 15807 4001
rect 15749 3992 15761 3995
rect 14884 3964 15761 3992
rect 14884 3952 14890 3964
rect 15749 3961 15761 3964
rect 15795 3961 15807 3995
rect 17236 3992 17264 4032
rect 17310 4020 17316 4072
rect 17368 4020 17374 4072
rect 18233 4063 18291 4069
rect 18233 4029 18245 4063
rect 18279 4060 18291 4063
rect 19153 4063 19211 4069
rect 18279 4032 19104 4060
rect 18279 4029 18291 4032
rect 18233 4023 18291 4029
rect 17954 3992 17960 4004
rect 15749 3955 15807 3961
rect 15856 3964 16896 3992
rect 17236 3964 17960 3992
rect 15856 3924 15884 3964
rect 11164 3896 15884 3924
rect 9456 3884 9462 3896
rect 15930 3884 15936 3936
rect 15988 3884 15994 3936
rect 16868 3924 16896 3964
rect 17954 3952 17960 3964
rect 18012 3952 18018 4004
rect 18966 3924 18972 3936
rect 16868 3896 18972 3924
rect 18966 3884 18972 3896
rect 19024 3884 19030 3936
rect 19076 3924 19104 4032
rect 19153 4029 19165 4063
rect 19199 4060 19211 4063
rect 19242 4060 19248 4072
rect 19199 4032 19248 4060
rect 19199 4029 19211 4032
rect 19153 4023 19211 4029
rect 19242 4020 19248 4032
rect 19300 4020 19306 4072
rect 19352 4060 19380 4100
rect 19702 4088 19708 4140
rect 19760 4128 19766 4140
rect 19797 4131 19855 4137
rect 19797 4128 19809 4131
rect 19760 4100 19809 4128
rect 19760 4088 19766 4100
rect 19797 4097 19809 4100
rect 19843 4097 19855 4131
rect 20438 4128 20444 4140
rect 19797 4091 19855 4097
rect 19904 4100 20444 4128
rect 19904 4060 19932 4100
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 22465 4131 22523 4137
rect 22465 4097 22477 4131
rect 22511 4128 22523 4131
rect 22646 4128 22652 4140
rect 22511 4100 22652 4128
rect 22511 4097 22523 4100
rect 22465 4091 22523 4097
rect 22646 4088 22652 4100
rect 22704 4088 22710 4140
rect 23290 4088 23296 4140
rect 23348 4128 23354 4140
rect 23385 4131 23443 4137
rect 23385 4128 23397 4131
rect 23348 4100 23397 4128
rect 23348 4088 23354 4100
rect 23385 4097 23397 4100
rect 23431 4097 23443 4131
rect 23385 4091 23443 4097
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 23641 4131 23699 4137
rect 23641 4128 23653 4131
rect 23532 4100 23653 4128
rect 23532 4088 23538 4100
rect 23641 4097 23653 4100
rect 23687 4097 23699 4131
rect 23641 4091 23699 4097
rect 25222 4088 25228 4140
rect 25280 4088 25286 4140
rect 27338 4128 27344 4140
rect 25516 4100 27344 4128
rect 19352 4032 19932 4060
rect 22741 4063 22799 4069
rect 22741 4029 22753 4063
rect 22787 4060 22799 4063
rect 23106 4060 23112 4072
rect 22787 4032 23112 4060
rect 22787 4029 22799 4032
rect 22741 4023 22799 4029
rect 23106 4020 23112 4032
rect 23164 4020 23170 4072
rect 24670 4020 24676 4072
rect 24728 4060 24734 4072
rect 25409 4063 25467 4069
rect 25409 4060 25421 4063
rect 24728 4032 25421 4060
rect 24728 4020 24734 4032
rect 25409 4029 25421 4032
rect 25455 4029 25467 4063
rect 25409 4023 25467 4029
rect 20070 3924 20076 3936
rect 19076 3896 20076 3924
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 25516 3924 25544 4100
rect 27338 4088 27344 4100
rect 27396 4088 27402 4140
rect 27522 4137 27528 4140
rect 27516 4128 27528 4137
rect 27483 4100 27528 4128
rect 27516 4091 27528 4100
rect 27522 4088 27528 4091
rect 27580 4088 27586 4140
rect 27890 4088 27896 4140
rect 27948 4128 27954 4140
rect 29089 4131 29147 4137
rect 29089 4128 29101 4131
rect 27948 4100 29101 4128
rect 27948 4088 27954 4100
rect 29089 4097 29101 4100
rect 29135 4097 29147 4131
rect 29196 4128 29224 4168
rect 30742 4156 30748 4208
rect 30800 4196 30806 4208
rect 31110 4196 31116 4208
rect 30800 4168 31116 4196
rect 30800 4156 30806 4168
rect 31110 4156 31116 4168
rect 31168 4156 31174 4208
rect 31573 4199 31631 4205
rect 31573 4165 31585 4199
rect 31619 4196 31631 4199
rect 31726 4196 31754 4236
rect 32677 4233 32689 4267
rect 32723 4264 32735 4267
rect 33318 4264 33324 4276
rect 32723 4236 33324 4264
rect 32723 4233 32735 4236
rect 32677 4227 32735 4233
rect 33318 4224 33324 4236
rect 33376 4224 33382 4276
rect 34238 4224 34244 4276
rect 34296 4264 34302 4276
rect 37366 4264 37372 4276
rect 34296 4236 37372 4264
rect 34296 4224 34302 4236
rect 37366 4224 37372 4236
rect 37424 4224 37430 4276
rect 37461 4267 37519 4273
rect 37461 4233 37473 4267
rect 37507 4264 37519 4267
rect 37826 4264 37832 4276
rect 37507 4236 37832 4264
rect 37507 4233 37519 4236
rect 37461 4227 37519 4233
rect 37826 4224 37832 4236
rect 37884 4224 37890 4276
rect 37921 4267 37979 4273
rect 37921 4233 37933 4267
rect 37967 4233 37979 4267
rect 37921 4227 37979 4233
rect 31619 4168 31984 4196
rect 31619 4165 31631 4168
rect 31573 4159 31631 4165
rect 29733 4131 29791 4137
rect 29733 4128 29745 4131
rect 29196 4100 29745 4128
rect 29089 4091 29147 4097
rect 29733 4097 29745 4100
rect 29779 4097 29791 4131
rect 31956 4128 31984 4168
rect 34606 4156 34612 4208
rect 34664 4156 34670 4208
rect 37734 4156 37740 4208
rect 37792 4196 37798 4208
rect 37936 4196 37964 4227
rect 38102 4224 38108 4276
rect 38160 4264 38166 4276
rect 38160 4236 41460 4264
rect 38160 4224 38166 4236
rect 37792 4168 37964 4196
rect 37792 4156 37798 4168
rect 38194 4156 38200 4208
rect 38252 4196 38258 4208
rect 41432 4205 41460 4236
rect 42058 4224 42064 4276
rect 42116 4264 42122 4276
rect 43346 4264 43352 4276
rect 42116 4236 43352 4264
rect 42116 4224 42122 4236
rect 43346 4224 43352 4236
rect 43404 4224 43410 4276
rect 53098 4224 53104 4276
rect 53156 4224 53162 4276
rect 39945 4199 40003 4205
rect 39945 4196 39957 4199
rect 38252 4168 39957 4196
rect 38252 4156 38258 4168
rect 39945 4165 39957 4168
rect 39991 4165 40003 4199
rect 40681 4199 40739 4205
rect 40681 4196 40693 4199
rect 39945 4159 40003 4165
rect 40052 4168 40693 4196
rect 33505 4131 33563 4137
rect 33505 4128 33517 4131
rect 31956 4100 33517 4128
rect 29733 4091 29791 4097
rect 33505 4097 33517 4100
rect 33551 4097 33563 4131
rect 33505 4091 33563 4097
rect 34425 4131 34483 4137
rect 34425 4097 34437 4131
rect 34471 4128 34483 4131
rect 34624 4128 34652 4156
rect 34471 4100 34652 4128
rect 34471 4097 34483 4100
rect 34425 4091 34483 4097
rect 35342 4088 35348 4140
rect 35400 4088 35406 4140
rect 35894 4088 35900 4140
rect 35952 4128 35958 4140
rect 36265 4131 36323 4137
rect 36265 4128 36277 4131
rect 35952 4100 36277 4128
rect 35952 4088 35958 4100
rect 36265 4097 36277 4100
rect 36311 4097 36323 4131
rect 36265 4091 36323 4097
rect 37826 4088 37832 4140
rect 37884 4088 37890 4140
rect 38749 4131 38807 4137
rect 38749 4097 38761 4131
rect 38795 4128 38807 4131
rect 39390 4128 39396 4140
rect 38795 4100 39396 4128
rect 38795 4097 38807 4100
rect 38749 4091 38807 4097
rect 39390 4088 39396 4100
rect 39448 4088 39454 4140
rect 40052 4128 40080 4168
rect 40681 4165 40693 4168
rect 40727 4165 40739 4199
rect 40681 4159 40739 4165
rect 41417 4199 41475 4205
rect 41417 4165 41429 4199
rect 41463 4165 41475 4199
rect 44361 4199 44419 4205
rect 44361 4196 44373 4199
rect 41417 4159 41475 4165
rect 42076 4168 44373 4196
rect 42076 4140 42104 4168
rect 44361 4165 44373 4168
rect 44407 4165 44419 4199
rect 44361 4159 44419 4165
rect 44818 4156 44824 4208
rect 44876 4196 44882 4208
rect 46569 4199 46627 4205
rect 46569 4196 46581 4199
rect 44876 4168 46581 4196
rect 44876 4156 44882 4168
rect 46569 4165 46581 4168
rect 46615 4165 46627 4199
rect 46569 4159 46627 4165
rect 51994 4156 52000 4208
rect 52052 4196 52058 4208
rect 52181 4199 52239 4205
rect 52181 4196 52193 4199
rect 52052 4168 52193 4196
rect 52052 4156 52058 4168
rect 52181 4165 52193 4168
rect 52227 4165 52239 4199
rect 52181 4159 52239 4165
rect 52822 4156 52828 4208
rect 52880 4196 52886 4208
rect 53009 4199 53067 4205
rect 53009 4196 53021 4199
rect 52880 4168 53021 4196
rect 52880 4156 52886 4168
rect 53009 4165 53021 4168
rect 53055 4165 53067 4199
rect 53009 4159 53067 4165
rect 53374 4156 53380 4208
rect 53432 4196 53438 4208
rect 53745 4199 53803 4205
rect 53745 4196 53757 4199
rect 53432 4168 53757 4196
rect 53432 4156 53438 4168
rect 53745 4165 53757 4168
rect 53791 4165 53803 4199
rect 53745 4159 53803 4165
rect 58161 4199 58219 4205
rect 58161 4165 58173 4199
rect 58207 4196 58219 4199
rect 58986 4196 58992 4208
rect 58207 4168 58992 4196
rect 58207 4165 58219 4168
rect 58161 4159 58219 4165
rect 58986 4156 58992 4168
rect 59044 4156 59050 4208
rect 39960 4100 40080 4128
rect 27249 4063 27307 4069
rect 27249 4029 27261 4063
rect 27295 4029 27307 4063
rect 27249 4023 27307 4029
rect 20772 3896 25544 3924
rect 27264 3924 27292 4023
rect 29638 4020 29644 4072
rect 29696 4060 29702 4072
rect 29917 4063 29975 4069
rect 29917 4060 29929 4063
rect 29696 4032 29929 4060
rect 29696 4020 29702 4032
rect 29917 4029 29929 4032
rect 29963 4029 29975 4063
rect 29917 4023 29975 4029
rect 32582 4020 32588 4072
rect 32640 4060 32646 4072
rect 32769 4063 32827 4069
rect 32769 4060 32781 4063
rect 32640 4032 32781 4060
rect 32640 4020 32646 4032
rect 32769 4029 32781 4032
rect 32815 4029 32827 4063
rect 32769 4023 32827 4029
rect 32858 4020 32864 4072
rect 32916 4020 32922 4072
rect 33134 4020 33140 4072
rect 33192 4060 33198 4072
rect 33689 4063 33747 4069
rect 33689 4060 33701 4063
rect 33192 4032 33701 4060
rect 33192 4020 33198 4032
rect 33689 4029 33701 4032
rect 33735 4029 33747 4063
rect 33689 4023 33747 4029
rect 34606 4020 34612 4072
rect 34664 4020 34670 4072
rect 34698 4020 34704 4072
rect 34756 4060 34762 4072
rect 35529 4063 35587 4069
rect 35529 4060 35541 4063
rect 34756 4032 35541 4060
rect 34756 4020 34762 4032
rect 35529 4029 35541 4032
rect 35575 4029 35587 4063
rect 35529 4023 35587 4029
rect 35618 4020 35624 4072
rect 35676 4060 35682 4072
rect 36449 4063 36507 4069
rect 36449 4060 36461 4063
rect 35676 4032 36461 4060
rect 35676 4020 35682 4032
rect 36449 4029 36461 4032
rect 36495 4029 36507 4063
rect 36449 4023 36507 4029
rect 38105 4063 38163 4069
rect 38105 4029 38117 4063
rect 38151 4060 38163 4063
rect 39301 4063 39359 4069
rect 39301 4060 39313 4063
rect 38151 4032 39313 4060
rect 38151 4029 38163 4032
rect 38105 4023 38163 4029
rect 39301 4029 39313 4032
rect 39347 4060 39359 4063
rect 39850 4060 39856 4072
rect 39347 4032 39856 4060
rect 39347 4029 39359 4032
rect 39301 4023 39359 4029
rect 31757 3995 31815 4001
rect 31757 3961 31769 3995
rect 31803 3992 31815 3995
rect 32122 3992 32128 4004
rect 31803 3964 32128 3992
rect 31803 3961 31815 3964
rect 31757 3955 31815 3961
rect 32122 3952 32128 3964
rect 32180 3952 32186 4004
rect 32876 3992 32904 4020
rect 32876 3964 37969 3992
rect 28442 3924 28448 3936
rect 27264 3896 28448 3924
rect 20772 3884 20778 3896
rect 28442 3884 28448 3896
rect 28500 3884 28506 3936
rect 28626 3884 28632 3936
rect 28684 3884 28690 3936
rect 30834 3884 30840 3936
rect 30892 3884 30898 3936
rect 31570 3884 31576 3936
rect 31628 3924 31634 3936
rect 32309 3927 32367 3933
rect 32309 3924 32321 3927
rect 31628 3896 32321 3924
rect 31628 3884 31634 3896
rect 32309 3893 32321 3896
rect 32355 3893 32367 3927
rect 37941 3924 37969 3964
rect 38120 3924 38148 4023
rect 39850 4020 39856 4032
rect 39908 4020 39914 4072
rect 38194 3952 38200 4004
rect 38252 3992 38258 4004
rect 39960 3992 39988 4100
rect 40126 4088 40132 4140
rect 40184 4128 40190 4140
rect 40865 4131 40923 4137
rect 40865 4128 40877 4131
rect 40184 4100 40877 4128
rect 40184 4088 40190 4100
rect 40865 4097 40877 4100
rect 40911 4097 40923 4131
rect 40865 4091 40923 4097
rect 41598 4088 41604 4140
rect 41656 4088 41662 4140
rect 42058 4088 42064 4140
rect 42116 4088 42122 4140
rect 42978 4088 42984 4140
rect 43036 4128 43042 4140
rect 43257 4131 43315 4137
rect 43257 4128 43269 4131
rect 43036 4100 43269 4128
rect 43036 4088 43042 4100
rect 43257 4097 43269 4100
rect 43303 4097 43315 4131
rect 43257 4091 43315 4097
rect 43625 4131 43683 4137
rect 43625 4097 43637 4131
rect 43671 4128 43683 4131
rect 44266 4128 44272 4140
rect 43671 4100 44272 4128
rect 43671 4097 43683 4100
rect 43625 4091 43683 4097
rect 44266 4088 44272 4100
rect 44324 4088 44330 4140
rect 44910 4088 44916 4140
rect 44968 4128 44974 4140
rect 45097 4131 45155 4137
rect 45097 4128 45109 4131
rect 44968 4100 45109 4128
rect 44968 4088 44974 4100
rect 45097 4097 45109 4100
rect 45143 4097 45155 4131
rect 45833 4131 45891 4137
rect 45833 4128 45845 4131
rect 45097 4091 45155 4097
rect 45204 4100 45845 4128
rect 42610 4020 42616 4072
rect 42668 4020 42674 4072
rect 43070 4020 43076 4072
rect 43128 4020 43134 4072
rect 43438 4020 43444 4072
rect 43496 4060 43502 4072
rect 43533 4063 43591 4069
rect 43533 4060 43545 4063
rect 43496 4032 43545 4060
rect 43496 4020 43502 4032
rect 43533 4029 43545 4032
rect 43579 4029 43591 4063
rect 43533 4023 43591 4029
rect 43990 4020 43996 4072
rect 44048 4060 44054 4072
rect 45204 4060 45232 4100
rect 45833 4097 45845 4100
rect 45879 4097 45891 4131
rect 45833 4091 45891 4097
rect 45922 4088 45928 4140
rect 45980 4128 45986 4140
rect 46017 4131 46075 4137
rect 46017 4128 46029 4131
rect 45980 4100 46029 4128
rect 45980 4088 45986 4100
rect 46017 4097 46029 4100
rect 46063 4097 46075 4131
rect 46017 4091 46075 4097
rect 46750 4088 46756 4140
rect 46808 4088 46814 4140
rect 48130 4088 48136 4140
rect 48188 4128 48194 4140
rect 48225 4131 48283 4137
rect 48225 4128 48237 4131
rect 48188 4100 48237 4128
rect 48188 4088 48194 4100
rect 48225 4097 48237 4100
rect 48271 4097 48283 4131
rect 48225 4091 48283 4097
rect 52362 4088 52368 4140
rect 52420 4128 52426 4140
rect 53929 4131 53987 4137
rect 53929 4128 53941 4131
rect 52420 4100 53941 4128
rect 52420 4088 52426 4100
rect 53929 4097 53941 4100
rect 53975 4097 53987 4131
rect 53929 4091 53987 4097
rect 54478 4088 54484 4140
rect 54536 4128 54542 4140
rect 54573 4131 54631 4137
rect 54573 4128 54585 4131
rect 54536 4100 54585 4128
rect 54536 4088 54542 4100
rect 54573 4097 54585 4100
rect 54619 4097 54631 4131
rect 54573 4091 54631 4097
rect 44048 4032 45232 4060
rect 44048 4020 44054 4032
rect 46382 4020 46388 4072
rect 46440 4060 46446 4072
rect 46440 4032 51074 4060
rect 46440 4020 46446 4032
rect 38252 3964 39988 3992
rect 40129 3995 40187 4001
rect 38252 3952 38258 3964
rect 40129 3961 40141 3995
rect 40175 3992 40187 3995
rect 40402 3992 40408 4004
rect 40175 3964 40408 3992
rect 40175 3961 40187 3964
rect 40129 3955 40187 3961
rect 40402 3952 40408 3964
rect 40460 3952 40466 4004
rect 41690 3952 41696 4004
rect 41748 3992 41754 4004
rect 47946 3992 47952 4004
rect 41748 3964 47952 3992
rect 41748 3952 41754 3964
rect 47946 3952 47952 3964
rect 48004 3952 48010 4004
rect 48406 3952 48412 4004
rect 48464 3952 48470 4004
rect 51046 3992 51074 4032
rect 52270 4020 52276 4072
rect 52328 4060 52334 4072
rect 58345 4063 58403 4069
rect 58345 4060 58357 4063
rect 52328 4032 58357 4060
rect 52328 4020 52334 4032
rect 58345 4029 58357 4032
rect 58391 4029 58403 4063
rect 58345 4023 58403 4029
rect 51046 3964 53604 3992
rect 37941 3896 38148 3924
rect 32309 3887 32367 3893
rect 43622 3884 43628 3936
rect 43680 3924 43686 3936
rect 44453 3927 44511 3933
rect 44453 3924 44465 3927
rect 43680 3896 44465 3924
rect 43680 3884 43686 3896
rect 44453 3893 44465 3896
rect 44499 3893 44511 3927
rect 44453 3887 44511 3893
rect 45186 3884 45192 3936
rect 45244 3884 45250 3936
rect 52270 3884 52276 3936
rect 52328 3884 52334 3936
rect 53576 3924 53604 3964
rect 53650 3952 53656 4004
rect 53708 3992 53714 4004
rect 54757 3995 54815 4001
rect 54757 3992 54769 3995
rect 53708 3964 54769 3992
rect 53708 3952 53714 3964
rect 54757 3961 54769 3964
rect 54803 3961 54815 3995
rect 54757 3955 54815 3961
rect 57422 3924 57428 3936
rect 53576 3896 57428 3924
rect 57422 3884 57428 3896
rect 57480 3884 57486 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 7524 3692 10732 3720
rect 7524 3680 7530 3692
rect 5258 3612 5264 3664
rect 5316 3612 5322 3664
rect 5997 3655 6055 3661
rect 5997 3621 6009 3655
rect 6043 3652 6055 3655
rect 6178 3652 6184 3664
rect 6043 3624 6184 3652
rect 6043 3621 6055 3624
rect 5997 3615 6055 3621
rect 6178 3612 6184 3624
rect 6236 3612 6242 3664
rect 7558 3612 7564 3664
rect 7616 3612 7622 3664
rect 8481 3655 8539 3661
rect 8481 3621 8493 3655
rect 8527 3621 8539 3655
rect 8481 3615 8539 3621
rect 6733 3587 6791 3593
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 8496 3584 8524 3615
rect 8570 3612 8576 3664
rect 8628 3612 8634 3664
rect 10704 3661 10732 3692
rect 10870 3680 10876 3732
rect 10928 3680 10934 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 13722 3720 13728 3732
rect 11112 3692 13728 3720
rect 11112 3680 11118 3692
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 16209 3723 16267 3729
rect 14108 3692 16160 3720
rect 10689 3655 10747 3661
rect 10689 3621 10701 3655
rect 10735 3621 10747 3655
rect 10689 3615 10747 3621
rect 12066 3612 12072 3664
rect 12124 3612 12130 3664
rect 12526 3612 12532 3664
rect 12584 3652 12590 3664
rect 13541 3655 13599 3661
rect 13541 3652 13553 3655
rect 12584 3624 13553 3652
rect 12584 3612 12590 3624
rect 13541 3621 13553 3624
rect 13587 3621 13599 3655
rect 14108 3652 14136 3692
rect 13541 3615 13599 3621
rect 13648 3624 14136 3652
rect 6779 3556 8524 3584
rect 9401 3587 9459 3593
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 9401 3553 9413 3587
rect 9447 3553 9459 3587
rect 9401 3547 9459 3553
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 13648 3584 13676 3624
rect 14182 3612 14188 3664
rect 14240 3652 14246 3664
rect 14553 3655 14611 3661
rect 14553 3652 14565 3655
rect 14240 3624 14565 3652
rect 14240 3612 14246 3624
rect 14553 3621 14565 3624
rect 14599 3621 14611 3655
rect 14553 3615 14611 3621
rect 14642 3612 14648 3664
rect 14700 3652 14706 3664
rect 16025 3655 16083 3661
rect 16025 3652 16037 3655
rect 14700 3624 16037 3652
rect 14700 3612 14706 3624
rect 16025 3621 16037 3624
rect 16071 3621 16083 3655
rect 16025 3615 16083 3621
rect 9723 3556 13676 3584
rect 13725 3587 13783 3593
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 13725 3553 13737 3587
rect 13771 3584 13783 3587
rect 14090 3584 14096 3596
rect 13771 3556 14096 3584
rect 13771 3553 13783 3556
rect 13725 3547 13783 3553
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 9416 3516 9444 3547
rect 14090 3544 14096 3556
rect 14148 3544 14154 3596
rect 14737 3587 14795 3593
rect 14737 3553 14749 3587
rect 14783 3584 14795 3587
rect 15194 3584 15200 3596
rect 14783 3556 15200 3584
rect 14783 3553 14795 3556
rect 14737 3547 14795 3553
rect 15194 3544 15200 3556
rect 15252 3544 15258 3596
rect 15749 3587 15807 3593
rect 15749 3553 15761 3587
rect 15795 3584 15807 3587
rect 15838 3584 15844 3596
rect 15795 3556 15844 3584
rect 15795 3553 15807 3556
rect 15749 3547 15807 3553
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 16132 3584 16160 3692
rect 16209 3689 16221 3723
rect 16255 3720 16267 3723
rect 16255 3692 23704 3720
rect 16255 3689 16267 3692
rect 16209 3683 16267 3689
rect 21085 3655 21143 3661
rect 21085 3621 21097 3655
rect 21131 3621 21143 3655
rect 23676 3652 23704 3692
rect 23750 3680 23756 3732
rect 23808 3720 23814 3732
rect 24581 3723 24639 3729
rect 24581 3720 24593 3723
rect 23808 3692 24593 3720
rect 23808 3680 23814 3692
rect 24581 3689 24593 3692
rect 24627 3689 24639 3723
rect 24581 3683 24639 3689
rect 24946 3680 24952 3732
rect 25004 3720 25010 3732
rect 25314 3720 25320 3732
rect 25004 3692 25320 3720
rect 25004 3680 25010 3692
rect 25314 3680 25320 3692
rect 25372 3720 25378 3732
rect 27246 3720 27252 3732
rect 25372 3692 27252 3720
rect 25372 3680 25378 3692
rect 27246 3680 27252 3692
rect 27304 3680 27310 3732
rect 27798 3680 27804 3732
rect 27856 3680 27862 3732
rect 28442 3680 28448 3732
rect 28500 3720 28506 3732
rect 31294 3720 31300 3732
rect 28500 3692 31300 3720
rect 28500 3680 28506 3692
rect 31294 3680 31300 3692
rect 31352 3680 31358 3732
rect 33318 3680 33324 3732
rect 33376 3720 33382 3732
rect 33597 3723 33655 3729
rect 33597 3720 33609 3723
rect 33376 3692 33609 3720
rect 33376 3680 33382 3692
rect 33597 3689 33609 3692
rect 33643 3689 33655 3723
rect 33597 3683 33655 3689
rect 36541 3723 36599 3729
rect 36541 3689 36553 3723
rect 36587 3720 36599 3723
rect 36630 3720 36636 3732
rect 36587 3692 36636 3720
rect 36587 3689 36599 3692
rect 36541 3683 36599 3689
rect 36630 3680 36636 3692
rect 36688 3680 36694 3732
rect 37016 3692 38148 3720
rect 30466 3652 30472 3664
rect 23676 3624 30472 3652
rect 21085 3615 21143 3621
rect 18601 3587 18659 3593
rect 18601 3584 18613 3587
rect 16132 3556 18613 3584
rect 18601 3553 18613 3556
rect 18647 3553 18659 3587
rect 18601 3547 18659 3553
rect 18785 3587 18843 3593
rect 18785 3553 18797 3587
rect 18831 3584 18843 3587
rect 19058 3584 19064 3596
rect 18831 3556 19064 3584
rect 18831 3553 18843 3556
rect 18785 3547 18843 3553
rect 1627 3488 9444 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 9582 3476 9588 3528
rect 9640 3476 9646 3528
rect 9769 3519 9827 3525
rect 9769 3485 9781 3519
rect 9815 3485 9827 3519
rect 9769 3479 9827 3485
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 1857 3451 1915 3457
rect 1857 3448 1869 3451
rect 992 3420 1869 3448
rect 992 3408 998 3420
rect 1857 3417 1869 3420
rect 1903 3417 1915 3451
rect 1857 3411 1915 3417
rect 5074 3408 5080 3460
rect 5132 3408 5138 3460
rect 5813 3451 5871 3457
rect 5813 3417 5825 3451
rect 5859 3448 5871 3451
rect 6549 3451 6607 3457
rect 5859 3420 6500 3448
rect 5859 3417 5871 3420
rect 5813 3411 5871 3417
rect 6472 3380 6500 3420
rect 6549 3417 6561 3451
rect 6595 3448 6607 3451
rect 7098 3448 7104 3460
rect 6595 3420 7104 3448
rect 6595 3417 6607 3420
rect 6549 3411 6607 3417
rect 7098 3408 7104 3420
rect 7156 3408 7162 3460
rect 7193 3451 7251 3457
rect 7193 3417 7205 3451
rect 7239 3448 7251 3451
rect 8113 3451 8171 3457
rect 8113 3448 8125 3451
rect 7239 3420 8125 3448
rect 7239 3417 7251 3420
rect 7193 3411 7251 3417
rect 8113 3417 8125 3420
rect 8159 3448 8171 3451
rect 8202 3448 8208 3460
rect 8159 3420 8208 3448
rect 8159 3417 8171 3420
rect 8113 3411 8171 3417
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 9490 3448 9496 3460
rect 8496 3420 9496 3448
rect 7282 3380 7288 3392
rect 6472 3352 7288 3380
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7653 3383 7711 3389
rect 7653 3349 7665 3383
rect 7699 3380 7711 3383
rect 8496 3380 8524 3420
rect 9490 3408 9496 3420
rect 9548 3408 9554 3460
rect 9784 3448 9812 3479
rect 9858 3476 9864 3528
rect 9916 3476 9922 3528
rect 12805 3519 12863 3525
rect 12805 3485 12817 3519
rect 12851 3516 12863 3519
rect 14826 3516 14832 3528
rect 12851 3488 14832 3516
rect 12851 3485 12863 3488
rect 12805 3479 12863 3485
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 17221 3519 17279 3525
rect 17221 3516 17233 3519
rect 16816 3488 17233 3516
rect 16816 3476 16822 3488
rect 17221 3485 17233 3488
rect 17267 3485 17279 3519
rect 17221 3479 17279 3485
rect 18506 3476 18512 3528
rect 18564 3476 18570 3528
rect 18616 3516 18644 3547
rect 19058 3544 19064 3556
rect 19116 3544 19122 3596
rect 19426 3544 19432 3596
rect 19484 3584 19490 3596
rect 19702 3584 19708 3596
rect 19484 3556 19708 3584
rect 19484 3544 19490 3556
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 21100 3516 21128 3615
rect 30466 3612 30472 3624
rect 30524 3612 30530 3664
rect 37016 3652 37044 3692
rect 36280 3624 37044 3652
rect 25130 3544 25136 3596
rect 25188 3544 25194 3596
rect 25961 3587 26019 3593
rect 25961 3584 25973 3587
rect 25240 3556 25973 3584
rect 18616 3488 21128 3516
rect 21729 3519 21787 3525
rect 21729 3485 21741 3519
rect 21775 3516 21787 3519
rect 21910 3516 21916 3528
rect 21775 3488 21916 3516
rect 21775 3485 21787 3488
rect 21729 3479 21787 3485
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 22646 3476 22652 3528
rect 22704 3516 22710 3528
rect 23290 3516 23296 3528
rect 22704 3488 23296 3516
rect 22704 3476 22710 3488
rect 23290 3476 23296 3488
rect 23348 3476 23354 3528
rect 23842 3476 23848 3528
rect 23900 3516 23906 3528
rect 25240 3516 25268 3556
rect 25961 3553 25973 3556
rect 26007 3553 26019 3587
rect 27982 3584 27988 3596
rect 25961 3547 26019 3553
rect 26988 3556 27988 3584
rect 23900 3488 25268 3516
rect 23900 3476 23906 3488
rect 25774 3476 25780 3528
rect 25832 3476 25838 3528
rect 26988 3460 27016 3556
rect 27982 3544 27988 3556
rect 28040 3544 28046 3596
rect 28258 3544 28264 3596
rect 28316 3544 28322 3596
rect 28445 3587 28503 3593
rect 28445 3553 28457 3587
rect 28491 3584 28503 3587
rect 28810 3584 28816 3596
rect 28491 3556 28816 3584
rect 28491 3553 28503 3556
rect 28445 3547 28503 3553
rect 28810 3544 28816 3556
rect 28868 3544 28874 3596
rect 31294 3544 31300 3596
rect 31352 3584 31358 3596
rect 32217 3587 32275 3593
rect 32217 3584 32229 3587
rect 31352 3556 32229 3584
rect 31352 3544 31358 3556
rect 32217 3553 32229 3556
rect 32263 3553 32275 3587
rect 32217 3547 32275 3553
rect 33410 3544 33416 3596
rect 33468 3584 33474 3596
rect 34606 3584 34612 3596
rect 33468 3556 34612 3584
rect 33468 3544 33474 3556
rect 34606 3544 34612 3556
rect 34664 3544 34670 3596
rect 27111 3519 27169 3525
rect 27111 3485 27123 3519
rect 27157 3516 27169 3519
rect 27157 3488 27292 3516
rect 27157 3485 27169 3488
rect 27111 3479 27169 3485
rect 10413 3451 10471 3457
rect 10413 3448 10425 3451
rect 9784 3420 10425 3448
rect 7699 3352 8524 3380
rect 7699 3349 7711 3352
rect 7653 3343 7711 3349
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 9784 3380 9812 3420
rect 10413 3417 10425 3420
rect 10459 3417 10471 3451
rect 10413 3411 10471 3417
rect 11885 3451 11943 3457
rect 11885 3417 11897 3451
rect 11931 3448 11943 3451
rect 11931 3420 12434 3448
rect 11931 3417 11943 3420
rect 11885 3411 11943 3417
rect 9364 3352 9812 3380
rect 12406 3380 12434 3420
rect 12618 3408 12624 3460
rect 12676 3408 12682 3460
rect 13262 3408 13268 3460
rect 13320 3448 13326 3460
rect 14277 3451 14335 3457
rect 14277 3448 14289 3451
rect 13320 3420 14289 3448
rect 13320 3408 13326 3420
rect 14277 3417 14289 3420
rect 14323 3417 14335 3451
rect 14277 3411 14335 3417
rect 17494 3408 17500 3460
rect 17552 3408 17558 3460
rect 19950 3451 20008 3457
rect 19950 3448 19962 3451
rect 18156 3420 19962 3448
rect 13354 3380 13360 3392
rect 12406 3352 13360 3380
rect 9364 3340 9370 3352
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 18156 3389 18184 3420
rect 19950 3417 19962 3420
rect 19996 3417 20008 3451
rect 19950 3411 20008 3417
rect 20088 3420 21220 3448
rect 18141 3383 18199 3389
rect 18141 3349 18153 3383
rect 18187 3349 18199 3383
rect 18141 3343 18199 3349
rect 19334 3340 19340 3392
rect 19392 3380 19398 3392
rect 20088 3380 20116 3420
rect 19392 3352 20116 3380
rect 21192 3380 21220 3420
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 22916 3451 22974 3457
rect 22916 3417 22928 3451
rect 22962 3448 22974 3451
rect 23198 3448 23204 3460
rect 22962 3420 23204 3448
rect 22962 3417 22974 3420
rect 22916 3411 22974 3417
rect 23198 3408 23204 3420
rect 23256 3408 23262 3460
rect 24949 3451 25007 3457
rect 24949 3448 24961 3451
rect 23492 3420 24961 3448
rect 23492 3380 23520 3420
rect 24949 3417 24961 3420
rect 24995 3417 25007 3451
rect 24949 3411 25007 3417
rect 26786 3408 26792 3460
rect 26844 3408 26850 3460
rect 26970 3408 26976 3460
rect 27028 3408 27034 3460
rect 27264 3448 27292 3488
rect 27338 3476 27344 3528
rect 27396 3476 27402 3528
rect 28626 3516 28632 3528
rect 27908 3488 28632 3516
rect 27908 3448 27936 3488
rect 28626 3476 28632 3488
rect 28684 3476 28690 3528
rect 30282 3476 30288 3528
rect 30340 3476 30346 3528
rect 30926 3476 30932 3528
rect 30984 3516 30990 3528
rect 31389 3519 31447 3525
rect 31389 3516 31401 3519
rect 30984 3488 31401 3516
rect 30984 3476 30990 3488
rect 31389 3485 31401 3488
rect 31435 3485 31447 3519
rect 31389 3479 31447 3485
rect 31570 3476 31576 3528
rect 31628 3476 31634 3528
rect 31757 3519 31815 3525
rect 31757 3485 31769 3519
rect 31803 3516 31815 3519
rect 32493 3519 32551 3525
rect 32493 3516 32505 3519
rect 31803 3488 32505 3516
rect 31803 3485 31815 3488
rect 31757 3479 31815 3485
rect 32493 3485 32505 3488
rect 32539 3485 32551 3519
rect 32493 3479 32551 3485
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34848 3488 34897 3516
rect 34848 3476 34854 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 34885 3479 34943 3485
rect 35894 3476 35900 3528
rect 35952 3476 35958 3528
rect 36045 3519 36103 3525
rect 36045 3485 36057 3519
rect 36091 3516 36103 3519
rect 36280 3516 36308 3624
rect 36998 3544 37004 3596
rect 37056 3544 37062 3596
rect 37277 3587 37335 3593
rect 37277 3553 37289 3587
rect 37323 3584 37335 3587
rect 38010 3584 38016 3596
rect 37323 3556 38016 3584
rect 37323 3553 37335 3556
rect 37277 3547 37335 3553
rect 38010 3544 38016 3556
rect 38068 3544 38074 3596
rect 38120 3584 38148 3692
rect 38194 3680 38200 3732
rect 38252 3720 38258 3732
rect 40862 3720 40868 3732
rect 38252 3692 40868 3720
rect 38252 3680 38258 3692
rect 40862 3680 40868 3692
rect 40920 3680 40926 3732
rect 41046 3680 41052 3732
rect 41104 3720 41110 3732
rect 41690 3720 41696 3732
rect 41104 3692 41696 3720
rect 41104 3680 41110 3692
rect 41690 3680 41696 3692
rect 41748 3680 41754 3732
rect 42702 3720 42708 3732
rect 41984 3692 42708 3720
rect 38286 3612 38292 3664
rect 38344 3652 38350 3664
rect 38381 3655 38439 3661
rect 38381 3652 38393 3655
rect 38344 3624 38393 3652
rect 38344 3612 38350 3624
rect 38381 3621 38393 3624
rect 38427 3621 38439 3655
rect 38381 3615 38439 3621
rect 39022 3612 39028 3664
rect 39080 3652 39086 3664
rect 40218 3652 40224 3664
rect 39080 3624 40224 3652
rect 39080 3612 39086 3624
rect 40218 3612 40224 3624
rect 40276 3612 40282 3664
rect 40402 3612 40408 3664
rect 40460 3612 40466 3664
rect 41984 3652 42012 3692
rect 42702 3680 42708 3692
rect 42760 3680 42766 3732
rect 44266 3680 44272 3732
rect 44324 3720 44330 3732
rect 45373 3723 45431 3729
rect 45373 3720 45385 3723
rect 44324 3692 45385 3720
rect 44324 3680 44330 3692
rect 45373 3689 45385 3692
rect 45419 3689 45431 3723
rect 45373 3683 45431 3689
rect 45554 3680 45560 3732
rect 45612 3720 45618 3732
rect 46109 3723 46167 3729
rect 46109 3720 46121 3723
rect 45612 3692 46121 3720
rect 45612 3680 45618 3692
rect 46109 3689 46121 3692
rect 46155 3689 46167 3723
rect 46109 3683 46167 3689
rect 47026 3680 47032 3732
rect 47084 3680 47090 3732
rect 47946 3680 47952 3732
rect 48004 3680 48010 3732
rect 48590 3680 48596 3732
rect 48648 3720 48654 3732
rect 48685 3723 48743 3729
rect 48685 3720 48697 3723
rect 48648 3692 48697 3720
rect 48648 3680 48654 3692
rect 48685 3689 48697 3692
rect 48731 3689 48743 3723
rect 48685 3683 48743 3689
rect 49418 3680 49424 3732
rect 49476 3680 49482 3732
rect 50154 3680 50160 3732
rect 50212 3720 50218 3732
rect 50525 3723 50583 3729
rect 50525 3720 50537 3723
rect 50212 3692 50537 3720
rect 50212 3680 50218 3692
rect 50525 3689 50537 3692
rect 50571 3689 50583 3723
rect 50525 3683 50583 3689
rect 51350 3680 51356 3732
rect 51408 3720 51414 3732
rect 51997 3723 52055 3729
rect 51997 3720 52009 3723
rect 51408 3692 52009 3720
rect 51408 3680 51414 3692
rect 51997 3689 52009 3692
rect 52043 3689 52055 3723
rect 51997 3683 52055 3689
rect 54202 3680 54208 3732
rect 54260 3680 54266 3732
rect 40880 3624 42012 3652
rect 42061 3655 42119 3661
rect 40586 3584 40592 3596
rect 38120 3556 40592 3584
rect 40586 3544 40592 3556
rect 40644 3544 40650 3596
rect 40880 3593 40908 3624
rect 42061 3621 42073 3655
rect 42107 3652 42119 3655
rect 42150 3652 42156 3664
rect 42107 3624 42156 3652
rect 42107 3621 42119 3624
rect 42061 3615 42119 3621
rect 42150 3612 42156 3624
rect 42208 3612 42214 3664
rect 45002 3652 45008 3664
rect 43640 3624 45008 3652
rect 40865 3587 40923 3593
rect 40865 3553 40877 3587
rect 40911 3553 40923 3587
rect 40865 3547 40923 3553
rect 41322 3544 41328 3596
rect 41380 3584 41386 3596
rect 42889 3587 42947 3593
rect 42889 3584 42901 3587
rect 41380 3556 42901 3584
rect 41380 3544 41386 3556
rect 42889 3553 42901 3556
rect 42935 3553 42947 3587
rect 42889 3547 42947 3553
rect 36091 3488 36308 3516
rect 36403 3519 36461 3525
rect 36091 3485 36103 3488
rect 36045 3479 36103 3485
rect 36403 3485 36415 3519
rect 36449 3516 36461 3519
rect 36906 3516 36912 3528
rect 36449 3488 36912 3516
rect 36449 3485 36461 3488
rect 36403 3479 36461 3485
rect 36906 3476 36912 3488
rect 36964 3476 36970 3528
rect 38838 3516 38844 3528
rect 37108 3488 38844 3516
rect 27264 3420 27936 3448
rect 27982 3408 27988 3460
rect 28040 3448 28046 3460
rect 28997 3451 29055 3457
rect 28997 3448 29009 3451
rect 28040 3420 29009 3448
rect 28040 3408 28046 3420
rect 28997 3417 29009 3420
rect 29043 3417 29055 3451
rect 28997 3411 29055 3417
rect 30190 3408 30196 3460
rect 30248 3448 30254 3460
rect 30561 3451 30619 3457
rect 30561 3448 30573 3451
rect 30248 3420 30573 3448
rect 30248 3408 30254 3420
rect 30561 3417 30573 3420
rect 30607 3417 30619 3451
rect 30561 3411 30619 3417
rect 33226 3408 33232 3460
rect 33284 3448 33290 3460
rect 35161 3451 35219 3457
rect 35161 3448 35173 3451
rect 33284 3420 35173 3448
rect 33284 3408 33290 3420
rect 35161 3417 35173 3420
rect 35207 3417 35219 3451
rect 35161 3411 35219 3417
rect 36173 3451 36231 3457
rect 36173 3417 36185 3451
rect 36219 3417 36231 3451
rect 36173 3411 36231 3417
rect 36265 3451 36323 3457
rect 36265 3417 36277 3451
rect 36311 3448 36323 3451
rect 37108 3448 37136 3488
rect 38838 3476 38844 3488
rect 38896 3476 38902 3528
rect 40770 3516 40776 3528
rect 39040 3488 40776 3516
rect 39040 3448 39068 3488
rect 40770 3476 40776 3488
rect 40828 3476 40834 3528
rect 41138 3476 41144 3528
rect 41196 3476 41202 3528
rect 41230 3476 41236 3528
rect 41288 3516 41294 3528
rect 43349 3519 43407 3525
rect 43349 3516 43361 3519
rect 41288 3488 43361 3516
rect 41288 3476 41294 3488
rect 43349 3485 43361 3488
rect 43395 3516 43407 3519
rect 43438 3516 43444 3528
rect 43395 3488 43444 3516
rect 43395 3485 43407 3488
rect 43349 3479 43407 3485
rect 43438 3476 43444 3488
rect 43496 3476 43502 3528
rect 43640 3525 43668 3624
rect 45002 3612 45008 3624
rect 45060 3612 45066 3664
rect 45094 3612 45100 3664
rect 45152 3652 45158 3664
rect 46014 3652 46020 3664
rect 45152 3624 46020 3652
rect 45152 3612 45158 3624
rect 46014 3612 46020 3624
rect 46072 3612 46078 3664
rect 48314 3612 48320 3664
rect 48372 3652 48378 3664
rect 52825 3655 52883 3661
rect 52825 3652 52837 3655
rect 48372 3624 52837 3652
rect 48372 3612 48378 3624
rect 52825 3621 52837 3624
rect 52871 3621 52883 3655
rect 52825 3615 52883 3621
rect 53834 3612 53840 3664
rect 53892 3652 53898 3664
rect 55677 3655 55735 3661
rect 55677 3652 55689 3655
rect 53892 3624 55689 3652
rect 53892 3612 53898 3624
rect 55677 3621 55689 3624
rect 55723 3621 55735 3655
rect 55677 3615 55735 3621
rect 52270 3584 52276 3596
rect 44284 3556 52276 3584
rect 43625 3519 43683 3525
rect 43625 3485 43637 3519
rect 43671 3485 43683 3519
rect 43625 3479 43683 3485
rect 43714 3476 43720 3528
rect 43772 3476 43778 3528
rect 44284 3525 44312 3556
rect 52270 3544 52276 3556
rect 52328 3544 52334 3596
rect 56870 3544 56876 3596
rect 56928 3544 56934 3596
rect 43993 3519 44051 3525
rect 43993 3485 44005 3519
rect 44039 3485 44051 3519
rect 43993 3479 44051 3485
rect 44269 3519 44327 3525
rect 44269 3485 44281 3519
rect 44315 3485 44327 3519
rect 44269 3479 44327 3485
rect 46017 3519 46075 3525
rect 46017 3485 46029 3519
rect 46063 3516 46075 3519
rect 46106 3516 46112 3528
rect 46063 3488 46112 3516
rect 46063 3485 46075 3488
rect 46017 3479 46075 3485
rect 36311 3420 37136 3448
rect 37936 3420 39068 3448
rect 36311 3417 36323 3420
rect 36265 3411 36323 3417
rect 21192 3352 23520 3380
rect 19392 3340 19398 3352
rect 24026 3340 24032 3392
rect 24084 3340 24090 3392
rect 25038 3340 25044 3392
rect 25096 3340 25102 3392
rect 25130 3340 25136 3392
rect 25188 3380 25194 3392
rect 26050 3380 26056 3392
rect 25188 3352 26056 3380
rect 25188 3340 25194 3352
rect 26050 3340 26056 3352
rect 26108 3380 26114 3392
rect 27157 3383 27215 3389
rect 27157 3380 27169 3383
rect 26108 3352 27169 3380
rect 26108 3340 26114 3352
rect 27157 3349 27169 3352
rect 27203 3349 27215 3383
rect 27157 3343 27215 3349
rect 27246 3340 27252 3392
rect 27304 3380 27310 3392
rect 28169 3383 28227 3389
rect 28169 3380 28181 3383
rect 27304 3352 28181 3380
rect 27304 3340 27310 3352
rect 28169 3349 28181 3352
rect 28215 3380 28227 3383
rect 29730 3380 29736 3392
rect 28215 3352 29736 3380
rect 28215 3349 28227 3352
rect 28169 3343 28227 3349
rect 29730 3340 29736 3352
rect 29788 3340 29794 3392
rect 31018 3340 31024 3392
rect 31076 3380 31082 3392
rect 32582 3380 32588 3392
rect 31076 3352 32588 3380
rect 31076 3340 31082 3352
rect 32582 3340 32588 3352
rect 32640 3340 32646 3392
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35618 3380 35624 3392
rect 34848 3352 35624 3380
rect 34848 3340 34854 3352
rect 35618 3340 35624 3352
rect 35676 3340 35682 3392
rect 36188 3380 36216 3411
rect 37936 3392 37964 3420
rect 39114 3408 39120 3460
rect 39172 3448 39178 3460
rect 39209 3451 39267 3457
rect 39209 3448 39221 3451
rect 39172 3420 39221 3448
rect 39172 3408 39178 3420
rect 39209 3417 39221 3420
rect 39255 3417 39267 3451
rect 39209 3411 39267 3417
rect 39390 3408 39396 3460
rect 39448 3448 39454 3460
rect 41877 3451 41935 3457
rect 41877 3448 41889 3451
rect 39448 3420 41889 3448
rect 39448 3408 39454 3420
rect 41877 3417 41889 3420
rect 41923 3417 41935 3451
rect 43898 3448 43904 3460
rect 41877 3411 41935 3417
rect 43640 3420 43904 3448
rect 37918 3380 37924 3392
rect 36188 3352 37924 3380
rect 37918 3340 37924 3352
rect 37976 3340 37982 3392
rect 38838 3340 38844 3392
rect 38896 3380 38902 3392
rect 39301 3383 39359 3389
rect 39301 3380 39313 3383
rect 38896 3352 39313 3380
rect 38896 3340 38902 3352
rect 39301 3349 39313 3352
rect 39347 3349 39359 3383
rect 39301 3343 39359 3349
rect 42978 3340 42984 3392
rect 43036 3380 43042 3392
rect 43640 3380 43668 3420
rect 43898 3408 43904 3420
rect 43956 3448 43962 3460
rect 44008 3448 44036 3479
rect 46106 3476 46112 3488
rect 46164 3476 46170 3528
rect 47578 3476 47584 3528
rect 47636 3516 47642 3528
rect 48501 3519 48559 3525
rect 48501 3516 48513 3519
rect 47636 3488 48513 3516
rect 47636 3476 47642 3488
rect 48501 3485 48513 3488
rect 48547 3485 48559 3519
rect 48501 3479 48559 3485
rect 48682 3476 48688 3528
rect 48740 3516 48746 3528
rect 49237 3519 49295 3525
rect 49237 3516 49249 3519
rect 48740 3488 49249 3516
rect 48740 3476 48746 3488
rect 49237 3485 49249 3488
rect 49283 3485 49295 3519
rect 49237 3479 49295 3485
rect 51258 3476 51264 3528
rect 51316 3516 51322 3528
rect 51905 3519 51963 3525
rect 51905 3516 51917 3519
rect 51316 3488 51917 3516
rect 51316 3476 51322 3488
rect 51905 3485 51917 3488
rect 51951 3485 51963 3519
rect 51905 3479 51963 3485
rect 53098 3476 53104 3528
rect 53156 3516 53162 3528
rect 54113 3519 54171 3525
rect 54113 3516 54125 3519
rect 53156 3488 54125 3516
rect 53156 3476 53162 3488
rect 54113 3485 54125 3488
rect 54159 3485 54171 3519
rect 54113 3479 54171 3485
rect 54754 3476 54760 3528
rect 54812 3516 54818 3528
rect 55493 3519 55551 3525
rect 55493 3516 55505 3519
rect 54812 3488 55505 3516
rect 54812 3476 54818 3488
rect 55493 3485 55505 3488
rect 55539 3485 55551 3519
rect 55493 3479 55551 3485
rect 43956 3420 44036 3448
rect 43956 3408 43962 3420
rect 44726 3408 44732 3460
rect 44784 3448 44790 3460
rect 45281 3451 45339 3457
rect 45281 3448 45293 3451
rect 44784 3420 45293 3448
rect 44784 3408 44790 3420
rect 45281 3417 45293 3420
rect 45327 3417 45339 3451
rect 45281 3411 45339 3417
rect 45370 3408 45376 3460
rect 45428 3448 45434 3460
rect 45428 3420 46244 3448
rect 45428 3408 45434 3420
rect 43036 3352 43668 3380
rect 43036 3340 43042 3352
rect 43714 3340 43720 3392
rect 43772 3380 43778 3392
rect 44174 3380 44180 3392
rect 43772 3352 44180 3380
rect 43772 3340 43778 3352
rect 44174 3340 44180 3352
rect 44232 3340 44238 3392
rect 46216 3380 46244 3420
rect 46750 3408 46756 3460
rect 46808 3448 46814 3460
rect 46937 3451 46995 3457
rect 46937 3448 46949 3451
rect 46808 3420 46949 3448
rect 46808 3408 46814 3420
rect 46937 3417 46949 3420
rect 46983 3417 46995 3451
rect 46937 3411 46995 3417
rect 47857 3451 47915 3457
rect 47857 3417 47869 3451
rect 47903 3417 47915 3451
rect 47857 3411 47915 3417
rect 47872 3380 47900 3411
rect 49786 3408 49792 3460
rect 49844 3448 49850 3460
rect 50433 3451 50491 3457
rect 50433 3448 50445 3451
rect 49844 3420 50445 3448
rect 49844 3408 49850 3420
rect 50433 3417 50445 3420
rect 50479 3417 50491 3451
rect 50433 3411 50491 3417
rect 50614 3408 50620 3460
rect 50672 3448 50678 3460
rect 51169 3451 51227 3457
rect 51169 3448 51181 3451
rect 50672 3420 51181 3448
rect 50672 3408 50678 3420
rect 51169 3417 51181 3420
rect 51215 3417 51227 3451
rect 51169 3411 51227 3417
rect 51718 3408 51724 3460
rect 51776 3448 51782 3460
rect 52641 3451 52699 3457
rect 52641 3448 52653 3451
rect 51776 3420 52653 3448
rect 51776 3408 51782 3420
rect 52641 3417 52653 3420
rect 52687 3417 52699 3451
rect 52641 3411 52699 3417
rect 53377 3451 53435 3457
rect 53377 3417 53389 3451
rect 53423 3417 53435 3451
rect 53377 3411 53435 3417
rect 46216 3352 47900 3380
rect 51074 3340 51080 3392
rect 51132 3380 51138 3392
rect 51261 3383 51319 3389
rect 51261 3380 51273 3383
rect 51132 3352 51273 3380
rect 51132 3340 51138 3352
rect 51261 3349 51273 3352
rect 51307 3349 51319 3383
rect 51261 3343 51319 3349
rect 52362 3340 52368 3392
rect 52420 3380 52426 3392
rect 53392 3380 53420 3411
rect 53742 3408 53748 3460
rect 53800 3448 53806 3460
rect 57118 3451 57176 3457
rect 57118 3448 57130 3451
rect 53800 3420 57130 3448
rect 53800 3408 53806 3420
rect 57118 3417 57130 3420
rect 57164 3417 57176 3451
rect 57118 3411 57176 3417
rect 52420 3352 53420 3380
rect 52420 3340 52426 3352
rect 53466 3340 53472 3392
rect 53524 3340 53530 3392
rect 57238 3340 57244 3392
rect 57296 3380 57302 3392
rect 58253 3383 58311 3389
rect 58253 3380 58265 3383
rect 57296 3352 58265 3380
rect 57296 3340 57302 3352
rect 58253 3349 58265 3352
rect 58299 3349 58311 3383
rect 58253 3343 58311 3349
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 5810 3176 5816 3188
rect 1596 3148 5816 3176
rect 1596 3049 1624 3148
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 6086 3176 6092 3188
rect 6012 3148 6092 3176
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 5166 3108 5172 3120
rect 4387 3080 5172 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 5166 3068 5172 3080
rect 5224 3068 5230 3120
rect 6012 3117 6040 3148
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 7098 3136 7104 3188
rect 7156 3176 7162 3188
rect 8570 3176 8576 3188
rect 7156 3148 8576 3176
rect 7156 3136 7162 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8849 3179 8907 3185
rect 8849 3145 8861 3179
rect 8895 3176 8907 3179
rect 9858 3176 9864 3188
rect 8895 3148 9864 3176
rect 8895 3145 8907 3148
rect 8849 3139 8907 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 12526 3136 12532 3188
rect 12584 3136 12590 3188
rect 13170 3136 13176 3188
rect 13228 3176 13234 3188
rect 13541 3179 13599 3185
rect 13541 3176 13553 3179
rect 13228 3148 13553 3176
rect 13228 3136 13234 3148
rect 13541 3145 13553 3148
rect 13587 3145 13599 3179
rect 15562 3176 15568 3188
rect 13541 3139 13599 3145
rect 14016 3148 15568 3176
rect 5997 3111 6055 3117
rect 5997 3077 6009 3111
rect 6043 3077 6055 3111
rect 5997 3071 6055 3077
rect 6932 3080 8156 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 6932 3040 6960 3080
rect 5859 3012 6960 3040
rect 7009 3043 7067 3049
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 7650 3040 7656 3052
rect 7055 3012 7656 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 934 2932 940 2984
rect 992 2972 998 2984
rect 1765 2975 1823 2981
rect 1765 2972 1777 2975
rect 992 2944 1777 2972
rect 992 2932 998 2944
rect 1765 2941 1777 2944
rect 1811 2941 1823 2975
rect 5092 2972 5120 3003
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3040 7803 3043
rect 8018 3040 8024 3052
rect 7791 3012 8024 3040
rect 7791 3009 7803 3012
rect 7745 3003 7803 3009
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 7558 2972 7564 2984
rect 5092 2944 7564 2972
rect 1765 2935 1823 2941
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 8128 2972 8156 3080
rect 8202 3068 8208 3120
rect 8260 3108 8266 3120
rect 8389 3111 8447 3117
rect 8389 3108 8401 3111
rect 8260 3080 8401 3108
rect 8260 3068 8266 3080
rect 8389 3077 8401 3080
rect 8435 3108 8447 3111
rect 8435 3080 9352 3108
rect 8435 3077 8447 3080
rect 8389 3071 8447 3077
rect 9214 3040 9220 3052
rect 8496 3012 9220 3040
rect 8496 2972 8524 3012
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 9324 3040 9352 3080
rect 9600 3080 13952 3108
rect 9324 3012 9444 3040
rect 8128 2944 8524 2972
rect 8588 2944 8800 2972
rect 5261 2907 5319 2913
rect 5261 2873 5273 2907
rect 5307 2904 5319 2907
rect 8588 2904 8616 2944
rect 5307 2876 8616 2904
rect 5307 2873 5319 2876
rect 5261 2867 5319 2873
rect 8662 2864 8668 2916
rect 8720 2864 8726 2916
rect 8772 2904 8800 2944
rect 9306 2932 9312 2984
rect 9364 2932 9370 2984
rect 9416 2972 9444 3012
rect 9490 3000 9496 3052
rect 9548 3000 9554 3052
rect 9600 3049 9628 3080
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 9766 3000 9772 3052
rect 9824 3000 9830 3052
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3040 12495 3043
rect 13722 3040 13728 3052
rect 12483 3012 13728 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 9677 2975 9735 2981
rect 9677 2972 9689 2975
rect 9416 2944 9689 2972
rect 9677 2941 9689 2944
rect 9723 2972 9735 2975
rect 10321 2975 10379 2981
rect 10321 2972 10333 2975
rect 9723 2944 10333 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 10321 2941 10333 2944
rect 10367 2941 10379 2975
rect 10321 2935 10379 2941
rect 13081 2975 13139 2981
rect 13081 2941 13093 2975
rect 13127 2972 13139 2975
rect 13262 2972 13268 2984
rect 13127 2944 13268 2972
rect 13127 2941 13139 2944
rect 13081 2935 13139 2941
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13538 2972 13544 2984
rect 13372 2944 13544 2972
rect 13372 2913 13400 2944
rect 13538 2932 13544 2944
rect 13596 2932 13602 2984
rect 13924 2972 13952 3080
rect 14016 3049 14044 3148
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 19058 3136 19064 3188
rect 19116 3176 19122 3188
rect 20346 3176 20352 3188
rect 19116 3148 20352 3176
rect 19116 3136 19122 3148
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 20438 3136 20444 3188
rect 20496 3176 20502 3188
rect 21085 3179 21143 3185
rect 21085 3176 21097 3179
rect 20496 3148 21097 3176
rect 20496 3136 20502 3148
rect 21085 3145 21097 3148
rect 21131 3145 21143 3179
rect 21085 3139 21143 3145
rect 23198 3136 23204 3188
rect 23256 3176 23262 3188
rect 23293 3179 23351 3185
rect 23293 3176 23305 3179
rect 23256 3148 23305 3176
rect 23256 3136 23262 3148
rect 23293 3145 23305 3148
rect 23339 3145 23351 3179
rect 23293 3139 23351 3145
rect 23658 3136 23664 3188
rect 23716 3136 23722 3188
rect 25038 3136 25044 3188
rect 25096 3176 25102 3188
rect 34238 3176 34244 3188
rect 25096 3148 34244 3176
rect 25096 3136 25102 3148
rect 34238 3136 34244 3148
rect 34296 3136 34302 3188
rect 34330 3136 34336 3188
rect 34388 3176 34394 3188
rect 34701 3179 34759 3185
rect 34701 3176 34713 3179
rect 34388 3148 34713 3176
rect 34388 3136 34394 3148
rect 34701 3145 34713 3148
rect 34747 3145 34759 3179
rect 34701 3139 34759 3145
rect 37642 3136 37648 3188
rect 37700 3176 37706 3188
rect 39390 3176 39396 3188
rect 37700 3148 39396 3176
rect 37700 3136 37706 3148
rect 39390 3136 39396 3148
rect 39448 3136 39454 3188
rect 39758 3136 39764 3188
rect 39816 3136 39822 3188
rect 40310 3136 40316 3188
rect 40368 3176 40374 3188
rect 40681 3179 40739 3185
rect 40681 3176 40693 3179
rect 40368 3148 40693 3176
rect 40368 3136 40374 3148
rect 40681 3145 40693 3148
rect 40727 3145 40739 3179
rect 40681 3139 40739 3145
rect 41782 3136 41788 3188
rect 41840 3136 41846 3188
rect 44358 3136 44364 3188
rect 44416 3176 44422 3188
rect 44453 3179 44511 3185
rect 44453 3176 44465 3179
rect 44416 3148 44465 3176
rect 44416 3136 44422 3148
rect 44453 3145 44465 3148
rect 44499 3145 44511 3179
rect 44453 3139 44511 3145
rect 44634 3136 44640 3188
rect 44692 3176 44698 3188
rect 45189 3179 45247 3185
rect 45189 3176 45201 3179
rect 44692 3148 45201 3176
rect 44692 3136 44698 3148
rect 45189 3145 45201 3148
rect 45235 3145 45247 3179
rect 45189 3139 45247 3145
rect 47486 3136 47492 3188
rect 47544 3176 47550 3188
rect 47949 3179 48007 3185
rect 47949 3176 47961 3179
rect 47544 3148 47961 3176
rect 47544 3136 47550 3148
rect 47949 3145 47961 3148
rect 47995 3145 48007 3179
rect 47949 3139 48007 3145
rect 48774 3136 48780 3188
rect 48832 3176 48838 3188
rect 48869 3179 48927 3185
rect 48869 3176 48881 3179
rect 48832 3148 48881 3176
rect 48832 3136 48838 3148
rect 48869 3145 48881 3148
rect 48915 3145 48927 3179
rect 48869 3139 48927 3145
rect 49789 3179 49847 3185
rect 49789 3145 49801 3179
rect 49835 3176 49847 3179
rect 49878 3176 49884 3188
rect 49835 3148 49884 3176
rect 49835 3145 49847 3148
rect 49789 3139 49847 3145
rect 49878 3136 49884 3148
rect 49936 3136 49942 3188
rect 52178 3136 52184 3188
rect 52236 3136 52242 3188
rect 54018 3136 54024 3188
rect 54076 3176 54082 3188
rect 54205 3179 54263 3185
rect 54205 3176 54217 3179
rect 54076 3148 54217 3176
rect 54076 3136 54082 3148
rect 54205 3145 54217 3148
rect 54251 3145 54263 3179
rect 54205 3139 54263 3145
rect 55214 3136 55220 3188
rect 55272 3176 55278 3188
rect 55309 3179 55367 3185
rect 55309 3176 55321 3179
rect 55272 3148 55321 3176
rect 55272 3136 55278 3148
rect 55309 3145 55321 3148
rect 55355 3145 55367 3179
rect 55309 3139 55367 3145
rect 57422 3136 57428 3188
rect 57480 3136 57486 3188
rect 23753 3111 23811 3117
rect 23753 3108 23765 3111
rect 14108 3080 23765 3108
rect 14001 3043 14059 3049
rect 14001 3009 14013 3043
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 14108 2972 14136 3080
rect 23753 3077 23765 3080
rect 23799 3108 23811 3111
rect 24026 3108 24032 3120
rect 23799 3080 24032 3108
rect 23799 3077 23811 3080
rect 23753 3071 23811 3077
rect 24026 3068 24032 3080
rect 24084 3068 24090 3120
rect 28534 3068 28540 3120
rect 28592 3068 28598 3120
rect 31294 3068 31300 3120
rect 31352 3108 31358 3120
rect 31352 3080 33364 3108
rect 31352 3068 31358 3080
rect 14458 3000 14464 3052
rect 14516 3040 14522 3052
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 14516 3012 14933 3040
rect 14516 3000 14522 3012
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 13924 2944 14136 2972
rect 14274 2932 14280 2984
rect 14332 2932 14338 2984
rect 14936 2972 14964 3003
rect 15838 3000 15844 3052
rect 15896 3000 15902 3052
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3040 17003 3043
rect 16991 3012 17816 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 15197 2975 15255 2981
rect 14936 2944 15056 2972
rect 10597 2907 10655 2913
rect 10597 2904 10609 2907
rect 8772 2876 10609 2904
rect 10597 2873 10609 2876
rect 10643 2873 10655 2907
rect 10597 2867 10655 2873
rect 10781 2907 10839 2913
rect 10781 2873 10793 2907
rect 10827 2904 10839 2907
rect 13357 2907 13415 2913
rect 10827 2876 13308 2904
rect 10827 2873 10839 2876
rect 10781 2867 10839 2873
rect 4433 2839 4491 2845
rect 4433 2805 4445 2839
rect 4479 2836 4491 2839
rect 6914 2836 6920 2848
rect 4479 2808 6920 2836
rect 4479 2805 4491 2808
rect 4433 2799 4491 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7101 2839 7159 2845
rect 7101 2805 7113 2839
rect 7147 2836 7159 2839
rect 7374 2836 7380 2848
rect 7147 2808 7380 2836
rect 7147 2805 7159 2808
rect 7101 2799 7159 2805
rect 7374 2796 7380 2808
rect 7432 2796 7438 2848
rect 7837 2839 7895 2845
rect 7837 2805 7849 2839
rect 7883 2836 7895 2839
rect 7926 2836 7932 2848
rect 7883 2808 7932 2836
rect 7883 2805 7895 2808
rect 7837 2799 7895 2805
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 8018 2796 8024 2848
rect 8076 2836 8082 2848
rect 10870 2836 10876 2848
rect 8076 2808 10876 2836
rect 8076 2796 8082 2808
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 13280 2836 13308 2876
rect 13357 2873 13369 2907
rect 13403 2873 13415 2907
rect 13357 2867 13415 2873
rect 14826 2836 14832 2848
rect 13280 2808 14832 2836
rect 14826 2796 14832 2808
rect 14884 2796 14890 2848
rect 15028 2836 15056 2944
rect 15197 2941 15209 2975
rect 15243 2972 15255 2975
rect 16022 2972 16028 2984
rect 15243 2944 16028 2972
rect 15243 2941 15255 2944
rect 15197 2935 15255 2941
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 16117 2975 16175 2981
rect 16117 2941 16129 2975
rect 16163 2972 16175 2975
rect 16298 2972 16304 2984
rect 16163 2944 16304 2972
rect 16163 2941 16175 2944
rect 16117 2935 16175 2941
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2972 17279 2975
rect 17586 2972 17592 2984
rect 17267 2944 17592 2972
rect 17267 2941 17279 2944
rect 17221 2935 17279 2941
rect 17586 2932 17592 2944
rect 17644 2932 17650 2984
rect 17788 2972 17816 3012
rect 17862 3000 17868 3052
rect 17920 3000 17926 3052
rect 18690 3000 18696 3052
rect 18748 3040 18754 3052
rect 18785 3043 18843 3049
rect 18785 3040 18797 3043
rect 18748 3012 18797 3040
rect 18748 3000 18754 3012
rect 18785 3009 18797 3012
rect 18831 3009 18843 3043
rect 18785 3003 18843 3009
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 19978 3049 19984 3052
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 19484 3012 19717 3040
rect 19484 3000 19490 3012
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 19972 3003 19984 3049
rect 19978 3000 19984 3003
rect 20036 3000 20042 3052
rect 20346 3000 20352 3052
rect 20404 3040 20410 3052
rect 21266 3040 21272 3052
rect 20404 3012 21272 3040
rect 20404 3000 20410 3012
rect 21266 3000 21272 3012
rect 21324 3000 21330 3052
rect 22373 3043 22431 3049
rect 22373 3009 22385 3043
rect 22419 3040 22431 3043
rect 22830 3040 22836 3052
rect 22419 3012 22836 3040
rect 22419 3009 22431 3012
rect 22373 3003 22431 3009
rect 22830 3000 22836 3012
rect 22888 3000 22894 3052
rect 25225 3043 25283 3049
rect 25225 3009 25237 3043
rect 25271 3040 25283 3043
rect 26145 3043 26203 3049
rect 25271 3012 26096 3040
rect 25271 3009 25283 3012
rect 25225 3003 25283 3009
rect 17954 2972 17960 2984
rect 17788 2944 17960 2972
rect 17954 2932 17960 2944
rect 18012 2932 18018 2984
rect 18138 2932 18144 2984
rect 18196 2932 18202 2984
rect 18966 2932 18972 2984
rect 19024 2932 19030 2984
rect 22649 2975 22707 2981
rect 22649 2941 22661 2975
rect 22695 2972 22707 2975
rect 23382 2972 23388 2984
rect 22695 2944 23388 2972
rect 22695 2941 22707 2944
rect 22649 2935 22707 2941
rect 23382 2932 23388 2944
rect 23440 2932 23446 2984
rect 23934 2932 23940 2984
rect 23992 2932 23998 2984
rect 25409 2975 25467 2981
rect 25409 2972 25421 2975
rect 25240 2944 25421 2972
rect 25240 2916 25268 2944
rect 25409 2941 25421 2944
rect 25455 2941 25467 2975
rect 25409 2935 25467 2941
rect 17494 2864 17500 2916
rect 17552 2904 17558 2916
rect 19426 2904 19432 2916
rect 17552 2876 19432 2904
rect 17552 2864 17558 2876
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 24946 2904 24952 2916
rect 22066 2876 24952 2904
rect 22066 2836 22094 2876
rect 24946 2864 24952 2876
rect 25004 2864 25010 2916
rect 25222 2864 25228 2916
rect 25280 2864 25286 2916
rect 26068 2904 26096 3012
rect 26145 3009 26157 3043
rect 26191 3040 26203 3043
rect 26970 3040 26976 3052
rect 26191 3012 26976 3040
rect 26191 3009 26203 3012
rect 26145 3003 26203 3009
rect 26970 3000 26976 3012
rect 27028 3000 27034 3052
rect 27522 3000 27528 3052
rect 27580 3000 27586 3052
rect 28442 3000 28448 3052
rect 28500 3000 28506 3052
rect 28552 3040 28580 3068
rect 28721 3043 28779 3049
rect 28721 3040 28733 3043
rect 28552 3012 28733 3040
rect 28721 3009 28733 3012
rect 28767 3009 28779 3043
rect 28721 3003 28779 3009
rect 30834 3000 30840 3052
rect 30892 3000 30898 3052
rect 33336 3049 33364 3080
rect 37918 3068 37924 3120
rect 37976 3068 37982 3120
rect 38562 3068 38568 3120
rect 38620 3108 38626 3120
rect 41046 3108 41052 3120
rect 38620 3080 41052 3108
rect 38620 3068 38626 3080
rect 41046 3068 41052 3080
rect 41104 3068 41110 3120
rect 42610 3068 42616 3120
rect 42668 3068 42674 3120
rect 43162 3068 43168 3120
rect 43220 3108 43226 3120
rect 44910 3108 44916 3120
rect 43220 3080 44916 3108
rect 43220 3068 43226 3080
rect 44910 3068 44916 3080
rect 44968 3068 44974 3120
rect 46753 3111 46811 3117
rect 46753 3077 46765 3111
rect 46799 3108 46811 3111
rect 47118 3108 47124 3120
rect 46799 3080 47124 3108
rect 46799 3077 46811 3080
rect 46753 3071 46811 3077
rect 47118 3068 47124 3080
rect 47176 3068 47182 3120
rect 49510 3068 49516 3120
rect 49568 3108 49574 3120
rect 50617 3111 50675 3117
rect 50617 3108 50629 3111
rect 49568 3080 50629 3108
rect 49568 3068 49574 3080
rect 50617 3077 50629 3080
rect 50663 3077 50675 3111
rect 50617 3071 50675 3077
rect 50890 3068 50896 3120
rect 50948 3108 50954 3120
rect 52089 3111 52147 3117
rect 52089 3108 52101 3111
rect 50948 3080 52101 3108
rect 50948 3068 50954 3080
rect 52089 3077 52101 3080
rect 52135 3077 52147 3111
rect 52089 3071 52147 3077
rect 53282 3068 53288 3120
rect 53340 3108 53346 3120
rect 56137 3111 56195 3117
rect 56137 3108 56149 3111
rect 53340 3080 56149 3108
rect 53340 3068 53346 3080
rect 56137 3077 56149 3080
rect 56183 3077 56195 3111
rect 56137 3071 56195 3077
rect 58158 3068 58164 3120
rect 58216 3068 58222 3120
rect 32309 3043 32367 3049
rect 32309 3040 32321 3043
rect 31128 3012 32321 3040
rect 26421 2975 26479 2981
rect 26421 2941 26433 2975
rect 26467 2972 26479 2975
rect 27338 2972 27344 2984
rect 26467 2944 27344 2972
rect 26467 2941 26479 2944
rect 26421 2935 26479 2941
rect 27338 2932 27344 2944
rect 27396 2932 27402 2984
rect 27798 2932 27804 2984
rect 27856 2932 27862 2984
rect 30558 2972 30564 2984
rect 28460 2944 30564 2972
rect 28460 2904 28488 2944
rect 30558 2932 30564 2944
rect 30616 2932 30622 2984
rect 30742 2932 30748 2984
rect 30800 2972 30806 2984
rect 31021 2975 31079 2981
rect 31021 2972 31033 2975
rect 30800 2944 31033 2972
rect 30800 2932 30806 2944
rect 31021 2941 31033 2944
rect 31067 2941 31079 2975
rect 31021 2935 31079 2941
rect 26068 2876 28488 2904
rect 29730 2864 29736 2916
rect 29788 2904 29794 2916
rect 29825 2907 29883 2913
rect 29825 2904 29837 2907
rect 29788 2876 29837 2904
rect 29788 2864 29794 2876
rect 29825 2873 29837 2876
rect 29871 2873 29883 2907
rect 29825 2867 29883 2873
rect 30098 2864 30104 2916
rect 30156 2904 30162 2916
rect 31128 2904 31156 3012
rect 32309 3009 32321 3012
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 33321 3043 33379 3049
rect 33321 3009 33333 3043
rect 33367 3040 33379 3043
rect 34514 3040 34520 3052
rect 33367 3012 34520 3040
rect 33367 3009 33379 3012
rect 33321 3003 33379 3009
rect 34514 3000 34520 3012
rect 34572 3000 34578 3052
rect 35434 3000 35440 3052
rect 35492 3000 35498 3052
rect 36170 3000 36176 3052
rect 36228 3040 36234 3052
rect 36357 3043 36415 3049
rect 36357 3040 36369 3043
rect 36228 3012 36369 3040
rect 36228 3000 36234 3012
rect 36357 3009 36369 3012
rect 36403 3009 36415 3043
rect 36357 3003 36415 3009
rect 37274 3000 37280 3052
rect 37332 3040 37338 3052
rect 37553 3043 37611 3049
rect 37553 3040 37565 3043
rect 37332 3012 37565 3040
rect 37332 3000 37338 3012
rect 37553 3009 37565 3012
rect 37599 3009 37611 3043
rect 37553 3003 37611 3009
rect 38654 3000 38660 3052
rect 38712 3000 38718 3052
rect 38856 3012 39068 3040
rect 31570 2932 31576 2984
rect 31628 2972 31634 2984
rect 32493 2975 32551 2981
rect 32493 2972 32505 2975
rect 31628 2944 32505 2972
rect 31628 2932 31634 2944
rect 32493 2941 32505 2944
rect 32539 2941 32551 2975
rect 32493 2935 32551 2941
rect 33594 2932 33600 2984
rect 33652 2932 33658 2984
rect 35618 2932 35624 2984
rect 35676 2932 35682 2984
rect 36538 2932 36544 2984
rect 36596 2932 36602 2984
rect 36906 2932 36912 2984
rect 36964 2972 36970 2984
rect 38856 2972 38884 3012
rect 36964 2944 38884 2972
rect 36964 2932 36970 2944
rect 38930 2932 38936 2984
rect 38988 2932 38994 2984
rect 30156 2876 31156 2904
rect 30156 2864 30162 2876
rect 38654 2864 38660 2916
rect 38712 2904 38718 2916
rect 38838 2904 38844 2916
rect 38712 2876 38844 2904
rect 38712 2864 38718 2876
rect 38838 2864 38844 2876
rect 38896 2864 38902 2916
rect 39040 2904 39068 3012
rect 39298 3000 39304 3052
rect 39356 3040 39362 3052
rect 39669 3043 39727 3049
rect 39669 3040 39681 3043
rect 39356 3012 39681 3040
rect 39356 3000 39362 3012
rect 39669 3009 39681 3012
rect 39715 3009 39727 3043
rect 39669 3003 39727 3009
rect 40126 3000 40132 3052
rect 40184 3040 40190 3052
rect 40589 3043 40647 3049
rect 40589 3040 40601 3043
rect 40184 3012 40601 3040
rect 40184 3000 40190 3012
rect 40589 3009 40601 3012
rect 40635 3009 40647 3043
rect 40589 3003 40647 3009
rect 41506 3000 41512 3052
rect 41564 3040 41570 3052
rect 41693 3043 41751 3049
rect 41693 3040 41705 3043
rect 41564 3012 41705 3040
rect 41564 3000 41570 3012
rect 41693 3009 41705 3012
rect 41739 3009 41751 3043
rect 41693 3003 41751 3009
rect 42978 3000 42984 3052
rect 43036 3040 43042 3052
rect 43254 3040 43260 3052
rect 43036 3012 43260 3040
rect 43036 3000 43042 3012
rect 43254 3000 43260 3012
rect 43312 3000 43318 3052
rect 43622 3000 43628 3052
rect 43680 3000 43686 3052
rect 43806 3000 43812 3052
rect 43864 3040 43870 3052
rect 44361 3043 44419 3049
rect 44361 3040 44373 3043
rect 43864 3012 44373 3040
rect 43864 3000 43870 3012
rect 44361 3009 44373 3012
rect 44407 3009 44419 3043
rect 44361 3003 44419 3009
rect 45002 3000 45008 3052
rect 45060 3000 45066 3052
rect 46198 3000 46204 3052
rect 46256 3040 46262 3052
rect 46385 3043 46443 3049
rect 46385 3040 46397 3043
rect 46256 3012 46397 3040
rect 46256 3000 46262 3012
rect 46385 3009 46397 3012
rect 46431 3009 46443 3043
rect 46385 3003 46443 3009
rect 47026 3000 47032 3052
rect 47084 3040 47090 3052
rect 47857 3043 47915 3049
rect 47857 3040 47869 3043
rect 47084 3012 47869 3040
rect 47084 3000 47090 3012
rect 47857 3009 47869 3012
rect 47903 3009 47915 3043
rect 47857 3003 47915 3009
rect 48406 3000 48412 3052
rect 48464 3040 48470 3052
rect 48777 3043 48835 3049
rect 48777 3040 48789 3043
rect 48464 3012 48789 3040
rect 48464 3000 48470 3012
rect 48777 3009 48789 3012
rect 48823 3009 48835 3043
rect 48777 3003 48835 3009
rect 48958 3000 48964 3052
rect 49016 3040 49022 3052
rect 49697 3043 49755 3049
rect 49697 3040 49709 3043
rect 49016 3012 49709 3040
rect 49016 3000 49022 3012
rect 49697 3009 49709 3012
rect 49743 3009 49755 3043
rect 49697 3003 49755 3009
rect 49804 3012 50936 3040
rect 40770 2932 40776 2984
rect 40828 2972 40834 2984
rect 42996 2972 43024 3000
rect 40828 2944 43024 2972
rect 43349 2975 43407 2981
rect 40828 2932 40834 2944
rect 43349 2941 43361 2975
rect 43395 2941 43407 2975
rect 43349 2935 43407 2941
rect 41230 2904 41236 2916
rect 39040 2876 41236 2904
rect 41230 2864 41236 2876
rect 41288 2864 41294 2916
rect 43364 2904 43392 2935
rect 43438 2932 43444 2984
rect 43496 2972 43502 2984
rect 43533 2975 43591 2981
rect 43533 2972 43545 2975
rect 43496 2944 43545 2972
rect 43496 2932 43502 2944
rect 43533 2941 43545 2944
rect 43579 2972 43591 2975
rect 43898 2972 43904 2984
rect 43579 2944 43904 2972
rect 43579 2941 43591 2944
rect 43533 2935 43591 2941
rect 43898 2932 43904 2944
rect 43956 2932 43962 2984
rect 45278 2932 45284 2984
rect 45336 2972 45342 2984
rect 49804 2972 49832 3012
rect 45336 2944 49832 2972
rect 45336 2932 45342 2944
rect 50801 2907 50859 2913
rect 50801 2904 50813 2907
rect 43364 2876 50813 2904
rect 50801 2873 50813 2876
rect 50847 2873 50859 2907
rect 50908 2904 50936 3012
rect 50982 3000 50988 3052
rect 51040 3040 51046 3052
rect 51353 3043 51411 3049
rect 51353 3040 51365 3043
rect 51040 3012 51365 3040
rect 51040 3000 51046 3012
rect 51353 3009 51365 3012
rect 51399 3009 51411 3043
rect 51353 3003 51411 3009
rect 51442 3000 51448 3052
rect 51500 3040 51506 3052
rect 53009 3043 53067 3049
rect 53009 3040 53021 3043
rect 51500 3012 53021 3040
rect 51500 3000 51506 3012
rect 53009 3009 53021 3012
rect 53055 3009 53067 3043
rect 53009 3003 53067 3009
rect 53926 3000 53932 3052
rect 53984 3040 53990 3052
rect 54113 3043 54171 3049
rect 54113 3040 54125 3043
rect 53984 3012 54125 3040
rect 53984 3000 53990 3012
rect 54113 3009 54125 3012
rect 54159 3009 54171 3043
rect 54113 3003 54171 3009
rect 54202 3000 54208 3052
rect 54260 3040 54266 3052
rect 55033 3043 55091 3049
rect 55033 3040 55045 3043
rect 54260 3012 55045 3040
rect 54260 3000 54266 3012
rect 55033 3009 55045 3012
rect 55079 3009 55091 3043
rect 55033 3003 55091 3009
rect 55306 3000 55312 3052
rect 55364 3040 55370 3052
rect 55861 3043 55919 3049
rect 55861 3040 55873 3043
rect 55364 3012 55873 3040
rect 55364 3000 55370 3012
rect 55861 3009 55873 3012
rect 55907 3009 55919 3043
rect 55861 3003 55919 3009
rect 57241 3043 57299 3049
rect 57241 3009 57253 3043
rect 57287 3040 57299 3043
rect 58250 3040 58256 3052
rect 57287 3012 58256 3040
rect 57287 3009 57299 3012
rect 57241 3003 57299 3009
rect 58250 3000 58256 3012
rect 58308 3000 58314 3052
rect 52086 2932 52092 2984
rect 52144 2972 52150 2984
rect 53193 2975 53251 2981
rect 53193 2972 53205 2975
rect 52144 2944 53205 2972
rect 52144 2932 52150 2944
rect 53193 2941 53205 2944
rect 53239 2941 53251 2975
rect 53193 2935 53251 2941
rect 57057 2975 57115 2981
rect 57057 2941 57069 2975
rect 57103 2972 57115 2975
rect 58345 2975 58403 2981
rect 58345 2972 58357 2975
rect 57103 2944 58357 2972
rect 57103 2941 57115 2944
rect 57057 2935 57115 2941
rect 58345 2941 58357 2944
rect 58391 2941 58403 2975
rect 58345 2935 58403 2941
rect 51537 2907 51595 2913
rect 51537 2904 51549 2907
rect 50908 2876 51549 2904
rect 50801 2867 50859 2873
rect 51537 2873 51549 2876
rect 51583 2873 51595 2907
rect 51537 2867 51595 2873
rect 15028 2808 22094 2836
rect 24765 2839 24823 2845
rect 24765 2805 24777 2839
rect 24811 2836 24823 2839
rect 26602 2836 26608 2848
rect 24811 2808 26608 2836
rect 24811 2805 24823 2808
rect 24765 2799 24823 2805
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 27522 2796 27528 2848
rect 27580 2836 27586 2848
rect 29086 2836 29092 2848
rect 27580 2808 29092 2836
rect 27580 2796 27586 2808
rect 29086 2796 29092 2808
rect 29144 2796 29150 2848
rect 37458 2796 37464 2848
rect 37516 2836 37522 2848
rect 40034 2836 40040 2848
rect 37516 2808 40040 2836
rect 37516 2796 37522 2808
rect 40034 2796 40040 2808
rect 40092 2796 40098 2848
rect 43070 2796 43076 2848
rect 43128 2836 43134 2848
rect 49694 2836 49700 2848
rect 43128 2808 49700 2836
rect 43128 2796 43134 2808
rect 49694 2796 49700 2808
rect 49752 2796 49758 2848
rect 50154 2796 50160 2848
rect 50212 2836 50218 2848
rect 50982 2836 50988 2848
rect 50212 2808 50988 2836
rect 50212 2796 50218 2808
rect 50982 2796 50988 2808
rect 51040 2796 51046 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 7190 2632 7196 2644
rect 3375 2604 7196 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 8478 2592 8484 2644
rect 8536 2592 8542 2644
rect 13630 2632 13636 2644
rect 10336 2604 13636 2632
rect 5997 2567 6055 2573
rect 5997 2533 6009 2567
rect 6043 2564 6055 2567
rect 7834 2564 7840 2576
rect 6043 2536 7840 2564
rect 6043 2533 6055 2536
rect 5997 2527 6055 2533
rect 7834 2524 7840 2536
rect 7892 2524 7898 2576
rect 8386 2524 8392 2576
rect 8444 2524 8450 2576
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2496 4583 2499
rect 8404 2496 8432 2524
rect 4571 2468 8432 2496
rect 4571 2465 4583 2468
rect 4525 2459 4583 2465
rect 1578 2388 1584 2440
rect 1636 2388 1642 2440
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 7834 2428 7840 2440
rect 4387 2400 7840 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 10134 2428 10140 2440
rect 8435 2400 10140 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2428 10287 2431
rect 10336 2428 10364 2604
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 14461 2635 14519 2641
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 17402 2632 17408 2644
rect 14507 2604 17408 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 17954 2592 17960 2644
rect 18012 2632 18018 2644
rect 19058 2632 19064 2644
rect 18012 2604 19064 2632
rect 18012 2592 18018 2604
rect 19058 2592 19064 2604
rect 19116 2592 19122 2644
rect 19978 2592 19984 2644
rect 20036 2592 20042 2644
rect 22189 2635 22247 2641
rect 22189 2601 22201 2635
rect 22235 2632 22247 2635
rect 25774 2632 25780 2644
rect 22235 2604 25780 2632
rect 22235 2601 22247 2604
rect 22189 2595 22247 2601
rect 25774 2592 25780 2604
rect 25832 2592 25838 2644
rect 25958 2592 25964 2644
rect 26016 2632 26022 2644
rect 26016 2604 30420 2632
rect 26016 2592 26022 2604
rect 10413 2567 10471 2573
rect 10413 2533 10425 2567
rect 10459 2564 10471 2567
rect 11054 2564 11060 2576
rect 10459 2536 11060 2564
rect 10459 2533 10471 2536
rect 10413 2527 10471 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 11149 2567 11207 2573
rect 11149 2533 11161 2567
rect 11195 2564 11207 2567
rect 14642 2564 14648 2576
rect 11195 2536 14648 2564
rect 11195 2533 11207 2536
rect 11149 2527 11207 2533
rect 14642 2524 14648 2536
rect 14700 2524 14706 2576
rect 21358 2564 21364 2576
rect 18432 2536 21364 2564
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 15010 2496 15016 2508
rect 12667 2468 15016 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 15010 2456 15016 2468
rect 15068 2456 15074 2508
rect 17037 2499 17095 2505
rect 17037 2465 17049 2499
rect 17083 2496 17095 2499
rect 17770 2496 17776 2508
rect 17083 2468 17776 2496
rect 17083 2465 17095 2468
rect 17037 2459 17095 2465
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 11238 2428 11244 2440
rect 10275 2400 10364 2428
rect 10428 2400 11244 2428
rect 10275 2397 10287 2400
rect 10229 2391 10287 2397
rect 934 2320 940 2372
rect 992 2360 998 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 992 2332 1869 2360
rect 992 2320 998 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 3234 2320 3240 2372
rect 3292 2320 3298 2372
rect 5077 2363 5135 2369
rect 5077 2329 5089 2363
rect 5123 2360 5135 2363
rect 5123 2332 5764 2360
rect 5123 2329 5135 2332
rect 5077 2323 5135 2329
rect 5169 2295 5227 2301
rect 5169 2261 5181 2295
rect 5215 2292 5227 2295
rect 5350 2292 5356 2304
rect 5215 2264 5356 2292
rect 5215 2261 5227 2264
rect 5169 2255 5227 2261
rect 5350 2252 5356 2264
rect 5408 2252 5414 2304
rect 5736 2292 5764 2332
rect 5810 2320 5816 2372
rect 5868 2320 5874 2372
rect 6914 2320 6920 2372
rect 6972 2320 6978 2372
rect 7098 2320 7104 2372
rect 7156 2320 7162 2372
rect 7650 2320 7656 2372
rect 7708 2320 7714 2372
rect 9493 2363 9551 2369
rect 9493 2329 9505 2363
rect 9539 2329 9551 2363
rect 9493 2323 9551 2329
rect 9677 2363 9735 2369
rect 9677 2329 9689 2363
rect 9723 2360 9735 2363
rect 10428 2360 10456 2400
rect 11238 2388 11244 2400
rect 11296 2388 11302 2440
rect 12342 2388 12348 2440
rect 12400 2388 12406 2440
rect 12986 2388 12992 2440
rect 13044 2428 13050 2440
rect 13265 2431 13323 2437
rect 13265 2428 13277 2431
rect 13044 2400 13277 2428
rect 13044 2388 13050 2400
rect 13265 2397 13277 2400
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 14918 2388 14924 2440
rect 14976 2388 14982 2440
rect 15470 2388 15476 2440
rect 15528 2428 15534 2440
rect 15841 2431 15899 2437
rect 15841 2428 15853 2431
rect 15528 2400 15853 2428
rect 15528 2388 15534 2400
rect 15841 2397 15853 2400
rect 15887 2397 15899 2431
rect 15841 2391 15899 2397
rect 17494 2388 17500 2440
rect 17552 2388 17558 2440
rect 18432 2437 18460 2536
rect 21358 2524 21364 2536
rect 21416 2524 21422 2576
rect 22664 2536 28856 2564
rect 20438 2456 20444 2508
rect 20496 2456 20502 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 21174 2496 21180 2508
rect 20671 2468 21180 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 21174 2456 21180 2468
rect 21232 2456 21238 2508
rect 18417 2431 18475 2437
rect 17696 2400 18368 2428
rect 9723 2332 10456 2360
rect 10965 2363 11023 2369
rect 9723 2329 9735 2332
rect 9677 2323 9735 2329
rect 10965 2329 10977 2363
rect 11011 2360 11023 2363
rect 13446 2360 13452 2372
rect 11011 2332 13452 2360
rect 11011 2329 11023 2332
rect 10965 2323 11023 2329
rect 6822 2292 6828 2304
rect 5736 2264 6828 2292
rect 6822 2252 6828 2264
rect 6880 2252 6886 2304
rect 7742 2252 7748 2304
rect 7800 2252 7806 2304
rect 9508 2292 9536 2323
rect 13446 2320 13452 2332
rect 13504 2320 13510 2372
rect 13541 2363 13599 2369
rect 13541 2329 13553 2363
rect 13587 2329 13599 2363
rect 13541 2323 13599 2329
rect 15197 2363 15255 2369
rect 15197 2329 15209 2363
rect 15243 2360 15255 2363
rect 16117 2363 16175 2369
rect 15243 2332 16068 2360
rect 15243 2329 15255 2332
rect 15197 2323 15255 2329
rect 11054 2292 11060 2304
rect 9508 2264 11060 2292
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 13556 2292 13584 2323
rect 15838 2292 15844 2304
rect 13556 2264 15844 2292
rect 15838 2252 15844 2264
rect 15896 2252 15902 2304
rect 16040 2292 16068 2332
rect 16117 2329 16129 2363
rect 16163 2360 16175 2363
rect 17696 2360 17724 2400
rect 16163 2332 17724 2360
rect 17773 2363 17831 2369
rect 16163 2329 16175 2332
rect 16117 2323 16175 2329
rect 17773 2329 17785 2363
rect 17819 2360 17831 2363
rect 18230 2360 18236 2372
rect 17819 2332 18236 2360
rect 17819 2329 17831 2332
rect 17773 2323 17831 2329
rect 18230 2320 18236 2332
rect 18288 2320 18294 2372
rect 18340 2360 18368 2400
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 20254 2428 20260 2440
rect 18417 2391 18475 2397
rect 18616 2400 20260 2428
rect 18616 2360 18644 2400
rect 20254 2388 20260 2400
rect 20312 2388 20318 2440
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2428 20407 2431
rect 20530 2428 20536 2440
rect 20395 2400 20536 2428
rect 20395 2397 20407 2400
rect 20349 2391 20407 2397
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 22094 2428 22100 2440
rect 21315 2400 22100 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 22094 2388 22100 2400
rect 22152 2388 22158 2440
rect 22664 2437 22692 2536
rect 24581 2499 24639 2505
rect 24581 2465 24593 2499
rect 24627 2496 24639 2499
rect 27430 2496 27436 2508
rect 24627 2468 27436 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 27430 2456 27436 2468
rect 27488 2456 27494 2508
rect 28166 2496 28172 2508
rect 27724 2468 28172 2496
rect 22649 2431 22707 2437
rect 22649 2397 22661 2431
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 23474 2388 23480 2440
rect 23532 2428 23538 2440
rect 23569 2431 23627 2437
rect 23569 2428 23581 2431
rect 23532 2400 23581 2428
rect 23532 2388 23538 2400
rect 23569 2397 23581 2400
rect 23615 2397 23627 2431
rect 23569 2391 23627 2397
rect 23658 2388 23664 2440
rect 23716 2428 23722 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 23716 2400 25237 2428
rect 23716 2388 23722 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2428 26203 2431
rect 27724 2428 27752 2468
rect 28166 2456 28172 2468
rect 28224 2456 28230 2508
rect 28828 2496 28856 2536
rect 28902 2524 28908 2576
rect 28960 2564 28966 2576
rect 30282 2564 30288 2576
rect 28960 2536 30288 2564
rect 28960 2524 28966 2536
rect 30282 2524 30288 2536
rect 30340 2524 30346 2576
rect 30392 2496 30420 2604
rect 30466 2592 30472 2644
rect 30524 2632 30530 2644
rect 43073 2635 43131 2641
rect 30524 2604 41414 2632
rect 30524 2592 30530 2604
rect 32122 2524 32128 2576
rect 32180 2564 32186 2576
rect 32180 2536 35848 2564
rect 32180 2524 32186 2536
rect 28828 2468 30328 2496
rect 30392 2468 32352 2496
rect 26191 2400 27752 2428
rect 27801 2431 27859 2437
rect 26191 2397 26203 2400
rect 26145 2391 26203 2397
rect 27801 2397 27813 2431
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 18340 2332 18644 2360
rect 18693 2363 18751 2369
rect 18693 2329 18705 2363
rect 18739 2360 18751 2363
rect 20714 2360 20720 2372
rect 18739 2332 20720 2360
rect 18739 2329 18751 2332
rect 18693 2323 18751 2329
rect 20714 2320 20720 2332
rect 20772 2320 20778 2372
rect 22925 2363 22983 2369
rect 22925 2329 22937 2363
rect 22971 2360 22983 2363
rect 23198 2360 23204 2372
rect 22971 2332 23204 2360
rect 22971 2329 22983 2332
rect 22925 2323 22983 2329
rect 23198 2320 23204 2332
rect 23256 2320 23262 2372
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 24762 2360 24768 2372
rect 23891 2332 24768 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 24762 2320 24768 2332
rect 24820 2320 24826 2372
rect 25498 2320 25504 2372
rect 25556 2320 25562 2372
rect 26418 2320 26424 2372
rect 26476 2320 26482 2372
rect 27614 2320 27620 2372
rect 27672 2360 27678 2372
rect 27816 2360 27844 2391
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28721 2431 28779 2437
rect 28721 2428 28733 2431
rect 28408 2400 28733 2428
rect 28408 2388 28414 2400
rect 28721 2397 28733 2400
rect 28767 2397 28779 2431
rect 28721 2391 28779 2397
rect 30006 2388 30012 2440
rect 30064 2428 30070 2440
rect 30193 2431 30251 2437
rect 30193 2428 30205 2431
rect 30064 2400 30205 2428
rect 30064 2388 30070 2400
rect 30193 2397 30205 2400
rect 30239 2397 30251 2431
rect 30193 2391 30251 2397
rect 27672 2332 27844 2360
rect 27672 2320 27678 2332
rect 18874 2292 18880 2304
rect 16040 2264 18880 2292
rect 18874 2252 18880 2264
rect 18932 2252 18938 2304
rect 19058 2252 19064 2304
rect 19116 2292 19122 2304
rect 21361 2295 21419 2301
rect 21361 2292 21373 2295
rect 19116 2264 21373 2292
rect 19116 2252 19122 2264
rect 21361 2261 21373 2264
rect 21407 2261 21419 2295
rect 21361 2255 21419 2261
rect 27157 2295 27215 2301
rect 27157 2261 27169 2295
rect 27203 2292 27215 2295
rect 27522 2292 27528 2304
rect 27203 2264 27528 2292
rect 27203 2261 27215 2264
rect 27157 2255 27215 2261
rect 27522 2252 27528 2264
rect 27580 2252 27586 2304
rect 27816 2292 27844 2332
rect 28077 2363 28135 2369
rect 28077 2329 28089 2363
rect 28123 2360 28135 2363
rect 28902 2360 28908 2372
rect 28123 2332 28908 2360
rect 28123 2329 28135 2332
rect 28077 2323 28135 2329
rect 28902 2320 28908 2332
rect 28960 2320 28966 2372
rect 28997 2363 29055 2369
rect 28997 2329 29009 2363
rect 29043 2360 29055 2363
rect 29914 2360 29920 2372
rect 29043 2332 29920 2360
rect 29043 2329 29055 2332
rect 28997 2323 29055 2329
rect 29914 2320 29920 2332
rect 29972 2320 29978 2372
rect 29822 2292 29828 2304
rect 27816 2264 29828 2292
rect 29822 2252 29828 2264
rect 29880 2252 29886 2304
rect 30300 2292 30328 2468
rect 31110 2388 31116 2440
rect 31168 2388 31174 2440
rect 32324 2437 32352 2468
rect 32309 2431 32367 2437
rect 32309 2397 32321 2431
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 32490 2388 32496 2440
rect 32548 2428 32554 2440
rect 33229 2431 33287 2437
rect 33229 2428 33241 2431
rect 32548 2400 33241 2428
rect 32548 2388 32554 2400
rect 33229 2397 33241 2400
rect 33275 2397 33287 2431
rect 33229 2391 33287 2397
rect 34882 2388 34888 2440
rect 34940 2388 34946 2440
rect 35820 2437 35848 2536
rect 39482 2524 39488 2576
rect 39540 2564 39546 2576
rect 41233 2567 41291 2573
rect 41233 2564 41245 2567
rect 39540 2536 41245 2564
rect 39540 2524 39546 2536
rect 41233 2533 41245 2536
rect 41279 2533 41291 2567
rect 41233 2527 41291 2533
rect 38654 2496 38660 2508
rect 37476 2468 38660 2496
rect 37476 2437 37504 2468
rect 38654 2456 38660 2468
rect 38712 2456 38718 2508
rect 35805 2431 35863 2437
rect 35805 2397 35817 2431
rect 35851 2397 35863 2431
rect 35805 2391 35863 2397
rect 37461 2431 37519 2437
rect 37461 2397 37473 2431
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 38381 2431 38439 2437
rect 38381 2397 38393 2431
rect 38427 2397 38439 2431
rect 38381 2391 38439 2397
rect 30466 2320 30472 2372
rect 30524 2320 30530 2372
rect 31018 2320 31024 2372
rect 31076 2360 31082 2372
rect 31389 2363 31447 2369
rect 31389 2360 31401 2363
rect 31076 2332 31401 2360
rect 31076 2320 31082 2332
rect 31389 2329 31401 2332
rect 31435 2329 31447 2363
rect 31389 2323 31447 2329
rect 32582 2320 32588 2372
rect 32640 2320 32646 2372
rect 33502 2320 33508 2372
rect 33560 2320 33566 2372
rect 35158 2320 35164 2372
rect 35216 2320 35222 2372
rect 36078 2320 36084 2372
rect 36136 2320 36142 2372
rect 37734 2320 37740 2372
rect 37792 2320 37798 2372
rect 32214 2292 32220 2304
rect 30300 2264 32220 2292
rect 32214 2252 32220 2264
rect 32272 2252 32278 2304
rect 35434 2252 35440 2304
rect 35492 2292 35498 2304
rect 38396 2292 38424 2391
rect 39114 2388 39120 2440
rect 39172 2428 39178 2440
rect 40037 2431 40095 2437
rect 40037 2428 40049 2431
rect 39172 2400 40049 2428
rect 39172 2388 39178 2400
rect 40037 2397 40049 2400
rect 40083 2397 40095 2431
rect 40037 2391 40095 2397
rect 38654 2320 38660 2372
rect 38712 2320 38718 2372
rect 38838 2320 38844 2372
rect 38896 2360 38902 2372
rect 40313 2363 40371 2369
rect 40313 2360 40325 2363
rect 38896 2332 40325 2360
rect 38896 2320 38902 2332
rect 40313 2329 40325 2332
rect 40359 2329 40371 2363
rect 40313 2323 40371 2329
rect 41046 2320 41052 2372
rect 41104 2320 41110 2372
rect 41386 2360 41414 2604
rect 43073 2601 43085 2635
rect 43119 2632 43131 2635
rect 44082 2632 44088 2644
rect 43119 2604 44088 2632
rect 43119 2601 43131 2604
rect 43073 2595 43131 2601
rect 44082 2592 44088 2604
rect 44140 2592 44146 2644
rect 44174 2592 44180 2644
rect 44232 2632 44238 2644
rect 45373 2635 45431 2641
rect 45373 2632 45385 2635
rect 44232 2604 45385 2632
rect 44232 2592 44238 2604
rect 45373 2601 45385 2604
rect 45419 2601 45431 2635
rect 45373 2595 45431 2601
rect 45830 2592 45836 2644
rect 45888 2632 45894 2644
rect 46201 2635 46259 2641
rect 46201 2632 46213 2635
rect 45888 2604 46213 2632
rect 45888 2592 45894 2604
rect 46201 2601 46213 2604
rect 46247 2601 46259 2635
rect 46201 2595 46259 2601
rect 47394 2592 47400 2644
rect 47452 2632 47458 2644
rect 47949 2635 48007 2641
rect 47949 2632 47961 2635
rect 47452 2604 47961 2632
rect 47452 2592 47458 2604
rect 47949 2601 47961 2604
rect 47995 2601 48007 2635
rect 47949 2595 48007 2601
rect 48866 2592 48872 2644
rect 48924 2592 48930 2644
rect 49694 2592 49700 2644
rect 49752 2632 49758 2644
rect 51997 2635 52055 2641
rect 51997 2632 52009 2635
rect 49752 2604 52009 2632
rect 49752 2592 49758 2604
rect 51997 2601 52009 2604
rect 52043 2601 52055 2635
rect 51997 2595 52055 2601
rect 58250 2592 58256 2644
rect 58308 2592 58314 2644
rect 51074 2564 51080 2576
rect 43088 2536 51080 2564
rect 43088 2428 43116 2536
rect 51074 2524 51080 2536
rect 51132 2524 51138 2576
rect 53466 2564 53472 2576
rect 51184 2536 53472 2564
rect 51184 2496 51212 2536
rect 53466 2524 53472 2536
rect 53524 2524 53530 2576
rect 43548 2468 51212 2496
rect 43257 2431 43315 2437
rect 43257 2428 43269 2431
rect 43088 2400 43269 2428
rect 43257 2397 43269 2400
rect 43303 2397 43315 2431
rect 43257 2391 43315 2397
rect 43346 2388 43352 2440
rect 43404 2428 43410 2440
rect 43441 2431 43499 2437
rect 43441 2428 43453 2431
rect 43404 2400 43453 2428
rect 43404 2388 43410 2400
rect 43441 2397 43453 2400
rect 43487 2397 43499 2431
rect 43441 2391 43499 2397
rect 43548 2360 43576 2468
rect 51810 2456 51816 2508
rect 51868 2496 51874 2508
rect 54021 2499 54079 2505
rect 54021 2496 54033 2499
rect 51868 2468 54033 2496
rect 51868 2456 51874 2468
rect 54021 2465 54033 2468
rect 54067 2465 54079 2499
rect 54021 2459 54079 2465
rect 55674 2456 55680 2508
rect 55732 2456 55738 2508
rect 43809 2431 43867 2437
rect 43809 2397 43821 2431
rect 43855 2397 43867 2431
rect 43809 2391 43867 2397
rect 41386 2332 43576 2360
rect 43824 2360 43852 2391
rect 43898 2388 43904 2440
rect 43956 2388 43962 2440
rect 44082 2388 44088 2440
rect 44140 2428 44146 2440
rect 51353 2431 51411 2437
rect 51353 2428 51365 2431
rect 44140 2400 51365 2428
rect 44140 2388 44146 2400
rect 51353 2397 51365 2400
rect 51399 2397 51411 2431
rect 51353 2391 51411 2397
rect 53834 2388 53840 2440
rect 53892 2388 53898 2440
rect 55214 2388 55220 2440
rect 55272 2428 55278 2440
rect 55493 2431 55551 2437
rect 55493 2428 55505 2431
rect 55272 2400 55505 2428
rect 55272 2388 55278 2400
rect 55493 2397 55505 2400
rect 55539 2397 55551 2431
rect 55493 2391 55551 2397
rect 57057 2431 57115 2437
rect 57057 2397 57069 2431
rect 57103 2428 57115 2431
rect 57238 2428 57244 2440
rect 57103 2400 57244 2428
rect 57103 2397 57115 2400
rect 57057 2391 57115 2397
rect 57238 2388 57244 2400
rect 57296 2388 57302 2440
rect 58161 2431 58219 2437
rect 58161 2397 58173 2431
rect 58207 2428 58219 2431
rect 58986 2428 58992 2440
rect 58207 2400 58992 2428
rect 58207 2397 58219 2400
rect 58161 2391 58219 2397
rect 58986 2388 58992 2400
rect 59044 2388 59050 2440
rect 45186 2360 45192 2372
rect 43824 2332 45192 2360
rect 45186 2320 45192 2332
rect 45244 2320 45250 2372
rect 45278 2320 45284 2372
rect 45336 2320 45342 2372
rect 45922 2320 45928 2372
rect 45980 2360 45986 2372
rect 46109 2363 46167 2369
rect 46109 2360 46121 2363
rect 45980 2332 46121 2360
rect 45980 2320 45986 2332
rect 46109 2329 46121 2332
rect 46155 2329 46167 2363
rect 46109 2323 46167 2329
rect 46290 2320 46296 2372
rect 46348 2360 46354 2372
rect 47029 2363 47087 2369
rect 47029 2360 47041 2363
rect 46348 2332 47041 2360
rect 46348 2320 46354 2332
rect 47029 2329 47041 2332
rect 47075 2329 47087 2363
rect 47029 2323 47087 2329
rect 47394 2320 47400 2372
rect 47452 2360 47458 2372
rect 47857 2363 47915 2369
rect 47857 2360 47869 2363
rect 47452 2332 47869 2360
rect 47452 2320 47458 2332
rect 47857 2329 47869 2332
rect 47903 2329 47915 2363
rect 47857 2323 47915 2329
rect 48774 2320 48780 2372
rect 48832 2320 48838 2372
rect 49694 2320 49700 2372
rect 49752 2360 49758 2372
rect 50433 2363 50491 2369
rect 50433 2360 50445 2363
rect 49752 2332 50445 2360
rect 49752 2320 49758 2332
rect 50433 2329 50445 2332
rect 50479 2329 50491 2363
rect 50433 2323 50491 2329
rect 51074 2320 51080 2372
rect 51132 2360 51138 2372
rect 51169 2363 51227 2369
rect 51169 2360 51181 2363
rect 51132 2332 51181 2360
rect 51132 2320 51138 2332
rect 51169 2329 51181 2332
rect 51215 2329 51227 2363
rect 51169 2323 51227 2329
rect 51902 2320 51908 2372
rect 51960 2320 51966 2372
rect 52546 2320 52552 2372
rect 52604 2360 52610 2372
rect 53009 2363 53067 2369
rect 53009 2360 53021 2363
rect 52604 2332 53021 2360
rect 52604 2320 52610 2332
rect 53009 2329 53021 2332
rect 53055 2329 53067 2363
rect 53009 2323 53067 2329
rect 57333 2363 57391 2369
rect 57333 2329 57345 2363
rect 57379 2360 57391 2363
rect 58894 2360 58900 2372
rect 57379 2332 58900 2360
rect 57379 2329 57391 2332
rect 57333 2323 57391 2329
rect 58894 2320 58900 2332
rect 58952 2320 58958 2372
rect 35492 2264 38424 2292
rect 35492 2252 35498 2264
rect 43530 2252 43536 2304
rect 43588 2292 43594 2304
rect 47121 2295 47179 2301
rect 47121 2292 47133 2295
rect 43588 2264 47133 2292
rect 43588 2252 43594 2264
rect 47121 2261 47133 2264
rect 47167 2261 47179 2295
rect 47121 2255 47179 2261
rect 47210 2252 47216 2304
rect 47268 2292 47274 2304
rect 50525 2295 50583 2301
rect 50525 2292 50537 2295
rect 47268 2264 50537 2292
rect 47268 2252 47274 2264
rect 50525 2261 50537 2264
rect 50571 2261 50583 2295
rect 50525 2255 50583 2261
rect 52454 2252 52460 2304
rect 52512 2292 52518 2304
rect 53101 2295 53159 2301
rect 53101 2292 53113 2295
rect 52512 2264 53113 2292
rect 52512 2252 52518 2264
rect 53101 2261 53113 2264
rect 53147 2261 53159 2295
rect 53101 2255 53159 2261
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 11146 2088 11152 2100
rect 7708 2060 11152 2088
rect 7708 2048 7714 2060
rect 11146 2048 11152 2060
rect 11204 2048 11210 2100
rect 12342 2048 12348 2100
rect 12400 2088 12406 2100
rect 15654 2088 15660 2100
rect 12400 2060 15660 2088
rect 12400 2048 12406 2060
rect 15654 2048 15660 2060
rect 15712 2048 15718 2100
rect 18230 2048 18236 2100
rect 18288 2088 18294 2100
rect 21634 2088 21640 2100
rect 18288 2060 21640 2088
rect 18288 2048 18294 2060
rect 21634 2048 21640 2060
rect 21692 2048 21698 2100
rect 23474 2048 23480 2100
rect 23532 2088 23538 2100
rect 40954 2088 40960 2100
rect 23532 2060 40960 2088
rect 23532 2048 23538 2060
rect 40954 2048 40960 2060
rect 41012 2048 41018 2100
rect 42426 2048 42432 2100
rect 42484 2088 42490 2100
rect 44082 2088 44088 2100
rect 42484 2060 44088 2088
rect 42484 2048 42490 2060
rect 44082 2048 44088 2060
rect 44140 2048 44146 2100
rect 7742 1980 7748 2032
rect 7800 2020 7806 2032
rect 12710 2020 12716 2032
rect 7800 1992 12716 2020
rect 7800 1980 7806 1992
rect 12710 1980 12716 1992
rect 12768 1980 12774 2032
rect 14366 1980 14372 2032
rect 14424 2020 14430 2032
rect 23658 2020 23664 2032
rect 14424 1992 23664 2020
rect 14424 1980 14430 1992
rect 23658 1980 23664 1992
rect 23716 1980 23722 2032
rect 26970 1980 26976 2032
rect 27028 2020 27034 2032
rect 34882 2020 34888 2032
rect 27028 1992 34888 2020
rect 27028 1980 27034 1992
rect 34882 1980 34888 1992
rect 34940 1980 34946 2032
rect 42702 1980 42708 2032
rect 42760 2020 42766 2032
rect 47210 2020 47216 2032
rect 42760 1992 47216 2020
rect 42760 1980 42766 1992
rect 47210 1980 47216 1992
rect 47268 1980 47274 2032
rect 6914 1912 6920 1964
rect 6972 1952 6978 1964
rect 10594 1952 10600 1964
rect 6972 1924 10600 1952
rect 6972 1912 6978 1924
rect 10594 1912 10600 1924
rect 10652 1912 10658 1964
rect 17494 1912 17500 1964
rect 17552 1952 17558 1964
rect 23014 1952 23020 1964
rect 17552 1924 23020 1952
rect 17552 1912 17558 1924
rect 23014 1912 23020 1924
rect 23072 1912 23078 1964
rect 9122 1844 9128 1896
rect 9180 1884 9186 1896
rect 27614 1884 27620 1896
rect 9180 1856 27620 1884
rect 9180 1844 9186 1856
rect 27614 1844 27620 1856
rect 27672 1844 27678 1896
rect 1578 1776 1584 1828
rect 1636 1816 1642 1828
rect 26786 1816 26792 1828
rect 1636 1788 26792 1816
rect 1636 1776 1642 1788
rect 26786 1776 26792 1788
rect 26844 1776 26850 1828
rect 7098 1708 7104 1760
rect 7156 1748 7162 1760
rect 12802 1748 12808 1760
rect 7156 1720 12808 1748
rect 7156 1708 7162 1720
rect 12802 1708 12808 1720
rect 12860 1708 12866 1760
rect 5350 1640 5356 1692
rect 5408 1680 5414 1692
rect 9398 1680 9404 1692
rect 5408 1652 9404 1680
rect 5408 1640 5414 1652
rect 9398 1640 9404 1652
rect 9456 1640 9462 1692
rect 10134 1640 10140 1692
rect 10192 1680 10198 1692
rect 11422 1680 11428 1692
rect 10192 1652 11428 1680
rect 10192 1640 10198 1652
rect 11422 1640 11428 1652
rect 11480 1640 11486 1692
rect 5810 1572 5816 1624
rect 5868 1612 5874 1624
rect 10042 1612 10048 1624
rect 5868 1584 10048 1612
rect 5868 1572 5874 1584
rect 10042 1572 10048 1584
rect 10100 1572 10106 1624
rect 14918 1300 14924 1352
rect 14976 1340 14982 1352
rect 37550 1340 37556 1352
rect 14976 1312 37556 1340
rect 14976 1300 14982 1312
rect 37550 1300 37556 1312
rect 37608 1300 37614 1352
rect 38746 1300 38752 1352
rect 38804 1340 38810 1352
rect 56502 1340 56508 1352
rect 38804 1312 56508 1340
rect 38804 1300 38810 1312
rect 56502 1300 56508 1312
rect 56560 1300 56566 1352
rect 39850 1232 39856 1284
rect 39908 1272 39914 1284
rect 43806 1272 43812 1284
rect 39908 1244 43812 1272
rect 39908 1232 39914 1244
rect 43806 1232 43812 1244
rect 43864 1232 43870 1284
rect 18138 1164 18144 1216
rect 18196 1204 18202 1216
rect 21358 1204 21364 1216
rect 18196 1176 21364 1204
rect 18196 1164 18202 1176
rect 21358 1164 21364 1176
rect 21416 1164 21422 1216
rect 32398 1164 32404 1216
rect 32456 1204 32462 1216
rect 36078 1204 36084 1216
rect 32456 1176 36084 1204
rect 32456 1164 32462 1176
rect 36078 1164 36084 1176
rect 36136 1164 36142 1216
rect 38746 1164 38752 1216
rect 38804 1204 38810 1216
rect 39206 1204 39212 1216
rect 38804 1176 39212 1204
rect 38804 1164 38810 1176
rect 39206 1164 39212 1176
rect 39264 1164 39270 1216
rect 40954 1164 40960 1216
rect 41012 1204 41018 1216
rect 45002 1204 45008 1216
rect 41012 1176 45008 1204
rect 41012 1164 41018 1176
rect 45002 1164 45008 1176
rect 45060 1164 45066 1216
rect 13446 1096 13452 1148
rect 13504 1136 13510 1148
rect 14458 1136 14464 1148
rect 13504 1108 14464 1136
rect 13504 1096 13510 1108
rect 14458 1096 14464 1108
rect 14516 1096 14522 1148
rect 17586 1096 17592 1148
rect 17644 1136 17650 1148
rect 20530 1136 20536 1148
rect 17644 1108 20536 1136
rect 17644 1096 17650 1108
rect 20530 1096 20536 1108
rect 20588 1096 20594 1148
rect 27798 1096 27804 1148
rect 27856 1136 27862 1148
rect 29086 1136 29092 1148
rect 27856 1108 29092 1136
rect 27856 1096 27862 1108
rect 29086 1096 29092 1108
rect 29144 1096 29150 1148
rect 33778 1096 33784 1148
rect 33836 1136 33842 1148
rect 36538 1136 36544 1148
rect 33836 1108 36544 1136
rect 33836 1096 33842 1108
rect 36538 1096 36544 1108
rect 36596 1096 36602 1148
rect 43438 1096 43444 1148
rect 43496 1136 43502 1148
rect 46106 1136 46112 1148
rect 43496 1108 46112 1136
rect 43496 1096 43502 1108
rect 46106 1096 46112 1108
rect 46164 1096 46170 1148
rect 12618 1028 12624 1080
rect 12676 1068 12682 1080
rect 14182 1068 14188 1080
rect 12676 1040 14188 1068
rect 12676 1028 12682 1040
rect 14182 1028 14188 1040
rect 14240 1028 14246 1080
rect 18966 1028 18972 1080
rect 19024 1068 19030 1080
rect 21910 1068 21916 1080
rect 19024 1040 21916 1068
rect 19024 1028 19030 1040
rect 21910 1028 21916 1040
rect 21968 1028 21974 1080
rect 27338 1028 27344 1080
rect 27396 1068 27402 1080
rect 28534 1068 28540 1080
rect 27396 1040 28540 1068
rect 27396 1028 27402 1040
rect 28534 1028 28540 1040
rect 28592 1028 28598 1080
rect 32122 1028 32128 1080
rect 32180 1068 32186 1080
rect 35158 1068 35164 1080
rect 32180 1040 35164 1068
rect 32180 1028 32186 1040
rect 35158 1028 35164 1040
rect 35216 1028 35222 1080
rect 42610 1028 42616 1080
rect 42668 1068 42674 1080
rect 44726 1068 44732 1080
rect 42668 1040 44732 1068
rect 42668 1028 42674 1040
rect 44726 1028 44732 1040
rect 44784 1028 44790 1080
rect 5074 960 5080 1012
rect 5132 1000 5138 1012
rect 6730 1000 6736 1012
rect 5132 972 6736 1000
rect 5132 960 5138 972
rect 6730 960 6736 972
rect 6788 960 6794 1012
rect 11054 960 11060 1012
rect 11112 1000 11118 1012
rect 12802 1000 12808 1012
rect 11112 972 12808 1000
rect 11112 960 11118 972
rect 12802 960 12808 972
rect 12860 960 12866 1012
rect 14274 960 14280 1012
rect 14332 1000 14338 1012
rect 15562 1000 15568 1012
rect 14332 972 15568 1000
rect 14332 960 14338 972
rect 15562 960 15568 972
rect 15620 960 15626 1012
rect 16298 960 16304 1012
rect 16356 1000 16362 1012
rect 16356 972 19196 1000
rect 16356 960 16362 972
rect 3234 892 3240 944
rect 3292 932 3298 944
rect 4522 932 4528 944
rect 3292 904 4528 932
rect 3292 892 3298 904
rect 4522 892 4528 904
rect 4580 892 4586 944
rect 5166 892 5172 944
rect 5224 932 5230 944
rect 6178 932 6184 944
rect 5224 904 6184 932
rect 5224 892 5230 904
rect 6178 892 6184 904
rect 6236 892 6242 944
rect 6914 892 6920 944
rect 6972 932 6978 944
rect 9490 932 9496 944
rect 6972 904 9496 932
rect 6972 892 6978 904
rect 9490 892 9496 904
rect 9548 892 9554 944
rect 13722 892 13728 944
rect 13780 932 13786 944
rect 14734 932 14740 944
rect 13780 904 14740 932
rect 13780 892 13786 904
rect 14734 892 14740 904
rect 14792 892 14798 944
rect 17310 892 17316 944
rect 17368 932 17374 944
rect 18322 932 18328 944
rect 17368 904 18328 932
rect 17368 892 17374 904
rect 18322 892 18328 904
rect 18380 892 18386 944
rect 19168 932 19196 972
rect 19242 960 19248 1012
rect 19300 1000 19306 1012
rect 20806 1000 20812 1012
rect 19300 972 20812 1000
rect 19300 960 19306 972
rect 20806 960 20812 972
rect 20864 960 20870 1012
rect 22002 960 22008 1012
rect 22060 1000 22066 1012
rect 23014 1000 23020 1012
rect 22060 972 23020 1000
rect 22060 960 22066 972
rect 23014 960 23020 972
rect 23072 960 23078 1012
rect 23198 960 23204 1012
rect 23256 1000 23262 1012
rect 24394 1000 24400 1012
rect 23256 972 24400 1000
rect 23256 960 23262 972
rect 24394 960 24400 972
rect 24452 960 24458 1012
rect 26418 960 26424 1012
rect 26476 1000 26482 1012
rect 28810 1000 28816 1012
rect 26476 972 28816 1000
rect 26476 960 26482 972
rect 28810 960 28816 972
rect 28868 960 28874 1012
rect 31846 960 31852 1012
rect 31904 1000 31910 1012
rect 33502 1000 33508 1012
rect 31904 972 33508 1000
rect 31904 960 31910 972
rect 33502 960 33508 972
rect 33560 960 33566 1012
rect 35618 1000 35624 1012
rect 33612 972 35624 1000
rect 19426 932 19432 944
rect 19168 904 19432 932
rect 19426 892 19432 904
rect 19484 892 19490 944
rect 20714 892 20720 944
rect 20772 932 20778 944
rect 22186 932 22192 944
rect 20772 904 22192 932
rect 20772 892 20778 904
rect 22186 892 22192 904
rect 22244 892 22250 944
rect 23382 892 23388 944
rect 23440 932 23446 944
rect 24118 932 24124 944
rect 23440 904 24124 932
rect 23440 892 23446 904
rect 24118 892 24124 904
rect 24176 892 24182 944
rect 27522 892 27528 944
rect 27580 932 27586 944
rect 28258 932 28264 944
rect 27580 904 28264 932
rect 27580 892 27586 904
rect 28258 892 28264 904
rect 28316 892 28322 944
rect 28902 892 28908 944
rect 28960 932 28966 944
rect 29362 932 29368 944
rect 28960 904 29368 932
rect 28960 892 28966 904
rect 29362 892 29368 904
rect 29420 892 29426 944
rect 31294 892 31300 944
rect 31352 932 31358 944
rect 32582 932 32588 944
rect 31352 904 32588 932
rect 31352 892 31358 904
rect 32582 892 32588 904
rect 32640 892 32646 944
rect 32950 892 32956 944
rect 33008 932 33014 944
rect 33612 932 33640 972
rect 35618 960 35624 972
rect 35676 960 35682 1012
rect 40678 960 40684 1012
rect 40736 1000 40742 1012
rect 45278 1000 45284 1012
rect 40736 972 45284 1000
rect 40736 960 40742 972
rect 45278 960 45284 972
rect 45336 960 45342 1012
rect 47302 960 47308 1012
rect 47360 1000 47366 1012
rect 48774 1000 48780 1012
rect 47360 972 48780 1000
rect 47360 960 47366 972
rect 48774 960 48780 972
rect 48832 960 48838 1012
rect 50062 960 50068 1012
rect 50120 1000 50126 1012
rect 51902 1000 51908 1012
rect 50120 972 51908 1000
rect 50120 960 50126 972
rect 51902 960 51908 972
rect 51960 960 51966 1012
rect 33008 904 33640 932
rect 33008 892 33014 904
rect 34054 892 34060 944
rect 34112 932 34118 944
rect 37734 932 37740 944
rect 34112 904 37740 932
rect 34112 892 34118 904
rect 37734 892 37740 904
rect 37792 892 37798 944
rect 39574 892 39580 944
rect 39632 932 39638 944
rect 41046 932 41052 944
rect 39632 904 41052 932
rect 39632 892 39638 904
rect 41046 892 41052 904
rect 41104 892 41110 944
rect 42334 892 42340 944
rect 42392 932 42398 944
rect 46290 932 46296 944
rect 42392 904 46296 932
rect 42392 892 42398 904
rect 46290 892 46296 904
rect 46348 892 46354 944
rect 46474 892 46480 944
rect 46532 932 46538 944
rect 47394 932 47400 944
rect 46532 904 47400 932
rect 46532 892 46538 904
rect 47394 892 47400 904
rect 47452 892 47458 944
rect 49234 892 49240 944
rect 49292 932 49298 944
rect 51074 932 51080 944
rect 49292 904 51080 932
rect 49292 892 49298 904
rect 51074 892 51080 904
rect 51132 892 51138 944
rect 47946 824 47952 876
rect 48004 864 48010 876
rect 49694 864 49700 876
rect 48004 836 49700 864
rect 48004 824 48010 836
rect 49694 824 49700 836
rect 49752 824 49758 876
rect 35250 348 35256 400
rect 35308 388 35314 400
rect 38930 388 38936 400
rect 35308 360 38936 388
rect 35308 348 35314 360
rect 38930 348 38936 360
rect 38988 348 38994 400
rect 34974 144 34980 196
rect 35032 184 35038 196
rect 38654 184 38660 196
rect 35032 156 38660 184
rect 35032 144 35038 156
rect 38654 144 38660 156
rect 38712 144 38718 196
rect 35526 76 35532 128
rect 35584 116 35590 128
rect 38838 116 38844 128
rect 35584 88 38844 116
rect 35584 76 35590 88
rect 38838 76 38844 88
rect 38896 76 38902 128
<< via1 >>
rect 30196 63248 30248 63300
rect 30472 63248 30524 63300
rect 32588 63248 32640 63300
rect 33324 63248 33376 63300
rect 34060 63248 34112 63300
rect 34796 63248 34848 63300
rect 39212 63248 39264 63300
rect 40132 63248 40184 63300
rect 40684 63248 40736 63300
rect 41604 63248 41656 63300
rect 43536 63112 43588 63164
rect 44364 63112 44416 63164
rect 30288 61684 30340 61736
rect 49424 61684 49476 61736
rect 9772 61616 9824 61668
rect 23480 61616 23532 61668
rect 33508 61616 33560 61668
rect 41788 61616 41840 61668
rect 5172 61548 5224 61600
rect 17868 61548 17920 61600
rect 28908 61548 28960 61600
rect 46848 61548 46900 61600
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 5172 61387 5224 61396
rect 5172 61353 5181 61387
rect 5181 61353 5215 61387
rect 5215 61353 5224 61387
rect 5172 61344 5224 61353
rect 8208 61344 8260 61396
rect 35992 61344 36044 61396
rect 36176 61344 36228 61396
rect 46848 61387 46900 61396
rect 46848 61353 46857 61387
rect 46857 61353 46891 61387
rect 46891 61353 46900 61387
rect 46848 61344 46900 61353
rect 49424 61387 49476 61396
rect 49424 61353 49433 61387
rect 49433 61353 49467 61387
rect 49467 61353 49476 61387
rect 49424 61344 49476 61353
rect 9772 61276 9824 61328
rect 19340 61276 19392 61328
rect 22100 61276 22152 61328
rect 26884 61276 26936 61328
rect 7656 61208 7708 61260
rect 18052 61208 18104 61260
rect 23020 61208 23072 61260
rect 940 61140 992 61192
rect 1032 61072 1084 61124
rect 4620 61140 4672 61192
rect 5080 61183 5132 61192
rect 5080 61149 5089 61183
rect 5089 61149 5123 61183
rect 5123 61149 5132 61183
rect 5080 61140 5132 61149
rect 5724 61183 5776 61192
rect 5724 61149 5733 61183
rect 5733 61149 5767 61183
rect 5767 61149 5776 61183
rect 5724 61140 5776 61149
rect 6644 61183 6696 61192
rect 6644 61149 6653 61183
rect 6653 61149 6687 61183
rect 6687 61149 6696 61183
rect 6644 61140 6696 61149
rect 7564 61183 7616 61192
rect 7564 61149 7573 61183
rect 7573 61149 7607 61183
rect 7607 61149 7616 61183
rect 7564 61140 7616 61149
rect 9680 61140 9732 61192
rect 10232 61183 10284 61192
rect 10232 61149 10241 61183
rect 10241 61149 10275 61183
rect 10275 61149 10284 61183
rect 10232 61140 10284 61149
rect 11152 61140 11204 61192
rect 11980 61183 12032 61192
rect 11980 61149 11989 61183
rect 11989 61149 12023 61183
rect 12023 61149 12032 61183
rect 11980 61140 12032 61149
rect 12716 61183 12768 61192
rect 12716 61149 12725 61183
rect 12725 61149 12759 61183
rect 12759 61149 12768 61183
rect 12716 61140 12768 61149
rect 14924 61183 14976 61192
rect 14924 61149 14933 61183
rect 14933 61149 14967 61183
rect 14967 61149 14976 61183
rect 14924 61140 14976 61149
rect 16120 61183 16172 61192
rect 16120 61149 16129 61183
rect 16129 61149 16163 61183
rect 16163 61149 16172 61183
rect 16120 61140 16172 61149
rect 17132 61183 17184 61192
rect 17132 61149 17141 61183
rect 17141 61149 17175 61183
rect 17175 61149 17184 61183
rect 17132 61140 17184 61149
rect 17960 61183 18012 61192
rect 17960 61149 17969 61183
rect 17969 61149 18003 61183
rect 18003 61149 18012 61183
rect 17960 61140 18012 61149
rect 18696 61183 18748 61192
rect 18696 61149 18705 61183
rect 18705 61149 18739 61183
rect 18739 61149 18748 61183
rect 18696 61140 18748 61149
rect 19800 61183 19852 61192
rect 19800 61149 19809 61183
rect 19809 61149 19843 61183
rect 19843 61149 19852 61183
rect 19800 61140 19852 61149
rect 20720 61140 20772 61192
rect 21272 61183 21324 61192
rect 21272 61149 21281 61183
rect 21281 61149 21315 61183
rect 21315 61149 21324 61183
rect 21272 61140 21324 61149
rect 22192 61140 22244 61192
rect 5632 61072 5684 61124
rect 6184 61072 6236 61124
rect 6920 61115 6972 61124
rect 6920 61081 6929 61115
rect 6929 61081 6963 61115
rect 6963 61081 6972 61115
rect 6920 61072 6972 61081
rect 9128 61072 9180 61124
rect 13636 61072 13688 61124
rect 15200 61115 15252 61124
rect 15200 61081 15209 61115
rect 15209 61081 15243 61115
rect 15243 61081 15252 61115
rect 15200 61072 15252 61081
rect 17500 61072 17552 61124
rect 19984 61115 20036 61124
rect 19984 61081 19993 61115
rect 19993 61081 20027 61115
rect 20027 61081 20036 61115
rect 19984 61072 20036 61081
rect 21180 61072 21232 61124
rect 32956 61208 33008 61260
rect 35900 61208 35952 61260
rect 23664 61140 23716 61192
rect 25136 61140 25188 61192
rect 26240 61183 26292 61192
rect 26240 61149 26249 61183
rect 26249 61149 26283 61183
rect 26283 61149 26292 61183
rect 26240 61140 26292 61149
rect 26608 61140 26660 61192
rect 28080 61140 28132 61192
rect 29828 61183 29880 61192
rect 29828 61149 29837 61183
rect 29837 61149 29871 61183
rect 29871 61149 29880 61183
rect 29828 61140 29880 61149
rect 31208 61183 31260 61192
rect 31208 61149 31217 61183
rect 31217 61149 31251 61183
rect 31251 61149 31260 61183
rect 31208 61140 31260 61149
rect 31760 61140 31812 61192
rect 33324 61183 33376 61192
rect 33324 61149 33333 61183
rect 33333 61149 33367 61183
rect 33367 61149 33376 61183
rect 33324 61140 33376 61149
rect 33508 61183 33560 61192
rect 33508 61149 33517 61183
rect 33517 61149 33551 61183
rect 33551 61149 33560 61183
rect 33508 61140 33560 61149
rect 34796 61140 34848 61192
rect 24768 61072 24820 61124
rect 28172 61072 28224 61124
rect 33232 61072 33284 61124
rect 34704 61072 34756 61124
rect 35900 61115 35952 61124
rect 35900 61081 35909 61115
rect 35909 61081 35943 61115
rect 35943 61081 35952 61115
rect 35900 61072 35952 61081
rect 35992 61072 36044 61124
rect 37280 61140 37332 61192
rect 37648 61140 37700 61192
rect 38752 61140 38804 61192
rect 40132 61183 40184 61192
rect 40132 61149 40141 61183
rect 40141 61149 40175 61183
rect 40175 61149 40184 61183
rect 40132 61140 40184 61149
rect 41604 61183 41656 61192
rect 41604 61149 41613 61183
rect 41613 61149 41647 61183
rect 41647 61149 41656 61183
rect 41604 61140 41656 61149
rect 42064 61140 42116 61192
rect 42800 61140 42852 61192
rect 38200 61072 38252 61124
rect 40040 61072 40092 61124
rect 41420 61072 41472 61124
rect 5908 61047 5960 61056
rect 5908 61013 5917 61047
rect 5917 61013 5951 61047
rect 5951 61013 5960 61047
rect 5908 61004 5960 61013
rect 12164 61047 12216 61056
rect 12164 61013 12173 61047
rect 12173 61013 12207 61047
rect 12207 61013 12216 61047
rect 12164 61004 12216 61013
rect 17316 61047 17368 61056
rect 17316 61013 17325 61047
rect 17325 61013 17359 61047
rect 17359 61013 17368 61047
rect 17316 61004 17368 61013
rect 18788 61047 18840 61056
rect 18788 61013 18797 61047
rect 18797 61013 18831 61047
rect 18831 61013 18840 61047
rect 18788 61004 18840 61013
rect 20996 61004 21048 61056
rect 22008 61004 22060 61056
rect 24676 61004 24728 61056
rect 25412 61047 25464 61056
rect 25412 61013 25421 61047
rect 25421 61013 25455 61047
rect 25455 61013 25464 61047
rect 25412 61004 25464 61013
rect 27344 61047 27396 61056
rect 27344 61013 27353 61047
rect 27353 61013 27387 61047
rect 27387 61013 27396 61047
rect 27344 61004 27396 61013
rect 28448 61004 28500 61056
rect 29920 61047 29972 61056
rect 29920 61013 29929 61047
rect 29929 61013 29963 61047
rect 29963 61013 29972 61047
rect 29920 61004 29972 61013
rect 31300 61047 31352 61056
rect 31300 61013 31309 61047
rect 31309 61013 31343 61047
rect 31343 61013 31352 61047
rect 31300 61004 31352 61013
rect 32588 61004 32640 61056
rect 33508 61004 33560 61056
rect 36084 61004 36136 61056
rect 39120 61047 39172 61056
rect 39120 61013 39129 61047
rect 39129 61013 39163 61047
rect 39163 61013 39172 61047
rect 39120 61004 39172 61013
rect 40224 61047 40276 61056
rect 40224 61013 40233 61047
rect 40233 61013 40267 61047
rect 40267 61013 40276 61047
rect 40224 61004 40276 61013
rect 40316 61004 40368 61056
rect 41696 61047 41748 61056
rect 41696 61013 41705 61047
rect 41705 61013 41739 61047
rect 41739 61013 41748 61047
rect 41696 61004 41748 61013
rect 42984 61072 43036 61124
rect 56692 61208 56744 61260
rect 58992 61208 59044 61260
rect 44364 61183 44416 61192
rect 44364 61149 44373 61183
rect 44373 61149 44407 61183
rect 44407 61149 44416 61183
rect 44364 61140 44416 61149
rect 44548 61140 44600 61192
rect 45560 61140 45612 61192
rect 44824 61072 44876 61124
rect 45744 61140 45796 61192
rect 47216 61140 47268 61192
rect 48320 61140 48372 61192
rect 48688 61140 48740 61192
rect 49792 61140 49844 61192
rect 51264 61140 51316 61192
rect 51632 61140 51684 61192
rect 53196 61183 53248 61192
rect 53196 61149 53205 61183
rect 53205 61149 53239 61183
rect 53239 61149 53248 61183
rect 53196 61140 53248 61149
rect 54116 61183 54168 61192
rect 54116 61149 54125 61183
rect 54125 61149 54159 61183
rect 54159 61149 54168 61183
rect 54116 61140 54168 61149
rect 55496 61183 55548 61192
rect 55496 61149 55505 61183
rect 55505 61149 55539 61183
rect 55539 61149 55548 61183
rect 55496 61140 55548 61149
rect 56048 61140 56100 61192
rect 57520 61140 57572 61192
rect 45376 61047 45428 61056
rect 45376 61013 45385 61047
rect 45385 61013 45419 61047
rect 45419 61013 45428 61047
rect 45376 61004 45428 61013
rect 49700 61072 49752 61124
rect 53472 61115 53524 61124
rect 53472 61081 53481 61115
rect 53481 61081 53515 61115
rect 53515 61081 53524 61115
rect 53472 61072 53524 61081
rect 55772 61115 55824 61124
rect 55772 61081 55781 61115
rect 55781 61081 55815 61115
rect 55815 61081 55824 61115
rect 55772 61072 55824 61081
rect 58348 61115 58400 61124
rect 58348 61081 58357 61115
rect 58357 61081 58391 61115
rect 58391 61081 58400 61115
rect 58348 61072 58400 61081
rect 46848 61004 46900 61056
rect 50068 61004 50120 61056
rect 50620 61004 50672 61056
rect 54300 61047 54352 61056
rect 54300 61013 54309 61047
rect 54309 61013 54343 61047
rect 54343 61013 54352 61047
rect 54300 61004 54352 61013
rect 56600 61047 56652 61056
rect 56600 61013 56609 61047
rect 56609 61013 56643 61047
rect 56643 61013 56652 61047
rect 56600 61004 56652 61013
rect 19574 60902 19626 60954
rect 19638 60902 19690 60954
rect 19702 60902 19754 60954
rect 19766 60902 19818 60954
rect 19830 60902 19882 60954
rect 50294 60902 50346 60954
rect 50358 60902 50410 60954
rect 50422 60902 50474 60954
rect 50486 60902 50538 60954
rect 50550 60902 50602 60954
rect 3240 60775 3292 60784
rect 3240 60741 3249 60775
rect 3249 60741 3283 60775
rect 3283 60741 3292 60775
rect 3240 60732 3292 60741
rect 3976 60775 4028 60784
rect 3976 60741 3985 60775
rect 3985 60741 4019 60775
rect 4019 60741 4028 60775
rect 3976 60732 4028 60741
rect 8392 60775 8444 60784
rect 8392 60741 8401 60775
rect 8401 60741 8435 60775
rect 8435 60741 8444 60775
rect 8392 60732 8444 60741
rect 13544 60775 13596 60784
rect 13544 60741 13553 60775
rect 13553 60741 13587 60775
rect 13587 60741 13596 60775
rect 13544 60732 13596 60741
rect 14280 60775 14332 60784
rect 14280 60741 14289 60775
rect 14289 60741 14323 60775
rect 14323 60741 14332 60775
rect 14280 60732 14332 60741
rect 15752 60775 15804 60784
rect 15752 60741 15761 60775
rect 15761 60741 15795 60775
rect 15795 60741 15804 60775
rect 15752 60732 15804 60741
rect 19432 60775 19484 60784
rect 19432 60741 19441 60775
rect 19441 60741 19475 60775
rect 19475 60741 19484 60775
rect 19432 60732 19484 60741
rect 22192 60732 22244 60784
rect 36176 60800 36228 60852
rect 24400 60732 24452 60784
rect 24676 60732 24728 60784
rect 40224 60800 40276 60852
rect 36360 60775 36412 60784
rect 36360 60741 36369 60775
rect 36369 60741 36403 60775
rect 36403 60741 36412 60775
rect 36360 60732 36412 60741
rect 41512 60775 41564 60784
rect 41512 60741 41521 60775
rect 41521 60741 41555 60775
rect 41555 60741 41564 60775
rect 41512 60732 41564 60741
rect 46664 60775 46716 60784
rect 46664 60741 46673 60775
rect 46673 60741 46707 60775
rect 46707 60741 46716 60775
rect 46664 60732 46716 60741
rect 50160 60732 50212 60784
rect 52644 60732 52696 60784
rect 940 60664 992 60716
rect 9036 60707 9088 60716
rect 9036 60673 9045 60707
rect 9045 60673 9079 60707
rect 9079 60673 9088 60707
rect 9036 60664 9088 60673
rect 17868 60664 17920 60716
rect 7932 60596 7984 60648
rect 18420 60596 18472 60648
rect 19616 60596 19668 60648
rect 22192 60596 22244 60648
rect 23664 60664 23716 60716
rect 27528 60707 27580 60716
rect 27528 60673 27537 60707
rect 27537 60673 27571 60707
rect 27571 60673 27580 60707
rect 27528 60664 27580 60673
rect 29000 60707 29052 60716
rect 29000 60673 29009 60707
rect 29009 60673 29043 60707
rect 29043 60673 29052 60707
rect 29000 60664 29052 60673
rect 30472 60707 30524 60716
rect 30472 60673 30481 60707
rect 30481 60673 30515 60707
rect 30515 60673 30524 60707
rect 30472 60664 30524 60673
rect 30564 60664 30616 60716
rect 4620 60528 4672 60580
rect 31208 60596 31260 60648
rect 54668 60707 54720 60716
rect 54668 60673 54677 60707
rect 54677 60673 54711 60707
rect 54711 60673 54720 60707
rect 54668 60664 54720 60673
rect 58900 60800 58952 60852
rect 56784 60732 56836 60784
rect 58992 60732 59044 60784
rect 56876 60707 56928 60716
rect 56876 60673 56885 60707
rect 56885 60673 56919 60707
rect 56919 60673 56928 60707
rect 56876 60664 56928 60673
rect 58072 60707 58124 60716
rect 58072 60673 58081 60707
rect 58081 60673 58115 60707
rect 58115 60673 58124 60707
rect 58072 60664 58124 60673
rect 3332 60503 3384 60512
rect 3332 60469 3341 60503
rect 3341 60469 3375 60503
rect 3375 60469 3384 60503
rect 3332 60460 3384 60469
rect 9220 60503 9272 60512
rect 9220 60469 9229 60503
rect 9229 60469 9263 60503
rect 9263 60469 9272 60503
rect 9220 60460 9272 60469
rect 15108 60460 15160 60512
rect 17868 60460 17920 60512
rect 20076 60460 20128 60512
rect 22284 60460 22336 60512
rect 24400 60460 24452 60512
rect 24676 60503 24728 60512
rect 24676 60469 24685 60503
rect 24685 60469 24719 60503
rect 24719 60469 24728 60503
rect 24676 60460 24728 60469
rect 24860 60460 24912 60512
rect 29000 60460 29052 60512
rect 29828 60460 29880 60512
rect 30012 60503 30064 60512
rect 30012 60469 30021 60503
rect 30021 60469 30055 60503
rect 30055 60469 30064 60503
rect 30012 60460 30064 60469
rect 42248 60528 42300 60580
rect 56692 60596 56744 60648
rect 58164 60528 58216 60580
rect 30932 60460 30984 60512
rect 35716 60460 35768 60512
rect 40960 60460 41012 60512
rect 44180 60460 44232 60512
rect 50436 60503 50488 60512
rect 50436 60469 50445 60503
rect 50445 60469 50479 60503
rect 50479 60469 50488 60503
rect 50436 60460 50488 60469
rect 53104 60503 53156 60512
rect 53104 60469 53113 60503
rect 53113 60469 53147 60503
rect 53147 60469 53156 60503
rect 53104 60460 53156 60469
rect 54852 60503 54904 60512
rect 54852 60469 54861 60503
rect 54861 60469 54895 60503
rect 54895 60469 54904 60503
rect 54852 60460 54904 60469
rect 55588 60503 55640 60512
rect 55588 60469 55597 60503
rect 55597 60469 55631 60503
rect 55631 60469 55640 60503
rect 55588 60460 55640 60469
rect 56324 60503 56376 60512
rect 56324 60469 56333 60503
rect 56333 60469 56367 60503
rect 56367 60469 56376 60503
rect 56324 60460 56376 60469
rect 57060 60503 57112 60512
rect 57060 60469 57069 60503
rect 57069 60469 57103 60503
rect 57103 60469 57112 60503
rect 57060 60460 57112 60469
rect 58256 60503 58308 60512
rect 58256 60469 58265 60503
rect 58265 60469 58299 60503
rect 58299 60469 58308 60503
rect 58256 60460 58308 60469
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 3332 60256 3384 60308
rect 20260 60256 20312 60308
rect 15108 60188 15160 60240
rect 19248 60188 19300 60240
rect 20168 60188 20220 60240
rect 21916 60188 21968 60240
rect 17868 60163 17920 60172
rect 17868 60129 17877 60163
rect 17877 60129 17911 60163
rect 17911 60129 17920 60163
rect 17868 60120 17920 60129
rect 18144 60120 18196 60172
rect 2596 60095 2648 60104
rect 2596 60061 2605 60095
rect 2605 60061 2639 60095
rect 2639 60061 2648 60095
rect 2596 60052 2648 60061
rect 5632 60052 5684 60104
rect 7748 60095 7800 60104
rect 7748 60061 7757 60095
rect 7757 60061 7791 60095
rect 7791 60061 7800 60095
rect 7748 60052 7800 60061
rect 940 59984 992 60036
rect 2044 60027 2096 60036
rect 2044 59993 2053 60027
rect 2053 59993 2087 60027
rect 2087 59993 2096 60027
rect 2044 59984 2096 59993
rect 7564 60027 7616 60036
rect 7564 59993 7573 60027
rect 7573 59993 7607 60027
rect 7607 59993 7616 60027
rect 7564 59984 7616 59993
rect 8208 59984 8260 60036
rect 2504 59916 2556 59968
rect 8024 59916 8076 59968
rect 17592 59916 17644 59968
rect 18420 60095 18472 60104
rect 18420 60061 18429 60095
rect 18429 60061 18463 60095
rect 18463 60061 18472 60095
rect 18420 60052 18472 60061
rect 18512 60052 18564 60104
rect 19616 60095 19668 60104
rect 19156 59984 19208 60036
rect 19616 60061 19625 60095
rect 19625 60061 19659 60095
rect 19659 60061 19668 60095
rect 19616 60052 19668 60061
rect 22008 60120 22060 60172
rect 19892 60095 19944 60104
rect 19892 60061 19895 60095
rect 19895 60061 19944 60095
rect 19892 60052 19944 60061
rect 19984 60052 20036 60104
rect 22284 60052 22336 60104
rect 58256 60256 58308 60308
rect 23296 60188 23348 60240
rect 30564 60188 30616 60240
rect 30748 60188 30800 60240
rect 41144 60188 41196 60240
rect 41236 60231 41288 60240
rect 41236 60197 41245 60231
rect 41245 60197 41279 60231
rect 41279 60197 41288 60231
rect 41236 60188 41288 60197
rect 41604 60188 41656 60240
rect 24860 60120 24912 60172
rect 22560 60095 22612 60104
rect 22560 60061 22569 60095
rect 22569 60061 22603 60095
rect 22603 60061 22612 60095
rect 22560 60052 22612 60061
rect 22836 60095 22888 60104
rect 22836 60061 22845 60095
rect 22845 60061 22879 60095
rect 22879 60061 22888 60095
rect 22836 60052 22888 60061
rect 23020 60095 23072 60104
rect 23020 60061 23029 60095
rect 23029 60061 23063 60095
rect 23063 60061 23072 60095
rect 23020 60052 23072 60061
rect 23204 60052 23256 60104
rect 29092 60120 29144 60172
rect 29184 60120 29236 60172
rect 28172 60095 28224 60104
rect 28172 60061 28182 60095
rect 28182 60061 28216 60095
rect 28216 60061 28224 60095
rect 28172 60052 28224 60061
rect 20812 60027 20864 60036
rect 20812 59993 20821 60027
rect 20821 59993 20855 60027
rect 20855 59993 20864 60027
rect 20812 59984 20864 59993
rect 20904 60027 20956 60036
rect 20904 59993 20913 60027
rect 20913 59993 20947 60027
rect 20947 59993 20956 60027
rect 20904 59984 20956 59993
rect 30196 60052 30248 60104
rect 30748 60095 30800 60104
rect 30748 60061 30757 60095
rect 30757 60061 30791 60095
rect 30791 60061 30800 60095
rect 30748 60052 30800 60061
rect 19892 59916 19944 59968
rect 19984 59916 20036 59968
rect 21272 59916 21324 59968
rect 21824 59959 21876 59968
rect 21824 59925 21833 59959
rect 21833 59925 21867 59959
rect 21867 59925 21876 59959
rect 21824 59916 21876 59925
rect 22284 59916 22336 59968
rect 23388 59916 23440 59968
rect 23664 59916 23716 59968
rect 23756 59916 23808 59968
rect 28908 59984 28960 60036
rect 30012 59984 30064 60036
rect 30932 60095 30984 60104
rect 30932 60061 30977 60095
rect 30977 60061 30984 60095
rect 30932 60052 30984 60061
rect 31116 60095 31168 60104
rect 31116 60061 31125 60095
rect 31125 60061 31159 60095
rect 31159 60061 31168 60095
rect 31116 60052 31168 60061
rect 31208 60052 31260 60104
rect 28632 59916 28684 59968
rect 28724 59959 28776 59968
rect 28724 59925 28733 59959
rect 28733 59925 28767 59959
rect 28767 59925 28776 59959
rect 28724 59916 28776 59925
rect 29092 59959 29144 59968
rect 29092 59925 29101 59959
rect 29101 59925 29135 59959
rect 29135 59925 29144 59959
rect 29092 59916 29144 59925
rect 30472 59959 30524 59968
rect 30472 59925 30481 59959
rect 30481 59925 30515 59959
rect 30515 59925 30524 59959
rect 30472 59916 30524 59925
rect 32220 59959 32272 59968
rect 32220 59925 32229 59959
rect 32229 59925 32263 59959
rect 32263 59925 32272 59959
rect 32220 59916 32272 59925
rect 32496 59916 32548 59968
rect 32956 60095 33008 60104
rect 32956 60061 32965 60095
rect 32965 60061 32999 60095
rect 32999 60061 33008 60095
rect 32956 60052 33008 60061
rect 34520 60052 34572 60104
rect 40960 60095 41012 60104
rect 40960 60061 40969 60095
rect 40969 60061 41003 60095
rect 41003 60061 41012 60095
rect 40960 60052 41012 60061
rect 41604 60052 41656 60104
rect 40868 60027 40920 60036
rect 40868 59993 40877 60027
rect 40877 59993 40911 60027
rect 40911 59993 40920 60027
rect 40868 59984 40920 59993
rect 42064 59984 42116 60036
rect 42248 60163 42300 60172
rect 42248 60129 42257 60163
rect 42257 60129 42291 60163
rect 42291 60129 42300 60163
rect 42248 60120 42300 60129
rect 42708 60163 42760 60172
rect 42708 60129 42717 60163
rect 42717 60129 42751 60163
rect 42751 60129 42760 60163
rect 42708 60120 42760 60129
rect 42432 60095 42484 60104
rect 42432 60061 42441 60095
rect 42441 60061 42475 60095
rect 42475 60061 42484 60095
rect 42432 60052 42484 60061
rect 50436 60120 50488 60172
rect 33048 59916 33100 59968
rect 42432 59916 42484 59968
rect 56232 60120 56284 60172
rect 56784 60052 56836 60104
rect 58992 60120 59044 60172
rect 57980 60052 58032 60104
rect 56692 60027 56744 60036
rect 56692 59993 56701 60027
rect 56701 59993 56735 60027
rect 56735 59993 56744 60027
rect 56692 59984 56744 59993
rect 59544 59984 59596 60036
rect 57336 59959 57388 59968
rect 57336 59925 57345 59959
rect 57345 59925 57379 59959
rect 57379 59925 57388 59959
rect 57336 59916 57388 59925
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 7748 59712 7800 59764
rect 19984 59712 20036 59764
rect 20904 59712 20956 59764
rect 55588 59712 55640 59764
rect 56232 59712 56284 59764
rect 58164 59712 58216 59764
rect 1584 59644 1636 59696
rect 7564 59644 7616 59696
rect 19156 59644 19208 59696
rect 21364 59644 21416 59696
rect 940 59576 992 59628
rect 18052 59576 18104 59628
rect 21180 59619 21232 59628
rect 21180 59585 21189 59619
rect 21189 59585 21223 59619
rect 21223 59585 21232 59619
rect 21180 59576 21232 59585
rect 21272 59619 21324 59628
rect 21272 59585 21281 59619
rect 21281 59585 21315 59619
rect 21315 59585 21324 59619
rect 21272 59576 21324 59585
rect 22100 59619 22152 59628
rect 22100 59585 22109 59619
rect 22109 59585 22143 59619
rect 22143 59585 22152 59619
rect 22100 59576 22152 59585
rect 20812 59508 20864 59560
rect 22836 59644 22888 59696
rect 29460 59644 29512 59696
rect 23296 59576 23348 59628
rect 23388 59619 23440 59628
rect 23388 59585 23397 59619
rect 23397 59585 23431 59619
rect 23431 59585 23440 59619
rect 23388 59576 23440 59585
rect 23480 59619 23532 59628
rect 23480 59585 23489 59619
rect 23489 59585 23523 59619
rect 23523 59585 23532 59619
rect 23480 59576 23532 59585
rect 23572 59619 23624 59628
rect 23572 59585 23586 59619
rect 23586 59585 23620 59619
rect 23620 59585 23624 59619
rect 23572 59576 23624 59585
rect 28356 59619 28408 59628
rect 28356 59585 28365 59619
rect 28365 59585 28399 59619
rect 28399 59585 28408 59619
rect 28356 59576 28408 59585
rect 28632 59619 28684 59628
rect 28632 59585 28641 59619
rect 28641 59585 28675 59619
rect 28675 59585 28684 59619
rect 30104 59687 30156 59696
rect 30104 59653 30113 59687
rect 30113 59653 30147 59687
rect 30147 59653 30156 59687
rect 30104 59644 30156 59653
rect 30288 59644 30340 59696
rect 28632 59576 28684 59585
rect 29736 59619 29788 59628
rect 29736 59585 29745 59619
rect 29745 59585 29779 59619
rect 29779 59585 29788 59619
rect 29736 59576 29788 59585
rect 29828 59619 29880 59628
rect 29828 59585 29838 59619
rect 29838 59585 29872 59619
rect 29872 59585 29880 59619
rect 29828 59576 29880 59585
rect 30012 59619 30064 59628
rect 30012 59585 30021 59619
rect 30021 59585 30055 59619
rect 30055 59585 30064 59619
rect 30012 59576 30064 59585
rect 30196 59619 30248 59628
rect 30196 59585 30210 59619
rect 30210 59585 30244 59619
rect 30244 59585 30248 59619
rect 30196 59576 30248 59585
rect 34520 59576 34572 59628
rect 22560 59440 22612 59492
rect 23388 59440 23440 59492
rect 24860 59440 24912 59492
rect 29644 59508 29696 59560
rect 30288 59440 30340 59492
rect 30380 59483 30432 59492
rect 30380 59449 30389 59483
rect 30389 59449 30423 59483
rect 30423 59449 30432 59483
rect 30380 59440 30432 59449
rect 1952 59415 2004 59424
rect 1952 59381 1961 59415
rect 1961 59381 1995 59415
rect 1995 59381 2004 59415
rect 1952 59372 2004 59381
rect 2320 59372 2372 59424
rect 19248 59372 19300 59424
rect 22468 59372 22520 59424
rect 22928 59372 22980 59424
rect 24492 59372 24544 59424
rect 29736 59372 29788 59424
rect 30012 59372 30064 59424
rect 30656 59415 30708 59424
rect 30656 59381 30665 59415
rect 30665 59381 30699 59415
rect 30699 59381 30708 59415
rect 30656 59372 30708 59381
rect 40868 59440 40920 59492
rect 42432 59644 42484 59696
rect 41788 59576 41840 59628
rect 58808 59644 58860 59696
rect 53104 59576 53156 59628
rect 58072 59619 58124 59628
rect 58072 59585 58081 59619
rect 58081 59585 58115 59619
rect 58115 59585 58124 59619
rect 58072 59576 58124 59585
rect 42708 59551 42760 59560
rect 42708 59517 42717 59551
rect 42717 59517 42751 59551
rect 42751 59517 42760 59551
rect 42708 59508 42760 59517
rect 42800 59508 42852 59560
rect 56324 59508 56376 59560
rect 57152 59440 57204 59492
rect 58716 59440 58768 59492
rect 32496 59372 32548 59424
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 1952 59032 2004 59084
rect 848 58964 900 59016
rect 19524 59100 19576 59152
rect 38844 59100 38896 59152
rect 58348 59100 58400 59152
rect 41604 59032 41656 59084
rect 19708 59007 19760 59016
rect 19708 58973 19717 59007
rect 19717 58973 19751 59007
rect 19751 58973 19760 59007
rect 19708 58964 19760 58973
rect 21364 58964 21416 59016
rect 23572 58964 23624 59016
rect 41512 59007 41564 59016
rect 41512 58973 41521 59007
rect 41521 58973 41555 59007
rect 41555 58973 41564 59007
rect 41512 58964 41564 58973
rect 50620 59032 50672 59084
rect 57152 59007 57204 59016
rect 57152 58973 57161 59007
rect 57161 58973 57195 59007
rect 57195 58973 57204 59007
rect 57152 58964 57204 58973
rect 58992 58964 59044 59016
rect 18512 58828 18564 58880
rect 58900 58896 58952 58948
rect 20076 58828 20128 58880
rect 41144 58871 41196 58880
rect 41144 58837 41153 58871
rect 41153 58837 41187 58871
rect 41187 58837 41196 58871
rect 41144 58828 41196 58837
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 2044 58624 2096 58676
rect 940 58488 992 58540
rect 34520 58488 34572 58540
rect 37924 58531 37976 58540
rect 3424 58420 3476 58472
rect 35808 58420 35860 58472
rect 37924 58497 37933 58531
rect 37933 58497 37967 58531
rect 37967 58497 37976 58531
rect 37924 58488 37976 58497
rect 38200 58531 38252 58540
rect 38200 58497 38209 58531
rect 38209 58497 38243 58531
rect 38243 58497 38252 58531
rect 38200 58488 38252 58497
rect 38292 58531 38344 58540
rect 38292 58497 38301 58531
rect 38301 58497 38335 58531
rect 38335 58497 38344 58531
rect 38292 58488 38344 58497
rect 38476 58488 38528 58540
rect 38844 58531 38896 58540
rect 38844 58497 38853 58531
rect 38853 58497 38887 58531
rect 38887 58497 38896 58531
rect 38844 58488 38896 58497
rect 58164 58599 58216 58608
rect 58164 58565 58173 58599
rect 58173 58565 58207 58599
rect 58207 58565 58216 58599
rect 58164 58556 58216 58565
rect 40040 58420 40092 58472
rect 49700 58488 49752 58540
rect 36912 58352 36964 58404
rect 38292 58352 38344 58404
rect 37556 58327 37608 58336
rect 37556 58293 37565 58327
rect 37565 58293 37599 58327
rect 37599 58293 37608 58327
rect 37556 58284 37608 58293
rect 37924 58284 37976 58336
rect 41604 58352 41656 58404
rect 42616 58284 42668 58336
rect 58256 58327 58308 58336
rect 58256 58293 58265 58327
rect 58265 58293 58299 58327
rect 58299 58293 58308 58327
rect 58256 58284 58308 58293
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 940 57876 992 57928
rect 35808 57944 35860 57996
rect 35716 57919 35768 57928
rect 35716 57885 35725 57919
rect 35725 57885 35759 57919
rect 35759 57885 35768 57919
rect 35716 57876 35768 57885
rect 6000 57808 6052 57860
rect 34796 57808 34848 57860
rect 35440 57740 35492 57792
rect 36268 57919 36320 57928
rect 36268 57885 36277 57919
rect 36277 57885 36311 57919
rect 36311 57885 36320 57919
rect 36268 57876 36320 57885
rect 58256 57876 58308 57928
rect 57980 57851 58032 57860
rect 57980 57817 57989 57851
rect 57989 57817 58023 57851
rect 58023 57817 58032 57851
rect 57980 57808 58032 57817
rect 58072 57783 58124 57792
rect 58072 57749 58081 57783
rect 58081 57749 58115 57783
rect 58115 57749 58124 57783
rect 58072 57740 58124 57749
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 940 57400 992 57452
rect 1768 57239 1820 57248
rect 1768 57205 1777 57239
rect 1777 57205 1811 57239
rect 1811 57205 1820 57239
rect 1768 57196 1820 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 33416 56992 33468 57044
rect 24860 56924 24912 56976
rect 36268 56924 36320 56976
rect 41144 56992 41196 57044
rect 43260 56992 43312 57044
rect 56508 56924 56560 56976
rect 22468 56788 22520 56840
rect 33048 56831 33100 56840
rect 33048 56797 33057 56831
rect 33057 56797 33091 56831
rect 33091 56797 33100 56831
rect 33048 56788 33100 56797
rect 33416 56831 33468 56840
rect 33416 56797 33425 56831
rect 33425 56797 33459 56831
rect 33459 56797 33468 56831
rect 33416 56788 33468 56797
rect 58992 56788 59044 56840
rect 940 56720 992 56772
rect 41420 56720 41472 56772
rect 55864 56720 55916 56772
rect 32680 56695 32732 56704
rect 32680 56661 32689 56695
rect 32689 56661 32723 56695
rect 32723 56661 32732 56695
rect 32680 56652 32732 56661
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 56508 56448 56560 56500
rect 58992 56380 59044 56432
rect 41512 56355 41564 56364
rect 41512 56321 41521 56355
rect 41521 56321 41555 56355
rect 41555 56321 41564 56355
rect 41512 56312 41564 56321
rect 46848 56312 46900 56364
rect 41420 56287 41472 56296
rect 41420 56253 41429 56287
rect 41429 56253 41463 56287
rect 41463 56253 41472 56287
rect 41420 56244 41472 56253
rect 41236 56176 41288 56228
rect 41604 56176 41656 56228
rect 41328 56108 41380 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 23572 55904 23624 55956
rect 30472 55904 30524 55956
rect 58348 55947 58400 55956
rect 58348 55913 58357 55947
rect 58357 55913 58391 55947
rect 58391 55913 58400 55947
rect 58348 55904 58400 55913
rect 1768 55836 1820 55888
rect 24124 55768 24176 55820
rect 30564 55768 30616 55820
rect 940 55632 992 55684
rect 24584 55675 24636 55684
rect 24584 55641 24593 55675
rect 24593 55641 24627 55675
rect 24627 55641 24636 55675
rect 24584 55632 24636 55641
rect 25688 55743 25740 55752
rect 25688 55709 25697 55743
rect 25697 55709 25731 55743
rect 25731 55709 25740 55743
rect 25688 55700 25740 55709
rect 29736 55675 29788 55684
rect 29736 55641 29745 55675
rect 29745 55641 29779 55675
rect 29779 55641 29788 55675
rect 29736 55632 29788 55641
rect 30380 55743 30432 55752
rect 30380 55709 30389 55743
rect 30389 55709 30423 55743
rect 30423 55709 30432 55743
rect 30380 55700 30432 55709
rect 30472 55743 30524 55752
rect 30472 55709 30481 55743
rect 30481 55709 30515 55743
rect 30515 55709 30524 55743
rect 30472 55700 30524 55709
rect 40040 55700 40092 55752
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 24308 55360 24360 55412
rect 25688 55360 25740 55412
rect 940 55224 992 55276
rect 23940 55224 23992 55276
rect 24032 55224 24084 55276
rect 24400 55267 24452 55276
rect 24400 55233 24409 55267
rect 24409 55233 24443 55267
rect 24443 55233 24452 55267
rect 24400 55224 24452 55233
rect 24768 55267 24820 55276
rect 24768 55233 24777 55267
rect 24777 55233 24811 55267
rect 24811 55233 24820 55267
rect 24768 55224 24820 55233
rect 24952 55267 25004 55276
rect 24952 55233 24961 55267
rect 24961 55233 24995 55267
rect 24995 55233 25004 55267
rect 24952 55224 25004 55233
rect 25320 55224 25372 55276
rect 41512 55360 41564 55412
rect 44180 55292 44232 55344
rect 41052 55267 41104 55276
rect 41052 55233 41061 55267
rect 41061 55233 41095 55267
rect 41095 55233 41104 55267
rect 41052 55224 41104 55233
rect 41236 55267 41288 55276
rect 41236 55233 41250 55267
rect 41250 55233 41284 55267
rect 41284 55233 41288 55267
rect 41236 55224 41288 55233
rect 42064 55224 42116 55276
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 28724 54680 28776 54732
rect 23572 54655 23624 54664
rect 23572 54621 23581 54655
rect 23581 54621 23615 54655
rect 23615 54621 23624 54655
rect 23572 54612 23624 54621
rect 940 54544 992 54596
rect 22100 54544 22152 54596
rect 24308 54612 24360 54664
rect 58348 54655 58400 54664
rect 58348 54621 58357 54655
rect 58357 54621 58391 54655
rect 58391 54621 58400 54655
rect 58348 54612 58400 54621
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 940 54136 992 54188
rect 1768 53975 1820 53984
rect 1768 53941 1777 53975
rect 1777 53941 1811 53975
rect 1811 53941 1820 53975
rect 1768 53932 1820 53941
rect 23572 53932 23624 53984
rect 24216 53932 24268 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 40132 53660 40184 53712
rect 24952 53592 25004 53644
rect 41052 53592 41104 53644
rect 21272 53456 21324 53508
rect 24400 53456 24452 53508
rect 1768 53388 1820 53440
rect 41236 53524 41288 53576
rect 44824 53456 44876 53508
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 24952 53184 25004 53236
rect 940 53048 992 53100
rect 23664 53048 23716 53100
rect 24400 53048 24452 53100
rect 45376 53048 45428 53100
rect 23848 52844 23900 52896
rect 58348 52887 58400 52896
rect 58348 52853 58357 52887
rect 58357 52853 58391 52887
rect 58391 52853 58400 52887
rect 58348 52844 58400 52853
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 24952 52683 25004 52692
rect 24952 52649 24961 52683
rect 24961 52649 24995 52683
rect 24995 52649 25004 52683
rect 24952 52640 25004 52649
rect 2044 52479 2096 52488
rect 2044 52445 2053 52479
rect 2053 52445 2087 52479
rect 2087 52445 2096 52479
rect 2044 52436 2096 52445
rect 940 52368 992 52420
rect 21456 52368 21508 52420
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 20260 52096 20312 52148
rect 940 51960 992 52012
rect 8024 52003 8076 52012
rect 8024 51969 8033 52003
rect 8033 51969 8067 52003
rect 8067 51969 8076 52003
rect 8024 51960 8076 51969
rect 8300 52003 8352 52012
rect 8300 51969 8309 52003
rect 8309 51969 8343 52003
rect 8343 51969 8352 52003
rect 8300 51960 8352 51969
rect 22192 51960 22244 52012
rect 22836 51960 22888 52012
rect 17868 51892 17920 51944
rect 7840 51799 7892 51808
rect 7840 51765 7849 51799
rect 7849 51765 7883 51799
rect 7883 51765 7892 51799
rect 7840 51756 7892 51765
rect 20536 51799 20588 51808
rect 20536 51765 20545 51799
rect 20545 51765 20579 51799
rect 20579 51765 20588 51799
rect 20536 51756 20588 51765
rect 24216 51756 24268 51808
rect 41144 51756 41196 51808
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 58348 51391 58400 51400
rect 58348 51357 58357 51391
rect 58357 51357 58391 51391
rect 58391 51357 58400 51391
rect 58348 51348 58400 51357
rect 940 51280 992 51332
rect 3976 51280 4028 51332
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 2688 50940 2740 50992
rect 3976 50983 4028 50992
rect 3976 50949 3985 50983
rect 3985 50949 4019 50983
rect 4019 50949 4028 50983
rect 3976 50940 4028 50949
rect 4068 50915 4120 50924
rect 4068 50881 4082 50915
rect 4082 50881 4116 50915
rect 4116 50881 4120 50915
rect 4068 50872 4120 50881
rect 4620 50804 4672 50856
rect 6276 50668 6328 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 27344 50396 27396 50448
rect 40776 50396 40828 50448
rect 6000 50328 6052 50380
rect 29552 50328 29604 50380
rect 32680 50328 32732 50380
rect 33232 50328 33284 50380
rect 36544 50328 36596 50380
rect 56600 50328 56652 50380
rect 57520 50260 57572 50312
rect 940 50192 992 50244
rect 2044 50192 2096 50244
rect 58992 50192 59044 50244
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 940 49784 992 49836
rect 4068 49784 4120 49836
rect 6828 49784 6880 49836
rect 8300 49784 8352 49836
rect 13084 49716 13136 49768
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 940 49172 992 49224
rect 57980 49147 58032 49156
rect 57980 49113 57989 49147
rect 57989 49113 58023 49147
rect 58023 49113 58032 49147
rect 57980 49104 58032 49113
rect 59452 49104 59504 49156
rect 6460 49036 6512 49088
rect 25412 49036 25464 49088
rect 43076 49036 43128 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 940 48696 992 48748
rect 1952 48560 2004 48612
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 17868 48220 17920 48272
rect 55956 48220 56008 48272
rect 58072 48220 58124 48272
rect 2044 48127 2096 48136
rect 2044 48093 2053 48127
rect 2053 48093 2087 48127
rect 2087 48093 2096 48127
rect 2044 48084 2096 48093
rect 4068 48152 4120 48204
rect 6828 48152 6880 48204
rect 9036 48152 9088 48204
rect 2412 48127 2464 48136
rect 2412 48093 2426 48127
rect 2426 48093 2460 48127
rect 2460 48093 2464 48127
rect 2412 48084 2464 48093
rect 57796 48084 57848 48136
rect 1584 47948 1636 48000
rect 58164 48059 58216 48068
rect 58164 48025 58173 48059
rect 58173 48025 58207 48059
rect 58207 48025 58216 48059
rect 58164 48016 58216 48025
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 31300 47744 31352 47796
rect 40408 47744 40460 47796
rect 30656 47676 30708 47728
rect 44088 47676 44140 47728
rect 940 47608 992 47660
rect 9128 47608 9180 47660
rect 34520 47608 34572 47660
rect 58072 47651 58124 47660
rect 58072 47617 58081 47651
rect 58081 47617 58115 47651
rect 58115 47617 58124 47651
rect 58072 47608 58124 47617
rect 3424 47540 3476 47592
rect 32220 47540 32272 47592
rect 1768 47447 1820 47456
rect 1768 47413 1777 47447
rect 1777 47413 1811 47447
rect 1811 47413 1820 47447
rect 1768 47404 1820 47413
rect 58808 47404 58860 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 8944 47132 8996 47184
rect 940 46996 992 47048
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 940 46520 992 46572
rect 36360 46316 36412 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 58164 46019 58216 46028
rect 58164 45985 58173 46019
rect 58173 45985 58207 46019
rect 58207 45985 58216 46019
rect 58164 45976 58216 45985
rect 57704 45908 57756 45960
rect 940 45840 992 45892
rect 15200 45772 15252 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 15200 45500 15252 45552
rect 17500 45543 17552 45552
rect 17500 45509 17509 45543
rect 17509 45509 17543 45543
rect 17543 45509 17552 45543
rect 17500 45500 17552 45509
rect 21088 45432 21140 45484
rect 9036 45296 9088 45348
rect 21456 45364 21508 45416
rect 33784 45500 33836 45552
rect 57060 45500 57112 45552
rect 36360 45475 36412 45484
rect 36360 45441 36369 45475
rect 36369 45441 36403 45475
rect 36403 45441 36412 45475
rect 36360 45432 36412 45441
rect 36636 45475 36688 45484
rect 36636 45441 36645 45475
rect 36645 45441 36679 45475
rect 36679 45441 36688 45475
rect 36636 45432 36688 45441
rect 37372 45432 37424 45484
rect 38016 45475 38068 45484
rect 38016 45441 38025 45475
rect 38025 45441 38059 45475
rect 38059 45441 38068 45475
rect 38016 45432 38068 45441
rect 38476 45475 38528 45484
rect 38476 45441 38479 45475
rect 38479 45441 38528 45475
rect 38476 45432 38528 45441
rect 58992 45432 59044 45484
rect 36912 45339 36964 45348
rect 36912 45305 36921 45339
rect 36921 45305 36955 45339
rect 36955 45305 36964 45339
rect 36912 45296 36964 45305
rect 17776 45271 17828 45280
rect 17776 45237 17785 45271
rect 17785 45237 17819 45271
rect 17819 45237 17828 45271
rect 17776 45228 17828 45237
rect 58440 45228 58492 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 35440 45067 35492 45076
rect 35440 45033 35449 45067
rect 35449 45033 35483 45067
rect 35483 45033 35492 45067
rect 35440 45024 35492 45033
rect 21272 44888 21324 44940
rect 35256 44956 35308 45008
rect 940 44820 992 44872
rect 1860 44863 1912 44872
rect 1860 44829 1869 44863
rect 1869 44829 1903 44863
rect 1903 44829 1912 44863
rect 1860 44820 1912 44829
rect 35072 44863 35124 44872
rect 35072 44829 35081 44863
rect 35081 44829 35115 44863
rect 35115 44829 35124 44863
rect 35072 44820 35124 44829
rect 35256 44863 35308 44872
rect 35256 44829 35270 44863
rect 35270 44829 35304 44863
rect 35304 44829 35308 44863
rect 35256 44820 35308 44829
rect 45744 44820 45796 44872
rect 56968 44863 57020 44872
rect 56968 44829 56977 44863
rect 56977 44829 57011 44863
rect 57011 44829 57020 44863
rect 56968 44820 57020 44829
rect 58992 44820 59044 44872
rect 9220 44752 9272 44804
rect 58716 44752 58768 44804
rect 58348 44684 58400 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 940 44344 992 44396
rect 9588 44208 9640 44260
rect 34704 44140 34756 44192
rect 35072 44140 35124 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 34244 43911 34296 43920
rect 34244 43877 34253 43911
rect 34253 43877 34287 43911
rect 34287 43877 34296 43911
rect 34244 43868 34296 43877
rect 9588 43732 9640 43784
rect 34060 43775 34112 43784
rect 34060 43741 34074 43775
rect 34074 43741 34108 43775
rect 34108 43741 34112 43775
rect 34060 43732 34112 43741
rect 53840 43732 53892 43784
rect 940 43664 992 43716
rect 33784 43664 33836 43716
rect 35900 43664 35952 43716
rect 58164 43707 58216 43716
rect 58164 43673 58173 43707
rect 58173 43673 58207 43707
rect 58207 43673 58216 43707
rect 58164 43664 58216 43673
rect 32312 43596 32364 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 940 43256 992 43308
rect 32312 43299 32364 43308
rect 32312 43265 32321 43299
rect 32321 43265 32355 43299
rect 32355 43265 32364 43299
rect 32312 43256 32364 43265
rect 32496 43299 32548 43308
rect 32496 43265 32505 43299
rect 32505 43265 32539 43299
rect 32539 43265 32548 43299
rect 32496 43256 32548 43265
rect 32680 43299 32732 43308
rect 32680 43265 32694 43299
rect 32694 43265 32728 43299
rect 32728 43265 32732 43299
rect 32680 43256 32732 43265
rect 54852 43256 54904 43308
rect 1768 43095 1820 43104
rect 1768 43061 1777 43095
rect 1777 43061 1811 43095
rect 1811 43061 1820 43095
rect 1768 43052 1820 43061
rect 31760 43052 31812 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 32680 42780 32732 42832
rect 24308 42712 24360 42764
rect 32496 42712 32548 42764
rect 33048 42687 33100 42696
rect 22192 42576 22244 42628
rect 24400 42576 24452 42628
rect 33048 42653 33057 42687
rect 33057 42653 33091 42687
rect 33091 42653 33100 42687
rect 33048 42644 33100 42653
rect 33140 42687 33192 42696
rect 33140 42653 33149 42687
rect 33149 42653 33183 42687
rect 33183 42653 33192 42687
rect 33140 42644 33192 42653
rect 33784 42712 33836 42764
rect 32036 42576 32088 42628
rect 33876 42687 33928 42696
rect 33876 42653 33885 42687
rect 33885 42653 33919 42687
rect 33919 42653 33928 42687
rect 33876 42644 33928 42653
rect 37280 42687 37332 42696
rect 37280 42653 37289 42687
rect 37289 42653 37323 42687
rect 37323 42653 37332 42687
rect 37280 42644 37332 42653
rect 58992 42644 59044 42696
rect 37372 42576 37424 42628
rect 54300 42576 54352 42628
rect 57980 42619 58032 42628
rect 57980 42585 57989 42619
rect 57989 42585 58023 42619
rect 58023 42585 58032 42619
rect 57980 42576 58032 42585
rect 58532 42576 58584 42628
rect 39304 42508 39356 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 37280 42304 37332 42356
rect 39396 42304 39448 42356
rect 940 42168 992 42220
rect 1768 42168 1820 42220
rect 33876 42168 33928 42220
rect 13084 42100 13136 42152
rect 23664 42100 23716 42152
rect 33140 42100 33192 42152
rect 33784 42100 33836 42152
rect 34060 42100 34112 42152
rect 6460 42032 6512 42084
rect 22560 42032 22612 42084
rect 2136 41964 2188 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 53564 41556 53616 41608
rect 58992 41556 59044 41608
rect 940 41488 992 41540
rect 6368 41488 6420 41540
rect 58716 41488 58768 41540
rect 50068 41420 50120 41472
rect 53840 41420 53892 41472
rect 58624 41420 58676 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 940 41080 992 41132
rect 21180 40876 21232 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 28448 40672 28500 40724
rect 41420 40672 41472 40724
rect 54668 40468 54720 40520
rect 940 40400 992 40452
rect 11704 40332 11756 40384
rect 56048 40332 56100 40384
rect 58992 40400 59044 40452
rect 58716 40332 58768 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 20904 40128 20956 40180
rect 58348 40128 58400 40180
rect 58716 40128 58768 40180
rect 1032 40060 1084 40112
rect 21088 40103 21140 40112
rect 21088 40069 21097 40103
rect 21097 40069 21131 40103
rect 21131 40069 21140 40103
rect 21088 40060 21140 40069
rect 21180 40103 21232 40112
rect 21180 40069 21189 40103
rect 21189 40069 21223 40103
rect 21223 40069 21232 40103
rect 21180 40060 21232 40069
rect 21640 39992 21692 40044
rect 2596 39788 2648 39840
rect 22284 39788 22336 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 2688 39516 2740 39568
rect 22652 39516 22704 39568
rect 2228 39448 2280 39500
rect 2320 39423 2372 39432
rect 2320 39389 2329 39423
rect 2329 39389 2363 39423
rect 2363 39389 2372 39423
rect 2320 39380 2372 39389
rect 2596 39423 2648 39432
rect 2596 39389 2605 39423
rect 2605 39389 2639 39423
rect 2639 39389 2648 39423
rect 2596 39380 2648 39389
rect 2688 39423 2740 39432
rect 2688 39389 2702 39423
rect 2702 39389 2736 39423
rect 2736 39389 2740 39423
rect 2688 39380 2740 39389
rect 58992 39380 59044 39432
rect 940 39312 992 39364
rect 29644 39312 29696 39364
rect 53472 39312 53524 39364
rect 57980 39355 58032 39364
rect 57980 39321 57989 39355
rect 57989 39321 58023 39355
rect 58023 39321 58032 39355
rect 57980 39312 58032 39321
rect 58348 39355 58400 39364
rect 58348 39321 58357 39355
rect 58357 39321 58391 39355
rect 58391 39321 58400 39355
rect 58348 39312 58400 39321
rect 3056 39244 3108 39296
rect 33508 39244 33560 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 1032 38904 1084 38956
rect 20536 38904 20588 38956
rect 22284 38947 22336 38956
rect 22284 38913 22293 38947
rect 22293 38913 22327 38947
rect 22327 38913 22336 38947
rect 22284 38904 22336 38913
rect 22468 38879 22520 38888
rect 22468 38845 22477 38879
rect 22477 38845 22511 38879
rect 22511 38845 22520 38879
rect 22468 38836 22520 38845
rect 19984 38768 20036 38820
rect 20260 38768 20312 38820
rect 23112 38811 23164 38820
rect 23112 38777 23121 38811
rect 23121 38777 23155 38811
rect 23155 38777 23164 38811
rect 23112 38768 23164 38777
rect 19432 38700 19484 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 16212 38496 16264 38548
rect 20904 38496 20956 38548
rect 21088 38496 21140 38548
rect 25320 38496 25372 38548
rect 1860 38428 1912 38480
rect 20996 38428 21048 38480
rect 23112 38428 23164 38480
rect 1676 38360 1728 38412
rect 1952 38292 2004 38344
rect 2412 38335 2464 38344
rect 2412 38301 2421 38335
rect 2421 38301 2455 38335
rect 2455 38301 2464 38335
rect 2412 38292 2464 38301
rect 3056 38403 3108 38412
rect 3056 38369 3065 38403
rect 3065 38369 3099 38403
rect 3099 38369 3108 38403
rect 3056 38360 3108 38369
rect 11704 38360 11756 38412
rect 2688 38292 2740 38344
rect 20352 38335 20404 38344
rect 20352 38301 20361 38335
rect 20361 38301 20395 38335
rect 20395 38301 20404 38335
rect 20352 38292 20404 38301
rect 2320 38267 2372 38276
rect 2320 38233 2329 38267
rect 2329 38233 2363 38267
rect 2363 38233 2372 38267
rect 2320 38224 2372 38233
rect 19248 38224 19300 38276
rect 20168 38224 20220 38276
rect 20720 38360 20772 38412
rect 23388 38428 23440 38480
rect 22928 38335 22980 38344
rect 22928 38301 22937 38335
rect 22937 38301 22971 38335
rect 22971 38301 22980 38335
rect 22928 38292 22980 38301
rect 26976 38360 27028 38412
rect 23388 38335 23440 38344
rect 23388 38301 23402 38335
rect 23402 38301 23436 38335
rect 23436 38301 23440 38335
rect 23388 38292 23440 38301
rect 46848 38292 46900 38344
rect 2596 38199 2648 38208
rect 2596 38165 2605 38199
rect 2605 38165 2639 38199
rect 2639 38165 2648 38199
rect 2596 38156 2648 38165
rect 20352 38156 20404 38208
rect 21732 38156 21784 38208
rect 23204 38267 23256 38276
rect 23204 38233 23213 38267
rect 23213 38233 23247 38267
rect 23247 38233 23256 38267
rect 23204 38224 23256 38233
rect 58164 38267 58216 38276
rect 58164 38233 58173 38267
rect 58173 38233 58207 38267
rect 58207 38233 58216 38267
rect 58164 38224 58216 38233
rect 23572 38199 23624 38208
rect 23572 38165 23581 38199
rect 23581 38165 23615 38199
rect 23615 38165 23624 38199
rect 23572 38156 23624 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 2596 37952 2648 38004
rect 16212 37952 16264 38004
rect 5908 37884 5960 37936
rect 19708 37927 19760 37936
rect 19708 37893 19714 37927
rect 19714 37893 19748 37927
rect 19748 37893 19760 37927
rect 19708 37884 19760 37893
rect 20812 37952 20864 38004
rect 20996 37995 21048 38004
rect 20996 37961 21005 37995
rect 21005 37961 21039 37995
rect 21039 37961 21048 37995
rect 20996 37952 21048 37961
rect 940 37816 992 37868
rect 16672 37816 16724 37868
rect 19340 37859 19392 37868
rect 19340 37825 19349 37859
rect 19349 37825 19383 37859
rect 19383 37825 19392 37859
rect 19340 37816 19392 37825
rect 1860 37723 1912 37732
rect 1860 37689 1869 37723
rect 1869 37689 1903 37723
rect 1903 37689 1912 37723
rect 1860 37680 1912 37689
rect 20720 37816 20772 37868
rect 20812 37859 20864 37868
rect 20812 37825 20821 37859
rect 20821 37825 20855 37859
rect 20855 37825 20864 37859
rect 20812 37816 20864 37825
rect 21088 37859 21140 37868
rect 21088 37825 21097 37859
rect 21097 37825 21131 37859
rect 21131 37825 21140 37859
rect 21088 37816 21140 37825
rect 21364 37816 21416 37868
rect 22836 37884 22888 37936
rect 24768 37884 24820 37936
rect 23020 37859 23072 37868
rect 23020 37825 23029 37859
rect 23029 37825 23063 37859
rect 23063 37825 23072 37859
rect 23020 37816 23072 37825
rect 20628 37748 20680 37800
rect 21456 37748 21508 37800
rect 19800 37680 19852 37732
rect 19984 37655 20036 37664
rect 19984 37621 19993 37655
rect 19993 37621 20027 37655
rect 20027 37621 20036 37655
rect 19984 37612 20036 37621
rect 20628 37655 20680 37664
rect 20628 37621 20637 37655
rect 20637 37621 20671 37655
rect 20671 37621 20680 37655
rect 20628 37612 20680 37621
rect 20812 37680 20864 37732
rect 23848 37816 23900 37868
rect 24124 37791 24176 37800
rect 24124 37757 24133 37791
rect 24133 37757 24167 37791
rect 24167 37757 24176 37791
rect 24124 37748 24176 37757
rect 24400 37748 24452 37800
rect 25136 37859 25188 37868
rect 25136 37825 25145 37859
rect 25145 37825 25179 37859
rect 25179 37825 25188 37859
rect 25136 37816 25188 37825
rect 25320 37859 25372 37868
rect 25320 37825 25329 37859
rect 25329 37825 25363 37859
rect 25363 37825 25372 37859
rect 25320 37816 25372 37825
rect 58072 37859 58124 37868
rect 58072 37825 58081 37859
rect 58081 37825 58115 37859
rect 58115 37825 58124 37859
rect 58072 37816 58124 37825
rect 28264 37748 28316 37800
rect 22836 37612 22888 37664
rect 24032 37612 24084 37664
rect 59176 37612 59228 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19248 37408 19300 37460
rect 21088 37408 21140 37460
rect 19800 37340 19852 37392
rect 20352 37340 20404 37392
rect 20720 37340 20772 37392
rect 22192 37340 22244 37392
rect 6000 37247 6052 37256
rect 6000 37213 6009 37247
rect 6009 37213 6043 37247
rect 6043 37213 6052 37247
rect 6000 37204 6052 37213
rect 6276 37247 6328 37256
rect 6276 37213 6285 37247
rect 6285 37213 6319 37247
rect 6319 37213 6328 37247
rect 6276 37204 6328 37213
rect 2412 37136 2464 37188
rect 5540 37111 5592 37120
rect 5540 37077 5549 37111
rect 5549 37077 5583 37111
rect 5583 37077 5592 37111
rect 5540 37068 5592 37077
rect 6736 37247 6788 37256
rect 6736 37213 6745 37247
rect 6745 37213 6779 37247
rect 6779 37213 6788 37247
rect 6736 37204 6788 37213
rect 19340 37204 19392 37256
rect 18880 37136 18932 37188
rect 20904 37272 20956 37324
rect 21088 37315 21140 37324
rect 21088 37281 21097 37315
rect 21097 37281 21131 37315
rect 21131 37281 21140 37315
rect 21088 37272 21140 37281
rect 31116 37272 31168 37324
rect 33508 37272 33560 37324
rect 20536 37204 20588 37256
rect 20168 37179 20220 37188
rect 20168 37145 20177 37179
rect 20177 37145 20211 37179
rect 20211 37145 20220 37179
rect 20168 37136 20220 37145
rect 28356 37204 28408 37256
rect 53472 37204 53524 37256
rect 53748 37247 53800 37256
rect 53748 37213 53757 37247
rect 53757 37213 53791 37247
rect 53791 37213 53800 37247
rect 53748 37204 53800 37213
rect 54484 37204 54536 37256
rect 20444 37068 20496 37120
rect 53840 37136 53892 37188
rect 56692 37136 56744 37188
rect 58164 37179 58216 37188
rect 58164 37145 58173 37179
rect 58173 37145 58207 37179
rect 58207 37145 58216 37179
rect 58164 37136 58216 37145
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 6000 36864 6052 36916
rect 42984 36864 43036 36916
rect 21824 36796 21876 36848
rect 940 36728 992 36780
rect 16580 36728 16632 36780
rect 18880 36771 18932 36780
rect 18880 36737 18889 36771
rect 18889 36737 18923 36771
rect 18923 36737 18932 36771
rect 18880 36728 18932 36737
rect 19248 36660 19300 36712
rect 19432 36728 19484 36780
rect 20720 36728 20772 36780
rect 23940 36728 23992 36780
rect 24124 36728 24176 36780
rect 21180 36660 21232 36712
rect 23848 36703 23900 36712
rect 23848 36669 23857 36703
rect 23857 36669 23891 36703
rect 23891 36669 23900 36703
rect 23848 36660 23900 36669
rect 57336 36796 57388 36848
rect 53656 36771 53708 36780
rect 53656 36737 53665 36771
rect 53665 36737 53699 36771
rect 53699 36737 53708 36771
rect 53656 36728 53708 36737
rect 53840 36771 53892 36780
rect 53840 36737 53849 36771
rect 53849 36737 53883 36771
rect 53883 36737 53892 36771
rect 53840 36728 53892 36737
rect 39948 36660 40000 36712
rect 21824 36592 21876 36644
rect 39120 36592 39172 36644
rect 40868 36592 40920 36644
rect 53472 36592 53524 36644
rect 3424 36524 3476 36576
rect 20996 36567 21048 36576
rect 20996 36533 21005 36567
rect 21005 36533 21039 36567
rect 21039 36533 21048 36567
rect 20996 36524 21048 36533
rect 21364 36567 21416 36576
rect 21364 36533 21373 36567
rect 21373 36533 21407 36567
rect 21407 36533 21416 36567
rect 21364 36524 21416 36533
rect 23480 36524 23532 36576
rect 24584 36524 24636 36576
rect 54208 36567 54260 36576
rect 54208 36533 54217 36567
rect 54217 36533 54251 36567
rect 54251 36533 54260 36567
rect 54208 36524 54260 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 6736 36320 6788 36372
rect 23480 36320 23532 36372
rect 23848 36363 23900 36372
rect 23848 36329 23857 36363
rect 23857 36329 23891 36363
rect 23891 36329 23900 36363
rect 23848 36320 23900 36329
rect 2412 36184 2464 36236
rect 2504 36159 2556 36168
rect 2504 36125 2513 36159
rect 2513 36125 2547 36159
rect 2547 36125 2556 36159
rect 2504 36116 2556 36125
rect 21364 36252 21416 36304
rect 21456 36252 21508 36304
rect 54208 36320 54260 36372
rect 20628 36184 20680 36236
rect 20720 36227 20772 36236
rect 20720 36193 20729 36227
rect 20729 36193 20763 36227
rect 20763 36193 20772 36227
rect 20720 36184 20772 36193
rect 940 36048 992 36100
rect 2228 36048 2280 36100
rect 2780 36091 2832 36100
rect 2780 36057 2789 36091
rect 2789 36057 2823 36091
rect 2823 36057 2832 36091
rect 2780 36048 2832 36057
rect 16672 36048 16724 36100
rect 19984 36048 20036 36100
rect 22284 36159 22336 36168
rect 22284 36125 22293 36159
rect 22293 36125 22327 36159
rect 22327 36125 22336 36159
rect 22284 36116 22336 36125
rect 22560 36159 22612 36168
rect 22560 36125 22569 36159
rect 22569 36125 22603 36159
rect 22603 36125 22612 36159
rect 22560 36116 22612 36125
rect 23572 36184 23624 36236
rect 23296 36159 23348 36168
rect 23296 36125 23305 36159
rect 23305 36125 23339 36159
rect 23339 36125 23348 36159
rect 23296 36116 23348 36125
rect 23388 36116 23440 36168
rect 24308 36116 24360 36168
rect 24584 36159 24636 36168
rect 24584 36125 24593 36159
rect 24593 36125 24627 36159
rect 24627 36125 24636 36159
rect 24584 36116 24636 36125
rect 22192 35980 22244 36032
rect 22744 35980 22796 36032
rect 23572 36091 23624 36100
rect 23572 36057 23581 36091
rect 23581 36057 23615 36091
rect 23615 36057 23624 36091
rect 23572 36048 23624 36057
rect 25228 36048 25280 36100
rect 57980 36091 58032 36100
rect 57980 36057 57989 36091
rect 57989 36057 58023 36091
rect 58023 36057 58032 36091
rect 57980 36048 58032 36057
rect 59268 36048 59320 36100
rect 24952 35980 25004 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 1584 35776 1636 35828
rect 20996 35776 21048 35828
rect 25136 35776 25188 35828
rect 18788 35708 18840 35760
rect 21088 35708 21140 35760
rect 940 35640 992 35692
rect 18880 35640 18932 35692
rect 20168 35640 20220 35692
rect 41696 35776 41748 35828
rect 21088 35572 21140 35624
rect 23388 35615 23440 35624
rect 23388 35581 23397 35615
rect 23397 35581 23431 35615
rect 23431 35581 23440 35615
rect 23388 35572 23440 35581
rect 40592 35683 40644 35692
rect 40592 35649 40601 35683
rect 40601 35649 40635 35683
rect 40635 35649 40644 35683
rect 40592 35640 40644 35649
rect 47676 35572 47728 35624
rect 39948 35504 40000 35556
rect 18880 35479 18932 35488
rect 18880 35445 18889 35479
rect 18889 35445 18923 35479
rect 18923 35445 18932 35479
rect 18880 35436 18932 35445
rect 33784 35436 33836 35488
rect 40592 35436 40644 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 22744 35275 22796 35284
rect 22744 35241 22753 35275
rect 22753 35241 22787 35275
rect 22787 35241 22796 35275
rect 22744 35232 22796 35241
rect 23572 35232 23624 35284
rect 37372 35232 37424 35284
rect 2780 35164 2832 35216
rect 22284 35164 22336 35216
rect 55680 35164 55732 35216
rect 21180 35028 21232 35080
rect 24400 35028 24452 35080
rect 26976 35028 27028 35080
rect 940 34960 992 35012
rect 22652 34960 22704 35012
rect 22928 34935 22980 34944
rect 22928 34901 22937 34935
rect 22937 34901 22971 34935
rect 22971 34901 22980 34935
rect 22928 34892 22980 34901
rect 40040 35071 40092 35080
rect 40040 35037 40049 35071
rect 40049 35037 40083 35071
rect 40083 35037 40092 35071
rect 40040 35028 40092 35037
rect 40316 35071 40368 35080
rect 40316 35037 40325 35071
rect 40325 35037 40359 35071
rect 40359 35037 40368 35071
rect 40316 35028 40368 35037
rect 40500 35028 40552 35080
rect 54944 35028 54996 35080
rect 37372 34960 37424 35012
rect 58164 35003 58216 35012
rect 58164 34969 58173 35003
rect 58173 34969 58207 35003
rect 58207 34969 58216 35003
rect 58164 34960 58216 34969
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 20260 34688 20312 34740
rect 22376 34688 22428 34740
rect 59360 34688 59412 34740
rect 19432 34620 19484 34672
rect 24860 34620 24912 34672
rect 58992 34552 59044 34604
rect 20076 34484 20128 34536
rect 23388 34484 23440 34536
rect 47584 34484 47636 34536
rect 54668 34484 54720 34536
rect 40040 34416 40092 34468
rect 44364 34416 44416 34468
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 21088 34144 21140 34196
rect 23572 34144 23624 34196
rect 23848 34144 23900 34196
rect 40040 34144 40092 34196
rect 40500 34144 40552 34196
rect 17316 34076 17368 34128
rect 940 33940 992 33992
rect 21916 34008 21968 34060
rect 21456 33983 21508 33992
rect 21456 33949 21463 33983
rect 21463 33949 21508 33983
rect 21456 33940 21508 33949
rect 21548 33983 21600 33992
rect 21548 33949 21557 33983
rect 21557 33949 21591 33983
rect 21591 33949 21600 33983
rect 21548 33940 21600 33949
rect 21824 33940 21876 33992
rect 22928 33983 22980 33992
rect 22928 33949 22937 33983
rect 22937 33949 22971 33983
rect 22971 33949 22980 33983
rect 22928 33940 22980 33949
rect 23112 33872 23164 33924
rect 23480 34076 23532 34128
rect 24492 33940 24544 33992
rect 24768 33983 24820 33992
rect 24768 33949 24775 33983
rect 24775 33949 24820 33983
rect 24768 33940 24820 33949
rect 24952 34008 25004 34060
rect 25044 33804 25096 33856
rect 35900 33804 35952 33856
rect 36544 33804 36596 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 2320 33532 2372 33584
rect 12164 33532 12216 33584
rect 22376 33575 22428 33584
rect 22376 33541 22385 33575
rect 22385 33541 22419 33575
rect 22419 33541 22428 33575
rect 22376 33532 22428 33541
rect 24860 33600 24912 33652
rect 31024 33600 31076 33652
rect 34704 33532 34756 33584
rect 38476 33600 38528 33652
rect 940 33464 992 33516
rect 20904 33507 20956 33516
rect 20904 33473 20913 33507
rect 20913 33473 20947 33507
rect 20947 33473 20956 33507
rect 20904 33464 20956 33473
rect 21088 33507 21140 33516
rect 21088 33473 21097 33507
rect 21097 33473 21131 33507
rect 21131 33473 21140 33507
rect 21088 33464 21140 33473
rect 21272 33507 21324 33516
rect 21272 33473 21281 33507
rect 21281 33473 21315 33507
rect 21315 33473 21324 33507
rect 21272 33464 21324 33473
rect 20352 33396 20404 33448
rect 20628 33396 20680 33448
rect 22284 33507 22336 33516
rect 22284 33473 22293 33507
rect 22293 33473 22327 33507
rect 22327 33473 22336 33507
rect 22284 33464 22336 33473
rect 23480 33464 23532 33516
rect 24952 33396 25004 33448
rect 23572 33328 23624 33380
rect 35900 33507 35952 33516
rect 35900 33473 35907 33507
rect 35907 33473 35952 33507
rect 35900 33464 35952 33473
rect 36084 33575 36136 33584
rect 36084 33541 36093 33575
rect 36093 33541 36127 33575
rect 36127 33541 36136 33575
rect 36084 33532 36136 33541
rect 40040 33464 40092 33516
rect 22652 33303 22704 33312
rect 22652 33269 22661 33303
rect 22661 33269 22695 33303
rect 22695 33269 22704 33303
rect 22652 33260 22704 33269
rect 23388 33260 23440 33312
rect 31024 33260 31076 33312
rect 37832 33260 37884 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 22652 32988 22704 33040
rect 58992 32920 59044 32972
rect 21732 32895 21784 32904
rect 21732 32861 21741 32895
rect 21741 32861 21775 32895
rect 21775 32861 21784 32895
rect 21732 32852 21784 32861
rect 23572 32852 23624 32904
rect 57428 32852 57480 32904
rect 940 32784 992 32836
rect 22560 32784 22612 32836
rect 58992 32784 59044 32836
rect 16580 32716 16632 32768
rect 54760 32716 54812 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 24768 32512 24820 32564
rect 54024 32512 54076 32564
rect 23296 32444 23348 32496
rect 53288 32444 53340 32496
rect 940 32376 992 32428
rect 1860 32376 1912 32428
rect 22008 32376 22060 32428
rect 24860 32419 24912 32428
rect 24860 32385 24869 32419
rect 24869 32385 24903 32419
rect 24903 32385 24912 32419
rect 24860 32376 24912 32385
rect 25044 32376 25096 32428
rect 37556 32376 37608 32428
rect 25228 32308 25280 32360
rect 23020 32172 23072 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 59544 31900 59596 31952
rect 16764 31764 16816 31816
rect 21824 31764 21876 31816
rect 23020 31807 23072 31816
rect 23020 31773 23029 31807
rect 23029 31773 23063 31807
rect 23063 31773 23072 31807
rect 23020 31764 23072 31773
rect 23388 31807 23440 31816
rect 23388 31773 23397 31807
rect 23397 31773 23431 31807
rect 23431 31773 23440 31807
rect 23388 31764 23440 31773
rect 48964 31764 49016 31816
rect 58992 31764 59044 31816
rect 23572 31671 23624 31680
rect 23572 31637 23581 31671
rect 23581 31637 23615 31671
rect 23615 31637 23624 31671
rect 23572 31628 23624 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 24308 31424 24360 31476
rect 24860 31467 24912 31476
rect 24860 31433 24869 31467
rect 24869 31433 24903 31467
rect 24903 31433 24912 31467
rect 24860 31424 24912 31433
rect 940 31288 992 31340
rect 24216 31331 24268 31340
rect 24216 31297 24225 31331
rect 24225 31297 24259 31331
rect 24259 31297 24268 31331
rect 24216 31288 24268 31297
rect 24400 31331 24452 31340
rect 24400 31297 24407 31331
rect 24407 31297 24452 31331
rect 24400 31288 24452 31297
rect 21548 31220 21600 31272
rect 23020 31220 23072 31272
rect 23480 31152 23532 31204
rect 24124 31152 24176 31204
rect 24216 31152 24268 31204
rect 58072 31331 58124 31340
rect 58072 31297 58081 31331
rect 58081 31297 58115 31331
rect 58115 31297 58124 31331
rect 58072 31288 58124 31297
rect 24952 31152 25004 31204
rect 47492 31152 47544 31204
rect 36360 31084 36412 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 24400 30880 24452 30932
rect 40684 30880 40736 30932
rect 19432 30812 19484 30864
rect 34796 30744 34848 30796
rect 940 30608 992 30660
rect 17776 30608 17828 30660
rect 22836 30719 22888 30728
rect 22836 30685 22845 30719
rect 22845 30685 22879 30719
rect 22879 30685 22888 30719
rect 22836 30676 22888 30685
rect 22008 30608 22060 30660
rect 23204 30719 23256 30728
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 23020 30651 23072 30660
rect 23020 30617 23029 30651
rect 23029 30617 23063 30651
rect 23063 30617 23072 30651
rect 23020 30608 23072 30617
rect 19156 30540 19208 30592
rect 19984 30540 20036 30592
rect 21916 30540 21968 30592
rect 23204 30540 23256 30592
rect 23388 30583 23440 30592
rect 23388 30549 23397 30583
rect 23397 30549 23431 30583
rect 23431 30549 23440 30583
rect 23388 30540 23440 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 19432 30379 19484 30388
rect 19432 30345 19441 30379
rect 19441 30345 19475 30379
rect 19475 30345 19484 30379
rect 19432 30336 19484 30345
rect 22836 30336 22888 30388
rect 25964 30336 26016 30388
rect 19156 30311 19208 30320
rect 19156 30277 19165 30311
rect 19165 30277 19199 30311
rect 19199 30277 19208 30311
rect 19156 30268 19208 30277
rect 9772 30200 9824 30252
rect 18788 30243 18840 30252
rect 18788 30209 18797 30243
rect 18797 30209 18831 30243
rect 18831 30209 18840 30243
rect 18788 30200 18840 30209
rect 18972 30243 19024 30252
rect 18972 30209 18979 30243
rect 18979 30209 19024 30243
rect 18972 30200 19024 30209
rect 19064 30243 19116 30252
rect 19064 30209 19073 30243
rect 19073 30209 19107 30243
rect 19107 30209 19116 30243
rect 19064 30200 19116 30209
rect 19248 30243 19300 30252
rect 19248 30209 19262 30243
rect 19262 30209 19296 30243
rect 19296 30209 19300 30243
rect 19248 30200 19300 30209
rect 940 30132 992 30184
rect 8944 29996 8996 30048
rect 22192 30243 22244 30252
rect 22192 30209 22201 30243
rect 22201 30209 22235 30243
rect 22235 30209 22244 30243
rect 22192 30200 22244 30209
rect 23204 30200 23256 30252
rect 23388 30243 23440 30252
rect 23388 30209 23397 30243
rect 23397 30209 23431 30243
rect 23431 30209 23440 30243
rect 23388 30200 23440 30209
rect 23572 30200 23624 30252
rect 23848 30243 23900 30252
rect 23848 30209 23857 30243
rect 23857 30209 23891 30243
rect 23891 30209 23900 30243
rect 23848 30200 23900 30209
rect 40592 30200 40644 30252
rect 40684 30200 40736 30252
rect 46480 30200 46532 30252
rect 22836 29996 22888 30048
rect 23112 30039 23164 30048
rect 23112 30005 23121 30039
rect 23121 30005 23155 30039
rect 23155 30005 23164 30039
rect 23112 29996 23164 30005
rect 30380 30132 30432 30184
rect 23664 29996 23716 30048
rect 23848 29996 23900 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 6368 29724 6420 29776
rect 27344 29792 27396 29844
rect 18788 29724 18840 29776
rect 24492 29724 24544 29776
rect 19064 29656 19116 29708
rect 22192 29656 22244 29708
rect 1952 29588 2004 29640
rect 23112 29656 23164 29708
rect 23204 29656 23256 29708
rect 25412 29656 25464 29708
rect 22652 29631 22704 29640
rect 22652 29597 22661 29631
rect 22661 29597 22695 29631
rect 22695 29597 22704 29631
rect 22652 29588 22704 29597
rect 22836 29631 22888 29640
rect 22836 29597 22845 29631
rect 22845 29597 22879 29631
rect 22879 29597 22888 29631
rect 22836 29588 22888 29597
rect 940 29520 992 29572
rect 21456 29520 21508 29572
rect 48872 29656 48924 29708
rect 58164 29699 58216 29708
rect 58164 29665 58173 29699
rect 58173 29665 58207 29699
rect 58207 29665 58216 29699
rect 58164 29656 58216 29665
rect 27068 29588 27120 29640
rect 40316 29588 40368 29640
rect 43352 29588 43404 29640
rect 56048 29588 56100 29640
rect 57244 29588 57296 29640
rect 58992 29520 59044 29572
rect 22928 29452 22980 29504
rect 33784 29452 33836 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 9772 29291 9824 29300
rect 9772 29257 9781 29291
rect 9781 29257 9815 29291
rect 9815 29257 9824 29291
rect 9772 29248 9824 29257
rect 19248 29248 19300 29300
rect 24308 29248 24360 29300
rect 9404 29155 9456 29164
rect 9404 29121 9413 29155
rect 9413 29121 9447 29155
rect 9447 29121 9456 29155
rect 9404 29112 9456 29121
rect 19064 29112 19116 29164
rect 24492 28976 24544 29028
rect 30840 28976 30892 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 1676 28636 1728 28688
rect 2596 28636 2648 28688
rect 940 28568 992 28620
rect 9404 28568 9456 28620
rect 2596 28543 2648 28552
rect 2596 28509 2606 28543
rect 2606 28509 2640 28543
rect 2640 28509 2648 28543
rect 21640 28568 21692 28620
rect 2596 28500 2648 28509
rect 54668 28500 54720 28552
rect 28264 28432 28316 28484
rect 49792 28432 49844 28484
rect 58164 28475 58216 28484
rect 58164 28441 58173 28475
rect 58173 28441 58207 28475
rect 58207 28441 58216 28475
rect 58164 28432 58216 28441
rect 25964 28364 26016 28416
rect 47400 28364 47452 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 2320 28024 2372 28076
rect 940 27956 992 28008
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 34244 27548 34296 27600
rect 35440 27548 35492 27600
rect 1584 27455 1636 27464
rect 1584 27421 1593 27455
rect 1593 27421 1627 27455
rect 1627 27421 1636 27455
rect 1584 27412 1636 27421
rect 58992 27412 59044 27464
rect 940 27344 992 27396
rect 34612 27276 34664 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 1584 27072 1636 27124
rect 2412 27004 2464 27056
rect 1676 26936 1728 26988
rect 2504 26979 2556 26988
rect 2504 26945 2513 26979
rect 2513 26945 2547 26979
rect 2547 26945 2556 26979
rect 2504 26936 2556 26945
rect 2596 26979 2648 26988
rect 2596 26945 2606 26979
rect 2606 26945 2640 26979
rect 2640 26945 2648 26979
rect 2596 26936 2648 26945
rect 940 26868 992 26920
rect 2136 26868 2188 26920
rect 21640 27004 21692 27056
rect 7840 26936 7892 26988
rect 23848 27004 23900 27056
rect 23480 26936 23532 26988
rect 23664 26936 23716 26988
rect 23204 26911 23256 26920
rect 23204 26877 23213 26911
rect 23213 26877 23247 26911
rect 23247 26877 23256 26911
rect 23204 26868 23256 26877
rect 24216 26979 24268 26988
rect 24216 26945 24225 26979
rect 24225 26945 24259 26979
rect 24259 26945 24268 26979
rect 24216 26936 24268 26945
rect 24400 26979 24452 26988
rect 24400 26945 24414 26979
rect 24414 26945 24448 26979
rect 24448 26945 24452 26979
rect 27068 27004 27120 27056
rect 24400 26936 24452 26945
rect 26884 26936 26936 26988
rect 27896 26936 27948 26988
rect 24400 26732 24452 26784
rect 30380 26868 30432 26920
rect 55220 26868 55272 26920
rect 48780 26732 48832 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 23664 26571 23716 26580
rect 23664 26537 23673 26571
rect 23673 26537 23707 26571
rect 23707 26537 23716 26571
rect 23664 26528 23716 26537
rect 29000 26392 29052 26444
rect 58164 26435 58216 26444
rect 58164 26401 58173 26435
rect 58173 26401 58207 26435
rect 58207 26401 58216 26435
rect 58164 26392 58216 26401
rect 23388 26367 23440 26376
rect 23388 26333 23397 26367
rect 23397 26333 23431 26367
rect 23431 26333 23440 26367
rect 23388 26324 23440 26333
rect 23572 26324 23624 26376
rect 24124 26324 24176 26376
rect 56324 26324 56376 26376
rect 18512 26256 18564 26308
rect 23940 26256 23992 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 940 25780 992 25832
rect 9404 25848 9456 25900
rect 10692 25891 10744 25900
rect 10692 25857 10701 25891
rect 10701 25857 10735 25891
rect 10735 25857 10744 25891
rect 10692 25848 10744 25857
rect 26884 25848 26936 25900
rect 58072 25891 58124 25900
rect 58072 25857 58081 25891
rect 58081 25857 58115 25891
rect 58115 25857 58124 25891
rect 58072 25848 58124 25857
rect 34060 25780 34112 25832
rect 39304 25780 39356 25832
rect 29000 25712 29052 25764
rect 44732 25712 44784 25764
rect 20628 25644 20680 25696
rect 47032 25644 47084 25696
rect 57980 25644 58032 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2504 25279 2556 25288
rect 2504 25245 2513 25279
rect 2513 25245 2547 25279
rect 2547 25245 2556 25279
rect 2504 25236 2556 25245
rect 2688 25279 2740 25288
rect 2688 25245 2701 25279
rect 2701 25245 2740 25279
rect 2688 25236 2740 25245
rect 52552 25236 52604 25288
rect 940 25168 992 25220
rect 58164 25211 58216 25220
rect 58164 25177 58173 25211
rect 58173 25177 58207 25211
rect 58207 25177 58216 25211
rect 58164 25168 58216 25177
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 47676 24828 47728 24880
rect 48412 24828 48464 24880
rect 2872 24760 2924 24812
rect 58072 24803 58124 24812
rect 58072 24769 58081 24803
rect 58081 24769 58115 24803
rect 58115 24769 58124 24803
rect 58072 24760 58124 24769
rect 940 24692 992 24744
rect 38844 24556 38896 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 2872 24395 2924 24404
rect 2872 24361 2881 24395
rect 2881 24361 2915 24395
rect 2915 24361 2924 24395
rect 2872 24352 2924 24361
rect 24768 24352 24820 24404
rect 42892 24352 42944 24404
rect 2688 24284 2740 24336
rect 17684 24284 17736 24336
rect 18880 24284 18932 24336
rect 39764 24284 39816 24336
rect 7932 24216 7984 24268
rect 31576 24216 31628 24268
rect 36176 24216 36228 24268
rect 54760 24216 54812 24268
rect 940 24080 992 24132
rect 2688 24191 2740 24200
rect 2688 24157 2697 24191
rect 2697 24157 2731 24191
rect 2731 24157 2740 24191
rect 2688 24148 2740 24157
rect 25596 24148 25648 24200
rect 35532 24148 35584 24200
rect 55864 24148 55916 24200
rect 12164 24080 12216 24132
rect 18972 24080 19024 24132
rect 51816 24080 51868 24132
rect 2504 24012 2556 24064
rect 2688 24012 2740 24064
rect 8944 24012 8996 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 19432 23672 19484 23724
rect 12808 23647 12860 23656
rect 12808 23613 12817 23647
rect 12817 23613 12851 23647
rect 12851 23613 12860 23647
rect 12808 23604 12860 23613
rect 23572 23604 23624 23656
rect 24768 23604 24820 23656
rect 19432 23468 19484 23520
rect 20444 23468 20496 23520
rect 27988 23468 28040 23520
rect 34612 23468 34664 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 12164 23307 12216 23316
rect 12164 23273 12173 23307
rect 12173 23273 12207 23307
rect 12207 23273 12216 23307
rect 12164 23264 12216 23273
rect 940 23128 992 23180
rect 10140 23060 10192 23112
rect 10692 23060 10744 23112
rect 12808 23060 12860 23112
rect 25596 23128 25648 23180
rect 29276 23128 29328 23180
rect 58992 23128 59044 23180
rect 24216 23060 24268 23112
rect 25872 23060 25924 23112
rect 57888 23103 57940 23112
rect 57888 23069 57897 23103
rect 57897 23069 57931 23103
rect 57931 23069 57940 23103
rect 57888 23060 57940 23069
rect 22468 22992 22520 23044
rect 33784 22992 33836 23044
rect 20904 22924 20956 22976
rect 39488 22924 39540 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 33784 22720 33836 22772
rect 59176 22720 59228 22772
rect 58164 22695 58216 22704
rect 58164 22661 58173 22695
rect 58173 22661 58207 22695
rect 58207 22661 58216 22695
rect 58164 22652 58216 22661
rect 9772 22584 9824 22636
rect 940 22516 992 22568
rect 18052 22584 18104 22636
rect 18788 22516 18840 22568
rect 16948 22380 17000 22432
rect 41972 22380 42024 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 6828 21972 6880 22024
rect 18880 22176 18932 22228
rect 9772 22083 9824 22092
rect 9772 22049 9781 22083
rect 9781 22049 9815 22083
rect 9815 22049 9824 22083
rect 9772 22040 9824 22049
rect 17960 22151 18012 22160
rect 17960 22117 17969 22151
rect 17969 22117 18003 22151
rect 18003 22117 18012 22151
rect 17960 22108 18012 22117
rect 36636 22108 36688 22160
rect 39580 22108 39632 22160
rect 17316 22040 17368 22092
rect 21364 22040 21416 22092
rect 57060 22040 57112 22092
rect 57428 22040 57480 22092
rect 940 21904 992 21956
rect 10140 21904 10192 21956
rect 17868 21972 17920 22024
rect 17408 21904 17460 21956
rect 21088 21972 21140 22024
rect 57152 21972 57204 22024
rect 18880 21904 18932 21956
rect 22744 21904 22796 21956
rect 23296 21904 23348 21956
rect 58164 21947 58216 21956
rect 58164 21913 58173 21947
rect 58173 21913 58207 21947
rect 58207 21913 58216 21947
rect 58164 21904 58216 21913
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 6828 21632 6880 21684
rect 6092 21496 6144 21548
rect 10140 21496 10192 21548
rect 15660 21564 15712 21616
rect 14096 21496 14148 21548
rect 17868 21564 17920 21616
rect 18236 21564 18288 21616
rect 18328 21539 18380 21548
rect 18328 21505 18337 21539
rect 18337 21505 18371 21539
rect 18371 21505 18380 21539
rect 18328 21496 18380 21505
rect 15384 21428 15436 21480
rect 16396 21360 16448 21412
rect 17408 21471 17460 21480
rect 17408 21437 17417 21471
rect 17417 21437 17451 21471
rect 17451 21437 17460 21471
rect 17408 21428 17460 21437
rect 21640 21632 21692 21684
rect 19616 21496 19668 21548
rect 20904 21564 20956 21616
rect 21824 21564 21876 21616
rect 20260 21496 20312 21548
rect 20812 21496 20864 21548
rect 23572 21539 23624 21548
rect 23572 21505 23581 21539
rect 23581 21505 23615 21539
rect 23615 21505 23624 21539
rect 23572 21496 23624 21505
rect 940 21292 992 21344
rect 13268 21292 13320 21344
rect 16580 21292 16632 21344
rect 16764 21292 16816 21344
rect 18236 21360 18288 21412
rect 19248 21428 19300 21480
rect 25964 21539 26016 21548
rect 25964 21505 25973 21539
rect 25973 21505 26007 21539
rect 26007 21505 26016 21539
rect 25964 21496 26016 21505
rect 28632 21539 28684 21548
rect 28632 21505 28641 21539
rect 28641 21505 28675 21539
rect 28675 21505 28684 21539
rect 28632 21496 28684 21505
rect 34796 21496 34848 21548
rect 21364 21360 21416 21412
rect 28908 21428 28960 21480
rect 19708 21292 19760 21344
rect 20168 21292 20220 21344
rect 20720 21292 20772 21344
rect 26424 21360 26476 21412
rect 39028 21496 39080 21548
rect 43720 21496 43772 21548
rect 58072 21539 58124 21548
rect 58072 21505 58081 21539
rect 58081 21505 58115 21539
rect 58115 21505 58124 21539
rect 58072 21496 58124 21505
rect 39212 21428 39264 21480
rect 42248 21428 42300 21480
rect 42340 21428 42392 21480
rect 57704 21428 57756 21480
rect 57888 21428 57940 21480
rect 23296 21292 23348 21344
rect 40040 21360 40092 21412
rect 33324 21292 33376 21344
rect 38568 21292 38620 21344
rect 42984 21335 43036 21344
rect 42984 21301 42993 21335
rect 42993 21301 43027 21335
rect 43027 21301 43036 21335
rect 42984 21292 43036 21301
rect 49056 21292 49108 21344
rect 57888 21292 57940 21344
rect 58256 21335 58308 21344
rect 58256 21301 58265 21335
rect 58265 21301 58299 21335
rect 58299 21301 58308 21335
rect 58256 21292 58308 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 13176 21088 13228 21140
rect 17316 21088 17368 21140
rect 18236 21088 18288 21140
rect 19616 21131 19668 21140
rect 19616 21097 19625 21131
rect 19625 21097 19659 21131
rect 19659 21097 19668 21131
rect 19616 21088 19668 21097
rect 11888 20884 11940 20936
rect 15200 21020 15252 21072
rect 18144 21020 18196 21072
rect 21088 21131 21140 21140
rect 21088 21097 21097 21131
rect 21097 21097 21131 21131
rect 21131 21097 21140 21131
rect 21088 21088 21140 21097
rect 23572 21088 23624 21140
rect 26148 21088 26200 21140
rect 14280 20927 14332 20936
rect 14280 20893 14289 20927
rect 14289 20893 14323 20927
rect 14323 20893 14332 20927
rect 14280 20884 14332 20893
rect 15384 20927 15436 20936
rect 15384 20893 15393 20927
rect 15393 20893 15427 20927
rect 15427 20893 15436 20927
rect 15384 20884 15436 20893
rect 16212 20816 16264 20868
rect 17224 20884 17276 20936
rect 18144 20927 18196 20936
rect 18144 20893 18153 20927
rect 18153 20893 18187 20927
rect 18187 20893 18196 20927
rect 18144 20884 18196 20893
rect 18788 20884 18840 20936
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 20168 20927 20220 20936
rect 20168 20893 20177 20927
rect 20177 20893 20211 20927
rect 20211 20893 20220 20927
rect 20168 20884 20220 20893
rect 20904 20927 20956 20936
rect 20904 20893 20913 20927
rect 20913 20893 20947 20927
rect 20947 20893 20956 20927
rect 20904 20884 20956 20893
rect 21640 20927 21692 20936
rect 21640 20893 21649 20927
rect 21649 20893 21683 20927
rect 21683 20893 21692 20927
rect 21640 20884 21692 20893
rect 23848 20884 23900 20936
rect 25688 21020 25740 21072
rect 26424 20995 26476 21004
rect 26424 20961 26433 20995
rect 26433 20961 26467 20995
rect 26467 20961 26476 20995
rect 26424 20952 26476 20961
rect 25596 20884 25648 20936
rect 25780 20884 25832 20936
rect 28632 21088 28684 21140
rect 38476 21088 38528 21140
rect 42340 21088 42392 21140
rect 29184 21020 29236 21072
rect 31668 21020 31720 21072
rect 57980 21088 58032 21140
rect 53380 21063 53432 21072
rect 53380 21029 53389 21063
rect 53389 21029 53423 21063
rect 53423 21029 53432 21063
rect 53380 21020 53432 21029
rect 26792 20884 26844 20936
rect 27804 20927 27856 20936
rect 27804 20893 27813 20927
rect 27813 20893 27847 20927
rect 27847 20893 27856 20927
rect 27804 20884 27856 20893
rect 28632 20884 28684 20936
rect 30656 20927 30708 20936
rect 30656 20893 30665 20927
rect 30665 20893 30699 20927
rect 30699 20893 30708 20927
rect 30656 20884 30708 20893
rect 30748 20927 30800 20936
rect 30748 20893 30757 20927
rect 30757 20893 30791 20927
rect 30791 20893 30800 20927
rect 30748 20884 30800 20893
rect 30932 20927 30984 20936
rect 30932 20893 30941 20927
rect 30941 20893 30975 20927
rect 30975 20893 30984 20927
rect 30932 20884 30984 20893
rect 31392 20927 31444 20936
rect 31392 20893 31401 20927
rect 31401 20893 31435 20927
rect 31435 20893 31444 20927
rect 31392 20884 31444 20893
rect 34796 20927 34848 20936
rect 34796 20893 34805 20927
rect 34805 20893 34839 20927
rect 34839 20893 34848 20927
rect 34796 20884 34848 20893
rect 35624 20884 35676 20936
rect 36544 20952 36596 21004
rect 41880 20952 41932 21004
rect 42248 20995 42300 21004
rect 42248 20961 42257 20995
rect 42257 20961 42291 20995
rect 42291 20961 42300 20995
rect 42248 20952 42300 20961
rect 59268 21020 59320 21072
rect 17960 20816 18012 20868
rect 18512 20816 18564 20868
rect 11980 20748 12032 20800
rect 14004 20748 14056 20800
rect 15292 20791 15344 20800
rect 15292 20757 15301 20791
rect 15301 20757 15335 20791
rect 15335 20757 15344 20791
rect 15292 20748 15344 20757
rect 17132 20748 17184 20800
rect 17500 20791 17552 20800
rect 17500 20757 17509 20791
rect 17509 20757 17543 20791
rect 17543 20757 17552 20791
rect 17500 20748 17552 20757
rect 18328 20748 18380 20800
rect 18972 20748 19024 20800
rect 24952 20791 25004 20800
rect 24952 20757 24961 20791
rect 24961 20757 24995 20791
rect 24995 20757 25004 20791
rect 24952 20748 25004 20757
rect 26792 20791 26844 20800
rect 26792 20757 26801 20791
rect 26801 20757 26835 20791
rect 26835 20757 26844 20791
rect 26792 20748 26844 20757
rect 27620 20748 27672 20800
rect 31668 20748 31720 20800
rect 35716 20791 35768 20800
rect 35716 20757 35725 20791
rect 35725 20757 35759 20791
rect 35759 20757 35768 20791
rect 35716 20748 35768 20757
rect 35992 20748 36044 20800
rect 38476 20927 38528 20936
rect 38476 20893 38485 20927
rect 38485 20893 38519 20927
rect 38519 20893 38528 20927
rect 38476 20884 38528 20893
rect 38568 20927 38620 20936
rect 38568 20893 38577 20927
rect 38577 20893 38611 20927
rect 38611 20893 38620 20927
rect 38568 20884 38620 20893
rect 41972 20884 42024 20936
rect 53840 20952 53892 21004
rect 45560 20884 45612 20936
rect 47860 20927 47912 20936
rect 47860 20893 47869 20927
rect 47869 20893 47903 20927
rect 47903 20893 47912 20927
rect 47860 20884 47912 20893
rect 43352 20859 43404 20868
rect 43352 20825 43361 20859
rect 43361 20825 43395 20859
rect 43395 20825 43404 20859
rect 43352 20816 43404 20825
rect 43812 20816 43864 20868
rect 47676 20859 47728 20868
rect 47676 20825 47685 20859
rect 47685 20825 47719 20859
rect 47719 20825 47728 20859
rect 47676 20816 47728 20825
rect 48964 20816 49016 20868
rect 49608 20816 49660 20868
rect 52920 20884 52972 20936
rect 53932 20927 53984 20936
rect 53932 20893 53941 20927
rect 53941 20893 53975 20927
rect 53975 20893 53984 20927
rect 53932 20884 53984 20893
rect 55680 20884 55732 20936
rect 56048 20927 56100 20936
rect 56048 20893 56057 20927
rect 56057 20893 56091 20927
rect 56091 20893 56100 20927
rect 56048 20884 56100 20893
rect 57888 20927 57940 20936
rect 57888 20893 57897 20927
rect 57897 20893 57931 20927
rect 57931 20893 57940 20927
rect 57888 20884 57940 20893
rect 37096 20791 37148 20800
rect 37096 20757 37105 20791
rect 37105 20757 37139 20791
rect 37139 20757 37148 20791
rect 37096 20748 37148 20757
rect 38752 20791 38804 20800
rect 38752 20757 38761 20791
rect 38761 20757 38795 20791
rect 38795 20757 38804 20791
rect 38752 20748 38804 20757
rect 41604 20748 41656 20800
rect 41880 20748 41932 20800
rect 42708 20748 42760 20800
rect 43628 20791 43680 20800
rect 43628 20757 43637 20791
rect 43637 20757 43671 20791
rect 43671 20757 43680 20791
rect 43628 20748 43680 20757
rect 48320 20748 48372 20800
rect 52644 20748 52696 20800
rect 54484 20816 54536 20868
rect 58992 20816 59044 20868
rect 53840 20748 53892 20800
rect 54208 20791 54260 20800
rect 54208 20757 54217 20791
rect 54217 20757 54251 20791
rect 54251 20757 54260 20791
rect 54208 20748 54260 20757
rect 56968 20748 57020 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 16212 20587 16264 20596
rect 16212 20553 16221 20587
rect 16221 20553 16255 20587
rect 16255 20553 16264 20587
rect 16212 20544 16264 20553
rect 18236 20544 18288 20596
rect 19432 20544 19484 20596
rect 11520 20476 11572 20528
rect 15200 20476 15252 20528
rect 3516 20408 3568 20460
rect 9312 20408 9364 20460
rect 10232 20451 10284 20460
rect 10232 20417 10241 20451
rect 10241 20417 10275 20451
rect 10275 20417 10284 20451
rect 10232 20408 10284 20417
rect 940 20340 992 20392
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 13176 20408 13228 20417
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 14004 20451 14056 20460
rect 14004 20417 14013 20451
rect 14013 20417 14047 20451
rect 14047 20417 14056 20451
rect 14004 20408 14056 20417
rect 15292 20451 15344 20460
rect 15292 20417 15301 20451
rect 15301 20417 15335 20451
rect 15335 20417 15344 20451
rect 15292 20408 15344 20417
rect 16948 20476 17000 20528
rect 18512 20519 18564 20528
rect 18512 20485 18521 20519
rect 18521 20485 18555 20519
rect 18555 20485 18564 20519
rect 18512 20476 18564 20485
rect 18972 20519 19024 20528
rect 18972 20485 18981 20519
rect 18981 20485 19015 20519
rect 19015 20485 19024 20519
rect 18972 20476 19024 20485
rect 16856 20451 16908 20460
rect 16856 20417 16865 20451
rect 16865 20417 16899 20451
rect 16899 20417 16908 20451
rect 16856 20408 16908 20417
rect 17132 20451 17184 20460
rect 17132 20417 17141 20451
rect 17141 20417 17175 20451
rect 17175 20417 17184 20451
rect 17132 20408 17184 20417
rect 19156 20408 19208 20460
rect 20168 20476 20220 20528
rect 22468 20587 22520 20596
rect 22468 20553 22477 20587
rect 22477 20553 22511 20587
rect 22511 20553 22520 20587
rect 22468 20544 22520 20553
rect 25596 20587 25648 20596
rect 25596 20553 25605 20587
rect 25605 20553 25639 20587
rect 25639 20553 25648 20587
rect 25596 20544 25648 20553
rect 27804 20544 27856 20596
rect 28448 20544 28500 20596
rect 28908 20544 28960 20596
rect 30748 20544 30800 20596
rect 31024 20587 31076 20596
rect 31024 20553 31033 20587
rect 31033 20553 31067 20587
rect 31067 20553 31076 20587
rect 31024 20544 31076 20553
rect 24952 20476 25004 20528
rect 25136 20476 25188 20528
rect 26792 20476 26844 20528
rect 37096 20544 37148 20596
rect 37280 20544 37332 20596
rect 12900 20340 12952 20392
rect 13084 20383 13136 20392
rect 13084 20349 13093 20383
rect 13093 20349 13127 20383
rect 13127 20349 13136 20383
rect 13084 20340 13136 20349
rect 13728 20340 13780 20392
rect 20904 20340 20956 20392
rect 20996 20383 21048 20392
rect 20996 20349 21005 20383
rect 21005 20349 21039 20383
rect 21039 20349 21048 20383
rect 20996 20340 21048 20349
rect 11704 20272 11756 20324
rect 8116 20204 8168 20256
rect 10324 20204 10376 20256
rect 10968 20204 11020 20256
rect 14188 20247 14240 20256
rect 14188 20213 14197 20247
rect 14197 20213 14231 20247
rect 14231 20213 14240 20247
rect 14188 20204 14240 20213
rect 15476 20247 15528 20256
rect 15476 20213 15485 20247
rect 15485 20213 15519 20247
rect 15519 20213 15528 20247
rect 15476 20204 15528 20213
rect 18880 20272 18932 20324
rect 18788 20204 18840 20256
rect 19248 20204 19300 20256
rect 20536 20272 20588 20324
rect 21732 20272 21784 20324
rect 22100 20408 22152 20460
rect 23848 20408 23900 20460
rect 20352 20204 20404 20256
rect 21364 20247 21416 20256
rect 21364 20213 21373 20247
rect 21373 20213 21407 20247
rect 21407 20213 21416 20247
rect 21364 20204 21416 20213
rect 22836 20204 22888 20256
rect 23204 20204 23256 20256
rect 23388 20340 23440 20392
rect 24860 20204 24912 20256
rect 25136 20247 25188 20256
rect 25136 20213 25145 20247
rect 25145 20213 25179 20247
rect 25179 20213 25188 20247
rect 25136 20204 25188 20213
rect 29000 20408 29052 20460
rect 35716 20476 35768 20528
rect 36084 20476 36136 20528
rect 40040 20587 40092 20596
rect 40040 20553 40049 20587
rect 40049 20553 40083 20587
rect 40083 20553 40092 20587
rect 40040 20544 40092 20553
rect 40684 20544 40736 20596
rect 44456 20544 44508 20596
rect 49608 20587 49660 20596
rect 49608 20553 49617 20587
rect 49617 20553 49651 20587
rect 49651 20553 49660 20587
rect 49608 20544 49660 20553
rect 56324 20587 56376 20596
rect 56324 20553 56333 20587
rect 56333 20553 56367 20587
rect 56367 20553 56376 20587
rect 56324 20544 56376 20553
rect 25504 20340 25556 20392
rect 26516 20340 26568 20392
rect 29092 20340 29144 20392
rect 30196 20408 30248 20460
rect 30656 20408 30708 20460
rect 33416 20451 33468 20460
rect 33416 20417 33425 20451
rect 33425 20417 33459 20451
rect 33459 20417 33468 20451
rect 33416 20408 33468 20417
rect 33600 20451 33652 20460
rect 33600 20417 33609 20451
rect 33609 20417 33643 20451
rect 33643 20417 33652 20451
rect 33600 20408 33652 20417
rect 35900 20408 35952 20460
rect 38752 20451 38804 20460
rect 38752 20417 38761 20451
rect 38761 20417 38795 20451
rect 38795 20417 38804 20451
rect 38752 20408 38804 20417
rect 41604 20451 41656 20460
rect 41604 20417 41613 20451
rect 41613 20417 41647 20451
rect 41647 20417 41656 20451
rect 41604 20408 41656 20417
rect 42800 20451 42852 20460
rect 42800 20417 42809 20451
rect 42809 20417 42843 20451
rect 42843 20417 42852 20451
rect 42800 20408 42852 20417
rect 30748 20340 30800 20392
rect 31116 20383 31168 20392
rect 31116 20349 31125 20383
rect 31125 20349 31159 20383
rect 31159 20349 31168 20383
rect 31116 20340 31168 20349
rect 31484 20340 31536 20392
rect 33324 20340 33376 20392
rect 32864 20272 32916 20324
rect 38384 20340 38436 20392
rect 37188 20272 37240 20324
rect 41696 20340 41748 20392
rect 39672 20272 39724 20324
rect 43720 20451 43772 20460
rect 43720 20417 43729 20451
rect 43729 20417 43763 20451
rect 43763 20417 43772 20451
rect 43720 20408 43772 20417
rect 43904 20451 43956 20460
rect 43904 20417 43913 20451
rect 43913 20417 43947 20451
rect 43947 20417 43956 20451
rect 43904 20408 43956 20417
rect 43996 20451 44048 20460
rect 43996 20417 44005 20451
rect 44005 20417 44039 20451
rect 44039 20417 44048 20451
rect 43996 20408 44048 20417
rect 44732 20476 44784 20528
rect 57704 20476 57756 20528
rect 43352 20340 43404 20392
rect 46756 20408 46808 20460
rect 48504 20451 48556 20460
rect 48504 20417 48538 20451
rect 48538 20417 48556 20451
rect 48504 20408 48556 20417
rect 50160 20408 50212 20460
rect 51632 20451 51684 20460
rect 51632 20417 51641 20451
rect 51641 20417 51675 20451
rect 51675 20417 51684 20451
rect 51632 20408 51684 20417
rect 46940 20340 46992 20392
rect 47676 20340 47728 20392
rect 48228 20383 48280 20392
rect 48228 20349 48237 20383
rect 48237 20349 48271 20383
rect 48271 20349 48280 20383
rect 48228 20340 48280 20349
rect 49240 20340 49292 20392
rect 51448 20383 51500 20392
rect 51448 20349 51457 20383
rect 51457 20349 51491 20383
rect 51491 20349 51500 20383
rect 51448 20340 51500 20349
rect 30748 20204 30800 20256
rect 35992 20204 36044 20256
rect 37096 20204 37148 20256
rect 41788 20247 41840 20256
rect 41788 20213 41797 20247
rect 41797 20213 41831 20247
rect 41831 20213 41840 20247
rect 41788 20204 41840 20213
rect 41880 20204 41932 20256
rect 52368 20272 52420 20324
rect 54208 20408 54260 20460
rect 55036 20408 55088 20460
rect 43996 20204 44048 20256
rect 45376 20204 45428 20256
rect 48412 20204 48464 20256
rect 50528 20204 50580 20256
rect 52460 20204 52512 20256
rect 54484 20315 54536 20324
rect 54484 20281 54493 20315
rect 54493 20281 54527 20315
rect 54527 20281 54536 20315
rect 54484 20272 54536 20281
rect 55864 20204 55916 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 8116 19975 8168 19984
rect 8116 19941 8125 19975
rect 8125 19941 8159 19975
rect 8159 19941 8168 19975
rect 8116 19932 8168 19941
rect 9312 20043 9364 20052
rect 9312 20009 9321 20043
rect 9321 20009 9355 20043
rect 9355 20009 9364 20043
rect 9312 20000 9364 20009
rect 10140 20000 10192 20052
rect 17960 20000 18012 20052
rect 20076 20000 20128 20052
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 7564 19796 7616 19848
rect 11244 19864 11296 19916
rect 11612 19907 11664 19916
rect 11612 19873 11621 19907
rect 11621 19873 11655 19907
rect 11655 19873 11664 19907
rect 11612 19864 11664 19873
rect 11888 19975 11940 19984
rect 11888 19941 11897 19975
rect 11897 19941 11931 19975
rect 11931 19941 11940 19975
rect 11888 19932 11940 19941
rect 13728 19975 13780 19984
rect 13728 19941 13737 19975
rect 13737 19941 13771 19975
rect 13771 19941 13780 19975
rect 13728 19932 13780 19941
rect 16396 19975 16448 19984
rect 16396 19941 16405 19975
rect 16405 19941 16439 19975
rect 16439 19941 16448 19975
rect 16396 19932 16448 19941
rect 20260 19932 20312 19984
rect 8392 19796 8444 19848
rect 9864 19839 9916 19848
rect 9864 19805 9873 19839
rect 9873 19805 9907 19839
rect 9907 19805 9916 19839
rect 9864 19796 9916 19805
rect 11152 19796 11204 19848
rect 11520 19839 11572 19848
rect 11520 19805 11529 19839
rect 11529 19805 11563 19839
rect 11563 19805 11572 19839
rect 11520 19796 11572 19805
rect 12348 19839 12400 19848
rect 12348 19805 12357 19839
rect 12357 19805 12391 19839
rect 12391 19805 12400 19839
rect 12348 19796 12400 19805
rect 16856 19864 16908 19916
rect 20076 19864 20128 19916
rect 23388 20000 23440 20052
rect 21732 19932 21784 19984
rect 24952 20000 25004 20052
rect 25136 20000 25188 20052
rect 26148 20000 26200 20052
rect 31024 20000 31076 20052
rect 42800 20000 42852 20052
rect 23204 19864 23256 19916
rect 13544 19796 13596 19848
rect 940 19728 992 19780
rect 6920 19728 6972 19780
rect 7104 19660 7156 19712
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 14372 19796 14424 19848
rect 17500 19796 17552 19848
rect 20812 19796 20864 19848
rect 21364 19796 21416 19848
rect 21732 19796 21784 19848
rect 24032 19907 24084 19916
rect 24032 19873 24041 19907
rect 24041 19873 24075 19907
rect 24075 19873 24084 19907
rect 24032 19864 24084 19873
rect 24860 19864 24912 19916
rect 25504 19864 25556 19916
rect 15108 19660 15160 19712
rect 15476 19728 15528 19780
rect 15568 19728 15620 19780
rect 19340 19728 19392 19780
rect 21456 19728 21508 19780
rect 24492 19796 24544 19848
rect 25780 19839 25832 19848
rect 25780 19805 25789 19839
rect 25789 19805 25823 19839
rect 25823 19805 25832 19839
rect 25780 19796 25832 19805
rect 42708 19975 42760 19984
rect 42708 19941 42717 19975
rect 42717 19941 42751 19975
rect 42751 19941 42760 19975
rect 43444 20000 43496 20052
rect 44732 20000 44784 20052
rect 47584 20043 47636 20052
rect 47584 20009 47593 20043
rect 47593 20009 47627 20043
rect 47627 20009 47636 20043
rect 47584 20000 47636 20009
rect 48504 20043 48556 20052
rect 48504 20009 48513 20043
rect 48513 20009 48547 20043
rect 48547 20009 48556 20043
rect 48504 20000 48556 20009
rect 50620 20000 50672 20052
rect 42708 19932 42760 19941
rect 24768 19728 24820 19780
rect 27528 19728 27580 19780
rect 15384 19660 15436 19712
rect 18880 19660 18932 19712
rect 19248 19660 19300 19712
rect 21640 19660 21692 19712
rect 22100 19703 22152 19712
rect 22100 19669 22109 19703
rect 22109 19669 22143 19703
rect 22143 19669 22152 19703
rect 22100 19660 22152 19669
rect 25136 19660 25188 19712
rect 27436 19660 27488 19712
rect 27988 19796 28040 19848
rect 28632 19864 28684 19916
rect 32864 19907 32916 19916
rect 30196 19796 30248 19848
rect 30288 19796 30340 19848
rect 32864 19873 32873 19907
rect 32873 19873 32907 19907
rect 32907 19873 32916 19907
rect 32864 19864 32916 19873
rect 37372 19864 37424 19916
rect 33600 19796 33652 19848
rect 37188 19796 37240 19848
rect 30932 19771 30984 19780
rect 30932 19737 30966 19771
rect 30966 19737 30984 19771
rect 30932 19728 30984 19737
rect 36084 19771 36136 19780
rect 36084 19737 36118 19771
rect 36118 19737 36136 19771
rect 36084 19728 36136 19737
rect 28080 19660 28132 19712
rect 33968 19660 34020 19712
rect 34336 19660 34388 19712
rect 36176 19660 36228 19712
rect 36268 19660 36320 19712
rect 40224 19796 40276 19848
rect 42892 19796 42944 19848
rect 45468 19864 45520 19916
rect 48412 19932 48464 19984
rect 49240 19932 49292 19984
rect 53564 20000 53616 20052
rect 53840 20000 53892 20052
rect 55128 20000 55180 20052
rect 56048 20043 56100 20052
rect 56048 20009 56057 20043
rect 56057 20009 56091 20043
rect 56091 20009 56100 20043
rect 56048 20000 56100 20009
rect 54944 19932 54996 19984
rect 48228 19864 48280 19916
rect 45376 19839 45428 19848
rect 45376 19805 45385 19839
rect 45385 19805 45419 19839
rect 45419 19805 45428 19839
rect 45376 19796 45428 19805
rect 46296 19796 46348 19848
rect 48320 19839 48372 19848
rect 48320 19805 48329 19839
rect 48329 19805 48363 19839
rect 48363 19805 48372 19839
rect 48320 19796 48372 19805
rect 52368 19907 52420 19916
rect 52368 19873 52377 19907
rect 52377 19873 52411 19907
rect 52411 19873 52420 19907
rect 52368 19864 52420 19873
rect 52460 19796 52512 19848
rect 54300 19839 54352 19848
rect 54300 19805 54309 19839
rect 54309 19805 54343 19839
rect 54343 19805 54352 19839
rect 54300 19796 54352 19805
rect 56324 19864 56376 19916
rect 55312 19796 55364 19848
rect 55496 19839 55548 19848
rect 55496 19805 55505 19839
rect 55505 19805 55539 19839
rect 55539 19805 55548 19839
rect 55496 19796 55548 19805
rect 40500 19771 40552 19780
rect 38200 19703 38252 19712
rect 38200 19669 38209 19703
rect 38209 19669 38243 19703
rect 38243 19669 38252 19703
rect 38200 19660 38252 19669
rect 40500 19737 40509 19771
rect 40509 19737 40543 19771
rect 40543 19737 40552 19771
rect 40500 19728 40552 19737
rect 40684 19771 40736 19780
rect 40684 19737 40693 19771
rect 40693 19737 40727 19771
rect 40727 19737 40736 19771
rect 40684 19728 40736 19737
rect 41788 19728 41840 19780
rect 42984 19728 43036 19780
rect 50528 19728 50580 19780
rect 45560 19660 45612 19712
rect 45928 19660 45980 19712
rect 52368 19728 52420 19780
rect 55956 19796 56008 19848
rect 56968 19796 57020 19848
rect 54668 19660 54720 19712
rect 54760 19660 54812 19712
rect 55128 19660 55180 19712
rect 57060 19660 57112 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 940 19388 992 19440
rect 7564 19456 7616 19508
rect 9680 19456 9732 19508
rect 10140 19499 10192 19508
rect 10140 19465 10149 19499
rect 10149 19465 10183 19499
rect 10183 19465 10192 19499
rect 10140 19456 10192 19465
rect 11152 19499 11204 19508
rect 11152 19465 11161 19499
rect 11161 19465 11195 19499
rect 11195 19465 11204 19499
rect 11152 19456 11204 19465
rect 6092 19252 6144 19304
rect 7104 19363 7156 19372
rect 7104 19329 7138 19363
rect 7138 19329 7156 19363
rect 7104 19320 7156 19329
rect 10692 19431 10744 19440
rect 10692 19397 10701 19431
rect 10701 19397 10735 19431
rect 10735 19397 10744 19431
rect 10692 19388 10744 19397
rect 11060 19388 11112 19440
rect 12072 19388 12124 19440
rect 12348 19388 12400 19440
rect 10048 19320 10100 19372
rect 11704 19363 11756 19372
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 14188 19320 14240 19372
rect 14372 19363 14424 19372
rect 14372 19329 14381 19363
rect 14381 19329 14415 19363
rect 14415 19329 14424 19363
rect 14372 19320 14424 19329
rect 15568 19388 15620 19440
rect 18144 19456 18196 19508
rect 19156 19456 19208 19508
rect 21640 19456 21692 19508
rect 24768 19499 24820 19508
rect 24768 19465 24777 19499
rect 24777 19465 24811 19499
rect 24811 19465 24820 19499
rect 24768 19456 24820 19465
rect 25596 19456 25648 19508
rect 15200 19320 15252 19372
rect 16580 19320 16632 19372
rect 19156 19363 19208 19372
rect 19156 19329 19165 19363
rect 19165 19329 19199 19363
rect 19199 19329 19208 19363
rect 19156 19320 19208 19329
rect 10968 19227 11020 19236
rect 10968 19193 10977 19227
rect 10977 19193 11011 19227
rect 11011 19193 11020 19227
rect 10968 19184 11020 19193
rect 11428 19184 11480 19236
rect 9680 19116 9732 19168
rect 12808 19116 12860 19168
rect 13360 19116 13412 19168
rect 17040 19295 17092 19304
rect 17040 19261 17049 19295
rect 17049 19261 17083 19295
rect 17083 19261 17092 19295
rect 17040 19252 17092 19261
rect 19340 19252 19392 19304
rect 20076 19363 20128 19372
rect 20076 19329 20085 19363
rect 20085 19329 20119 19363
rect 20119 19329 20128 19363
rect 20076 19320 20128 19329
rect 20168 19320 20220 19372
rect 20904 19320 20956 19372
rect 21180 19320 21232 19372
rect 22100 19320 22152 19372
rect 23388 19363 23440 19372
rect 23388 19329 23397 19363
rect 23397 19329 23431 19363
rect 23431 19329 23440 19363
rect 26516 19388 26568 19440
rect 23388 19320 23440 19329
rect 25136 19320 25188 19372
rect 25596 19363 25648 19372
rect 25596 19329 25605 19363
rect 25605 19329 25639 19363
rect 25639 19329 25648 19363
rect 25596 19320 25648 19329
rect 25780 19320 25832 19372
rect 25964 19320 26016 19372
rect 26148 19320 26200 19372
rect 27528 19388 27580 19440
rect 30288 19363 30340 19372
rect 30288 19329 30297 19363
rect 30297 19329 30331 19363
rect 30331 19329 30340 19363
rect 30288 19320 30340 19329
rect 30564 19363 30616 19372
rect 30564 19329 30598 19363
rect 30598 19329 30616 19363
rect 30564 19320 30616 19329
rect 31668 19499 31720 19508
rect 31668 19465 31677 19499
rect 31677 19465 31711 19499
rect 31711 19465 31720 19499
rect 31668 19456 31720 19465
rect 33416 19456 33468 19508
rect 33968 19499 34020 19508
rect 33968 19465 33977 19499
rect 33977 19465 34011 19499
rect 34011 19465 34020 19499
rect 33968 19456 34020 19465
rect 34060 19499 34112 19508
rect 34060 19465 34069 19499
rect 34069 19465 34103 19499
rect 34103 19465 34112 19499
rect 34060 19456 34112 19465
rect 35900 19499 35952 19508
rect 35900 19465 35909 19499
rect 35909 19465 35943 19499
rect 35943 19465 35952 19499
rect 35900 19456 35952 19465
rect 40500 19456 40552 19508
rect 41328 19456 41380 19508
rect 31392 19388 31444 19440
rect 36268 19431 36320 19440
rect 36268 19397 36277 19431
rect 36277 19397 36311 19431
rect 36311 19397 36320 19431
rect 36268 19388 36320 19397
rect 43352 19456 43404 19508
rect 45928 19456 45980 19508
rect 46848 19499 46900 19508
rect 46848 19465 46857 19499
rect 46857 19465 46891 19499
rect 46891 19465 46900 19499
rect 46848 19456 46900 19465
rect 46940 19456 46992 19508
rect 49700 19456 49752 19508
rect 43628 19388 43680 19440
rect 47860 19388 47912 19440
rect 48136 19388 48188 19440
rect 32496 19320 32548 19372
rect 33968 19320 34020 19372
rect 36360 19363 36412 19372
rect 36360 19329 36369 19363
rect 36369 19329 36403 19363
rect 36403 19329 36412 19363
rect 36360 19320 36412 19329
rect 21364 19252 21416 19304
rect 22468 19252 22520 19304
rect 25412 19252 25464 19304
rect 36544 19295 36596 19304
rect 36544 19261 36553 19295
rect 36553 19261 36587 19295
rect 36587 19261 36596 19295
rect 39212 19320 39264 19372
rect 41696 19363 41748 19372
rect 41696 19329 41705 19363
rect 41705 19329 41739 19363
rect 41739 19329 41748 19363
rect 41696 19320 41748 19329
rect 41880 19363 41932 19372
rect 41880 19329 41889 19363
rect 41889 19329 41923 19363
rect 41923 19329 41932 19363
rect 41880 19320 41932 19329
rect 42892 19363 42944 19372
rect 42892 19329 42901 19363
rect 42901 19329 42935 19363
rect 42935 19329 42944 19363
rect 42892 19320 42944 19329
rect 45468 19363 45520 19372
rect 45468 19329 45477 19363
rect 45477 19329 45511 19363
rect 45511 19329 45520 19363
rect 45468 19320 45520 19329
rect 45744 19363 45796 19372
rect 45744 19329 45778 19363
rect 45778 19329 45796 19363
rect 45744 19320 45796 19329
rect 47676 19320 47728 19372
rect 49792 19363 49844 19372
rect 49792 19329 49801 19363
rect 49801 19329 49835 19363
rect 49835 19329 49844 19363
rect 49792 19320 49844 19329
rect 51632 19499 51684 19508
rect 51632 19465 51641 19499
rect 51641 19465 51675 19499
rect 51675 19465 51684 19499
rect 51632 19456 51684 19465
rect 55036 19456 55088 19508
rect 50528 19388 50580 19440
rect 51264 19431 51316 19440
rect 51264 19397 51273 19431
rect 51273 19397 51307 19431
rect 51307 19397 51316 19431
rect 51264 19388 51316 19397
rect 53564 19388 53616 19440
rect 36544 19252 36596 19261
rect 18328 19184 18380 19236
rect 13912 19116 13964 19168
rect 17316 19116 17368 19168
rect 19892 19116 19944 19168
rect 21916 19184 21968 19236
rect 21088 19116 21140 19168
rect 21180 19116 21232 19168
rect 21548 19116 21600 19168
rect 27436 19184 27488 19236
rect 24492 19116 24544 19168
rect 25228 19116 25280 19168
rect 25780 19159 25832 19168
rect 25780 19125 25789 19159
rect 25789 19125 25823 19159
rect 25823 19125 25832 19159
rect 25780 19116 25832 19125
rect 28080 19116 28132 19168
rect 29276 19116 29328 19168
rect 40040 19252 40092 19304
rect 40500 19252 40552 19304
rect 42340 19252 42392 19304
rect 50620 19252 50672 19304
rect 50988 19252 51040 19304
rect 54760 19363 54812 19372
rect 54760 19329 54769 19363
rect 54769 19329 54803 19363
rect 54803 19329 54812 19363
rect 54760 19320 54812 19329
rect 37832 19116 37884 19168
rect 40960 19116 41012 19168
rect 49700 19184 49752 19236
rect 51448 19184 51500 19236
rect 55496 19184 55548 19236
rect 55680 19184 55732 19236
rect 50160 19116 50212 19168
rect 50436 19116 50488 19168
rect 58624 19116 58676 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 8392 18912 8444 18964
rect 9036 18844 9088 18896
rect 9588 18912 9640 18964
rect 10232 18912 10284 18964
rect 11612 18912 11664 18964
rect 13912 18912 13964 18964
rect 16580 18955 16632 18964
rect 16580 18921 16589 18955
rect 16589 18921 16623 18955
rect 16623 18921 16632 18955
rect 16580 18912 16632 18921
rect 18788 18955 18840 18964
rect 18788 18921 18797 18955
rect 18797 18921 18831 18955
rect 18831 18921 18840 18955
rect 18788 18912 18840 18921
rect 20904 18912 20956 18964
rect 21088 18912 21140 18964
rect 9312 18844 9364 18896
rect 11888 18844 11940 18896
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 5264 18708 5316 18760
rect 7104 18708 7156 18760
rect 940 18640 992 18692
rect 6736 18640 6788 18692
rect 6920 18640 6972 18692
rect 10232 18819 10284 18828
rect 10232 18785 10241 18819
rect 10241 18785 10275 18819
rect 10275 18785 10284 18819
rect 10232 18776 10284 18785
rect 12072 18819 12124 18828
rect 12072 18785 12081 18819
rect 12081 18785 12115 18819
rect 12115 18785 12124 18819
rect 12072 18776 12124 18785
rect 8208 18751 8260 18760
rect 8208 18717 8217 18751
rect 8217 18717 8251 18751
rect 8251 18717 8260 18751
rect 8208 18708 8260 18717
rect 8392 18751 8444 18760
rect 8392 18717 8401 18751
rect 8401 18717 8435 18751
rect 8435 18717 8444 18751
rect 8392 18708 8444 18717
rect 10140 18708 10192 18760
rect 10048 18640 10100 18692
rect 11428 18751 11480 18760
rect 11428 18717 11437 18751
rect 11437 18717 11471 18751
rect 11471 18717 11480 18751
rect 11428 18708 11480 18717
rect 13176 18708 13228 18760
rect 14832 18819 14884 18828
rect 14832 18785 14841 18819
rect 14841 18785 14875 18819
rect 14875 18785 14884 18819
rect 14832 18776 14884 18785
rect 15568 18708 15620 18760
rect 25780 18912 25832 18964
rect 5724 18572 5776 18624
rect 8392 18572 8444 18624
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9312 18572 9364 18581
rect 9956 18572 10008 18624
rect 10692 18572 10744 18624
rect 12164 18640 12216 18692
rect 15476 18640 15528 18692
rect 13176 18572 13228 18624
rect 16948 18708 17000 18760
rect 18512 18708 18564 18760
rect 24676 18887 24728 18896
rect 24676 18853 24685 18887
rect 24685 18853 24719 18887
rect 24719 18853 24728 18887
rect 24676 18844 24728 18853
rect 20352 18776 20404 18828
rect 22652 18776 22704 18828
rect 19340 18640 19392 18692
rect 20720 18708 20772 18760
rect 21364 18751 21416 18760
rect 21364 18717 21373 18751
rect 21373 18717 21407 18751
rect 21407 18717 21416 18751
rect 21364 18708 21416 18717
rect 23204 18708 23256 18760
rect 25688 18708 25740 18760
rect 29184 18912 29236 18964
rect 30564 18912 30616 18964
rect 43720 18912 43772 18964
rect 43904 18912 43956 18964
rect 45744 18912 45796 18964
rect 46296 18912 46348 18964
rect 48504 18912 48556 18964
rect 50528 18912 50580 18964
rect 54300 18844 54352 18896
rect 26516 18819 26568 18828
rect 26516 18785 26525 18819
rect 26525 18785 26559 18819
rect 26559 18785 26568 18819
rect 26516 18776 26568 18785
rect 27528 18776 27580 18828
rect 29460 18776 29512 18828
rect 29736 18776 29788 18828
rect 27804 18708 27856 18760
rect 28448 18708 28500 18760
rect 28816 18751 28868 18760
rect 28816 18717 28819 18751
rect 28819 18717 28868 18751
rect 28816 18708 28868 18717
rect 30196 18751 30248 18760
rect 30196 18717 30205 18751
rect 30205 18717 30239 18751
rect 30239 18717 30248 18751
rect 30196 18708 30248 18717
rect 20168 18640 20220 18692
rect 17960 18572 18012 18624
rect 19248 18572 19300 18624
rect 21180 18572 21232 18624
rect 24952 18683 25004 18692
rect 24952 18649 24961 18683
rect 24961 18649 24995 18683
rect 24995 18649 25004 18683
rect 24952 18640 25004 18649
rect 25228 18683 25280 18692
rect 25228 18649 25237 18683
rect 25237 18649 25271 18683
rect 25271 18649 25280 18683
rect 25228 18640 25280 18649
rect 24860 18572 24912 18624
rect 27252 18640 27304 18692
rect 27712 18572 27764 18624
rect 28540 18683 28592 18692
rect 28540 18649 28549 18683
rect 28549 18649 28583 18683
rect 28583 18649 28592 18683
rect 28540 18640 28592 18649
rect 30012 18572 30064 18624
rect 30748 18776 30800 18828
rect 31392 18819 31444 18828
rect 31392 18785 31401 18819
rect 31401 18785 31435 18819
rect 31435 18785 31444 18819
rect 31392 18776 31444 18785
rect 31484 18819 31536 18828
rect 31484 18785 31493 18819
rect 31493 18785 31527 18819
rect 31527 18785 31536 18819
rect 31484 18776 31536 18785
rect 37372 18819 37424 18828
rect 37372 18785 37381 18819
rect 37381 18785 37415 18819
rect 37415 18785 37424 18819
rect 37372 18776 37424 18785
rect 40500 18776 40552 18828
rect 41236 18819 41288 18828
rect 41236 18785 41245 18819
rect 41245 18785 41279 18819
rect 41279 18785 41288 18819
rect 41236 18776 41288 18785
rect 31668 18708 31720 18760
rect 32404 18751 32456 18760
rect 32404 18717 32413 18751
rect 32413 18717 32447 18751
rect 32447 18717 32456 18751
rect 32404 18708 32456 18717
rect 37096 18751 37148 18760
rect 37096 18717 37105 18751
rect 37105 18717 37139 18751
rect 37139 18717 37148 18751
rect 37096 18708 37148 18717
rect 38844 18708 38896 18760
rect 40960 18751 41012 18760
rect 40960 18717 40969 18751
rect 40969 18717 41003 18751
rect 41003 18717 41012 18751
rect 40960 18708 41012 18717
rect 32956 18640 33008 18692
rect 42524 18751 42576 18760
rect 42524 18717 42533 18751
rect 42533 18717 42567 18751
rect 42567 18717 42576 18751
rect 42524 18708 42576 18717
rect 37096 18572 37148 18624
rect 39120 18615 39172 18624
rect 39120 18581 39129 18615
rect 39129 18581 39163 18615
rect 39163 18581 39172 18615
rect 39120 18572 39172 18581
rect 40500 18572 40552 18624
rect 41144 18572 41196 18624
rect 42708 18708 42760 18760
rect 43720 18708 43772 18760
rect 42800 18683 42852 18692
rect 42800 18649 42809 18683
rect 42809 18649 42843 18683
rect 42843 18649 42852 18683
rect 42800 18640 42852 18649
rect 42892 18683 42944 18692
rect 42892 18649 42901 18683
rect 42901 18649 42935 18683
rect 42935 18649 42944 18683
rect 42892 18640 42944 18649
rect 43628 18683 43680 18692
rect 43628 18649 43637 18683
rect 43637 18649 43671 18683
rect 43671 18649 43680 18683
rect 43628 18640 43680 18649
rect 45376 18751 45428 18760
rect 45376 18717 45385 18751
rect 45385 18717 45419 18751
rect 45419 18717 45428 18751
rect 45376 18708 45428 18717
rect 46020 18708 46072 18760
rect 49792 18776 49844 18828
rect 55496 18819 55548 18828
rect 55496 18785 55505 18819
rect 55505 18785 55539 18819
rect 55539 18785 55548 18819
rect 55496 18776 55548 18785
rect 46572 18708 46624 18760
rect 46664 18708 46716 18760
rect 48412 18708 48464 18760
rect 48688 18751 48740 18760
rect 48688 18717 48697 18751
rect 48697 18717 48731 18751
rect 48731 18717 48740 18751
rect 48688 18708 48740 18717
rect 55680 18751 55732 18760
rect 55680 18717 55689 18751
rect 55689 18717 55723 18751
rect 55723 18717 55732 18751
rect 55680 18708 55732 18717
rect 42708 18572 42760 18624
rect 43168 18615 43220 18624
rect 43168 18581 43177 18615
rect 43177 18581 43211 18615
rect 43211 18581 43220 18615
rect 43168 18572 43220 18581
rect 43444 18572 43496 18624
rect 46112 18572 46164 18624
rect 47584 18640 47636 18692
rect 47768 18640 47820 18692
rect 50068 18640 50120 18692
rect 52368 18640 52420 18692
rect 58992 18708 59044 18760
rect 46940 18572 46992 18624
rect 47676 18572 47728 18624
rect 48964 18572 49016 18624
rect 56140 18572 56192 18624
rect 58072 18615 58124 18624
rect 58072 18581 58081 18615
rect 58081 18581 58115 18615
rect 58115 18581 58124 18615
rect 58072 18572 58124 18581
rect 58992 18572 59044 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 8116 18368 8168 18420
rect 6092 18300 6144 18352
rect 9864 18368 9916 18420
rect 12164 18411 12216 18420
rect 12164 18377 12173 18411
rect 12173 18377 12207 18411
rect 12207 18377 12216 18411
rect 12164 18368 12216 18377
rect 5724 18275 5776 18284
rect 5724 18241 5733 18275
rect 5733 18241 5767 18275
rect 5767 18241 5776 18275
rect 5724 18232 5776 18241
rect 9956 18300 10008 18352
rect 10140 18300 10192 18352
rect 15476 18368 15528 18420
rect 16396 18368 16448 18420
rect 18328 18368 18380 18420
rect 25596 18368 25648 18420
rect 25688 18368 25740 18420
rect 27252 18411 27304 18420
rect 27252 18377 27261 18411
rect 27261 18377 27295 18411
rect 27295 18377 27304 18411
rect 27252 18368 27304 18377
rect 27620 18411 27672 18420
rect 27620 18377 27629 18411
rect 27629 18377 27663 18411
rect 27663 18377 27672 18411
rect 27620 18368 27672 18377
rect 29736 18368 29788 18420
rect 13360 18300 13412 18352
rect 6920 18164 6972 18216
rect 7104 18207 7156 18216
rect 7104 18173 7113 18207
rect 7113 18173 7147 18207
rect 7147 18173 7156 18207
rect 7104 18164 7156 18173
rect 9680 18232 9732 18284
rect 10324 18275 10376 18284
rect 10324 18241 10333 18275
rect 10333 18241 10367 18275
rect 10367 18241 10376 18275
rect 10324 18232 10376 18241
rect 11980 18275 12032 18284
rect 11980 18241 11989 18275
rect 11989 18241 12023 18275
rect 12023 18241 12032 18275
rect 11980 18232 12032 18241
rect 12900 18275 12952 18284
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 13176 18232 13228 18284
rect 13268 18275 13320 18284
rect 13268 18241 13277 18275
rect 13277 18241 13311 18275
rect 13311 18241 13320 18275
rect 13268 18232 13320 18241
rect 8484 18207 8536 18216
rect 8484 18173 8493 18207
rect 8493 18173 8527 18207
rect 8527 18173 8536 18207
rect 8484 18164 8536 18173
rect 9312 18164 9364 18216
rect 14464 18275 14516 18284
rect 14464 18241 14473 18275
rect 14473 18241 14507 18275
rect 14507 18241 14516 18275
rect 14464 18232 14516 18241
rect 17040 18232 17092 18284
rect 17960 18232 18012 18284
rect 19524 18275 19576 18284
rect 19524 18241 19533 18275
rect 19533 18241 19567 18275
rect 19567 18241 19576 18275
rect 19524 18232 19576 18241
rect 16764 18164 16816 18216
rect 19616 18164 19668 18216
rect 20168 18164 20220 18216
rect 21548 18300 21600 18352
rect 20720 18232 20772 18284
rect 21640 18232 21692 18284
rect 22100 18232 22152 18284
rect 24216 18232 24268 18284
rect 25596 18232 25648 18284
rect 28080 18232 28132 18284
rect 29460 18275 29512 18284
rect 29460 18241 29469 18275
rect 29469 18241 29503 18275
rect 29503 18241 29512 18275
rect 29460 18232 29512 18241
rect 29552 18275 29604 18284
rect 29552 18241 29561 18275
rect 29561 18241 29595 18275
rect 29595 18241 29604 18275
rect 29552 18232 29604 18241
rect 29736 18275 29788 18284
rect 29736 18241 29745 18275
rect 29745 18241 29779 18275
rect 29779 18241 29788 18275
rect 29736 18232 29788 18241
rect 43168 18368 43220 18420
rect 46020 18368 46072 18420
rect 48320 18368 48372 18420
rect 12624 18096 12676 18148
rect 14096 18096 14148 18148
rect 14556 18096 14608 18148
rect 6552 18028 6604 18080
rect 9588 18028 9640 18080
rect 14464 18028 14516 18080
rect 15292 18028 15344 18080
rect 18512 18096 18564 18148
rect 21916 18164 21968 18216
rect 26148 18164 26200 18216
rect 27712 18207 27764 18216
rect 27712 18173 27721 18207
rect 27721 18173 27755 18207
rect 27755 18173 27764 18207
rect 27712 18164 27764 18173
rect 24308 18096 24360 18148
rect 24492 18139 24544 18148
rect 24492 18105 24501 18139
rect 24501 18105 24535 18139
rect 24535 18105 24544 18139
rect 24492 18096 24544 18105
rect 25136 18096 25188 18148
rect 25964 18096 26016 18148
rect 19248 18028 19300 18080
rect 19340 18028 19392 18080
rect 20260 18028 20312 18080
rect 20720 18028 20772 18080
rect 22652 18028 22704 18080
rect 27712 18028 27764 18080
rect 30012 18232 30064 18284
rect 32220 18300 32272 18352
rect 32404 18300 32456 18352
rect 30748 18207 30800 18216
rect 30748 18173 30757 18207
rect 30757 18173 30791 18207
rect 30791 18173 30800 18207
rect 30748 18164 30800 18173
rect 32956 18232 33008 18284
rect 34060 18300 34112 18352
rect 41236 18300 41288 18352
rect 41512 18300 41564 18352
rect 38660 18232 38712 18284
rect 32404 18164 32456 18216
rect 32588 18207 32640 18216
rect 32588 18173 32597 18207
rect 32597 18173 32631 18207
rect 32631 18173 32640 18207
rect 32588 18164 32640 18173
rect 32680 18207 32732 18216
rect 32680 18173 32689 18207
rect 32689 18173 32723 18207
rect 32723 18173 32732 18207
rect 32680 18164 32732 18173
rect 32772 18207 32824 18216
rect 32772 18173 32781 18207
rect 32781 18173 32815 18207
rect 32815 18173 32824 18207
rect 32772 18164 32824 18173
rect 33876 18164 33928 18216
rect 35348 18164 35400 18216
rect 38844 18207 38896 18216
rect 38844 18173 38853 18207
rect 38853 18173 38887 18207
rect 38887 18173 38896 18207
rect 38844 18164 38896 18173
rect 39120 18275 39172 18284
rect 39120 18241 39129 18275
rect 39129 18241 39163 18275
rect 39163 18241 39172 18275
rect 39120 18232 39172 18241
rect 42432 18232 42484 18284
rect 40960 18164 41012 18216
rect 42892 18343 42944 18352
rect 42892 18309 42901 18343
rect 42901 18309 42935 18343
rect 42935 18309 42944 18343
rect 42892 18300 42944 18309
rect 43628 18300 43680 18352
rect 44732 18300 44784 18352
rect 46112 18343 46164 18352
rect 46112 18309 46121 18343
rect 46121 18309 46155 18343
rect 46155 18309 46164 18343
rect 46112 18300 46164 18309
rect 46848 18300 46900 18352
rect 42984 18275 43036 18284
rect 42984 18241 42993 18275
rect 42993 18241 43027 18275
rect 43027 18241 43036 18275
rect 42984 18232 43036 18241
rect 44180 18232 44232 18284
rect 42892 18164 42944 18216
rect 47124 18232 47176 18284
rect 48504 18232 48556 18284
rect 49976 18368 50028 18420
rect 55680 18368 55732 18420
rect 57244 18411 57296 18420
rect 57244 18377 57253 18411
rect 57253 18377 57287 18411
rect 57287 18377 57296 18411
rect 57244 18368 57296 18377
rect 58716 18368 58768 18420
rect 56140 18343 56192 18352
rect 56140 18309 56174 18343
rect 56174 18309 56192 18343
rect 56140 18300 56192 18309
rect 48964 18275 49016 18284
rect 46572 18164 46624 18216
rect 48136 18164 48188 18216
rect 48964 18241 48998 18275
rect 48998 18241 49016 18275
rect 48964 18232 49016 18241
rect 54576 18275 54628 18284
rect 54576 18241 54585 18275
rect 54585 18241 54619 18275
rect 54619 18241 54628 18275
rect 54576 18232 54628 18241
rect 54760 18275 54812 18284
rect 54760 18241 54769 18275
rect 54769 18241 54803 18275
rect 54803 18241 54812 18275
rect 54760 18232 54812 18241
rect 54944 18275 54996 18284
rect 54944 18241 54953 18275
rect 54953 18241 54987 18275
rect 54987 18241 54996 18275
rect 54944 18232 54996 18241
rect 55864 18207 55916 18216
rect 55864 18173 55873 18207
rect 55873 18173 55907 18207
rect 55907 18173 55916 18207
rect 55864 18164 55916 18173
rect 28080 18028 28132 18080
rect 32220 18028 32272 18080
rect 32680 18028 32732 18080
rect 33968 18071 34020 18080
rect 33968 18037 33977 18071
rect 33977 18037 34011 18071
rect 34011 18037 34020 18071
rect 33968 18028 34020 18037
rect 42432 18028 42484 18080
rect 42524 18028 42576 18080
rect 58716 18096 58768 18148
rect 43444 18028 43496 18080
rect 52092 18028 52144 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 5264 17824 5316 17876
rect 10232 17824 10284 17876
rect 10324 17824 10376 17876
rect 13268 17824 13320 17876
rect 14280 17824 14332 17876
rect 15200 17824 15252 17876
rect 16764 17867 16816 17876
rect 16764 17833 16773 17867
rect 16773 17833 16807 17867
rect 16807 17833 16816 17867
rect 16764 17824 16816 17833
rect 16948 17824 17000 17876
rect 18696 17824 18748 17876
rect 24492 17824 24544 17876
rect 24952 17824 25004 17876
rect 23664 17756 23716 17808
rect 940 17688 992 17740
rect 8116 17731 8168 17740
rect 8116 17697 8125 17731
rect 8125 17697 8159 17731
rect 8159 17697 8168 17731
rect 8116 17688 8168 17697
rect 6460 17620 6512 17672
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 6552 17620 6604 17629
rect 9956 17688 10008 17740
rect 10324 17688 10376 17740
rect 10048 17663 10100 17672
rect 10048 17629 10057 17663
rect 10057 17629 10091 17663
rect 10091 17629 10100 17663
rect 10048 17620 10100 17629
rect 14832 17620 14884 17672
rect 15108 17663 15160 17672
rect 15108 17629 15117 17663
rect 15117 17629 15151 17663
rect 15151 17629 15160 17663
rect 15108 17620 15160 17629
rect 18696 17688 18748 17740
rect 18788 17688 18840 17740
rect 16212 17620 16264 17672
rect 6736 17527 6788 17536
rect 6736 17493 6745 17527
rect 6745 17493 6779 17527
rect 6779 17493 6788 17527
rect 6736 17484 6788 17493
rect 8576 17484 8628 17536
rect 17776 17484 17828 17536
rect 18052 17620 18104 17672
rect 19432 17663 19484 17672
rect 19432 17629 19441 17663
rect 19441 17629 19475 17663
rect 19475 17629 19484 17663
rect 19432 17620 19484 17629
rect 19616 17663 19668 17672
rect 19616 17629 19625 17663
rect 19625 17629 19659 17663
rect 19659 17629 19668 17663
rect 19616 17620 19668 17629
rect 23296 17688 23348 17740
rect 20904 17663 20956 17672
rect 20904 17629 20913 17663
rect 20913 17629 20947 17663
rect 20947 17629 20956 17663
rect 20904 17620 20956 17629
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 28540 17756 28592 17808
rect 24216 17688 24268 17740
rect 18144 17552 18196 17604
rect 18696 17484 18748 17536
rect 20444 17552 20496 17604
rect 23940 17620 23992 17672
rect 21548 17552 21600 17604
rect 24308 17552 24360 17604
rect 25596 17731 25648 17740
rect 25596 17697 25605 17731
rect 25605 17697 25639 17731
rect 25639 17697 25648 17731
rect 25596 17688 25648 17697
rect 27068 17663 27120 17672
rect 27068 17629 27077 17663
rect 27077 17629 27111 17663
rect 27111 17629 27120 17663
rect 27068 17620 27120 17629
rect 27344 17663 27396 17672
rect 27344 17629 27353 17663
rect 27353 17629 27387 17663
rect 27387 17629 27396 17663
rect 27344 17620 27396 17629
rect 27896 17688 27948 17740
rect 25044 17552 25096 17604
rect 21088 17484 21140 17536
rect 24676 17527 24728 17536
rect 24676 17493 24685 17527
rect 24685 17493 24719 17527
rect 24719 17493 24728 17527
rect 24676 17484 24728 17493
rect 24860 17527 24912 17536
rect 24860 17493 24869 17527
rect 24869 17493 24903 17527
rect 24903 17493 24912 17527
rect 24860 17484 24912 17493
rect 25228 17484 25280 17536
rect 25412 17484 25464 17536
rect 27160 17484 27212 17536
rect 27344 17484 27396 17536
rect 27988 17620 28040 17672
rect 28356 17663 28408 17672
rect 28356 17629 28363 17663
rect 28363 17629 28408 17663
rect 28356 17620 28408 17629
rect 29828 17799 29880 17808
rect 29828 17765 29837 17799
rect 29837 17765 29871 17799
rect 29871 17765 29880 17799
rect 29828 17756 29880 17765
rect 32772 17824 32824 17876
rect 37188 17824 37240 17876
rect 38844 17824 38896 17876
rect 38936 17824 38988 17876
rect 31024 17688 31076 17740
rect 28724 17484 28776 17536
rect 30012 17663 30064 17672
rect 30012 17629 30021 17663
rect 30021 17629 30055 17663
rect 30055 17629 30064 17663
rect 30012 17620 30064 17629
rect 28908 17552 28960 17604
rect 31944 17620 31996 17672
rect 32496 17731 32548 17740
rect 32496 17697 32505 17731
rect 32505 17697 32539 17731
rect 32539 17697 32548 17731
rect 32496 17688 32548 17697
rect 33876 17688 33928 17740
rect 34060 17731 34112 17740
rect 34060 17697 34069 17731
rect 34069 17697 34103 17731
rect 34103 17697 34112 17731
rect 34060 17688 34112 17697
rect 33784 17663 33836 17672
rect 33784 17629 33793 17663
rect 33793 17629 33827 17663
rect 33827 17629 33836 17663
rect 33784 17620 33836 17629
rect 34796 17620 34848 17672
rect 38752 17799 38804 17808
rect 38752 17765 38761 17799
rect 38761 17765 38795 17799
rect 38795 17765 38804 17799
rect 38752 17756 38804 17765
rect 41236 17756 41288 17808
rect 48688 17756 48740 17808
rect 53012 17867 53064 17876
rect 53012 17833 53021 17867
rect 53021 17833 53055 17867
rect 53055 17833 53064 17867
rect 53012 17824 53064 17833
rect 54484 17824 54536 17876
rect 57152 17824 57204 17876
rect 39212 17688 39264 17740
rect 39856 17688 39908 17740
rect 40224 17731 40276 17740
rect 40224 17697 40233 17731
rect 40233 17697 40267 17731
rect 40267 17697 40276 17731
rect 40224 17688 40276 17697
rect 48136 17688 48188 17740
rect 40500 17663 40552 17672
rect 30288 17484 30340 17536
rect 31392 17484 31444 17536
rect 33692 17552 33744 17604
rect 32772 17484 32824 17536
rect 33232 17484 33284 17536
rect 33876 17527 33928 17536
rect 33876 17493 33885 17527
rect 33885 17493 33919 17527
rect 33919 17493 33928 17527
rect 33876 17484 33928 17493
rect 36912 17552 36964 17604
rect 38660 17552 38712 17604
rect 39212 17595 39264 17604
rect 39212 17561 39221 17595
rect 39221 17561 39255 17595
rect 39255 17561 39264 17595
rect 39212 17552 39264 17561
rect 40500 17629 40534 17663
rect 40534 17629 40552 17663
rect 40500 17620 40552 17629
rect 47952 17663 48004 17672
rect 47952 17629 47961 17663
rect 47961 17629 47995 17663
rect 47995 17629 48004 17663
rect 47952 17620 48004 17629
rect 38936 17484 38988 17536
rect 46940 17552 46992 17604
rect 49976 17552 50028 17604
rect 50988 17663 51040 17672
rect 50988 17629 50997 17663
rect 50997 17629 51031 17663
rect 51031 17629 51040 17663
rect 50988 17620 51040 17629
rect 51632 17663 51684 17672
rect 51632 17629 51641 17663
rect 51641 17629 51675 17663
rect 51675 17629 51684 17663
rect 51632 17620 51684 17629
rect 54760 17688 54812 17740
rect 53012 17620 53064 17672
rect 53840 17620 53892 17672
rect 55864 17688 55916 17740
rect 58256 17620 58308 17672
rect 51908 17595 51960 17604
rect 51908 17561 51942 17595
rect 51942 17561 51960 17595
rect 51908 17552 51960 17561
rect 56324 17552 56376 17604
rect 51080 17484 51132 17536
rect 51632 17484 51684 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 8484 17280 8536 17332
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 6460 17212 6512 17264
rect 11152 17212 11204 17264
rect 17960 17323 18012 17332
rect 17960 17289 17969 17323
rect 17969 17289 18003 17323
rect 18003 17289 18012 17323
rect 17960 17280 18012 17289
rect 18880 17280 18932 17332
rect 19156 17280 19208 17332
rect 20996 17280 21048 17332
rect 24952 17323 25004 17332
rect 24952 17289 24961 17323
rect 24961 17289 24995 17323
rect 24995 17289 25004 17323
rect 24952 17280 25004 17289
rect 25228 17323 25280 17332
rect 25228 17289 25237 17323
rect 25237 17289 25271 17323
rect 25271 17289 25280 17323
rect 25228 17280 25280 17289
rect 2412 17144 2464 17196
rect 8576 17187 8628 17196
rect 8576 17153 8585 17187
rect 8585 17153 8619 17187
rect 8619 17153 8628 17187
rect 8576 17144 8628 17153
rect 15292 17187 15344 17196
rect 15292 17153 15301 17187
rect 15301 17153 15335 17187
rect 15335 17153 15344 17187
rect 15292 17144 15344 17153
rect 15568 17144 15620 17196
rect 940 17076 992 17128
rect 17776 17187 17828 17196
rect 17776 17153 17785 17187
rect 17785 17153 17819 17187
rect 17819 17153 17828 17187
rect 17776 17144 17828 17153
rect 18788 17144 18840 17196
rect 19340 17187 19392 17196
rect 19340 17153 19349 17187
rect 19349 17153 19383 17187
rect 19383 17153 19392 17187
rect 19340 17144 19392 17153
rect 22652 17212 22704 17264
rect 24676 17212 24728 17264
rect 25412 17255 25464 17264
rect 25412 17221 25421 17255
rect 25421 17221 25455 17255
rect 25455 17221 25464 17255
rect 25412 17212 25464 17221
rect 26056 17212 26108 17264
rect 28172 17255 28224 17264
rect 28172 17221 28181 17255
rect 28181 17221 28215 17255
rect 28215 17221 28224 17255
rect 28172 17212 28224 17221
rect 28448 17212 28500 17264
rect 33692 17212 33744 17264
rect 33968 17212 34020 17264
rect 38292 17323 38344 17332
rect 38292 17289 38301 17323
rect 38301 17289 38335 17323
rect 38335 17289 38344 17323
rect 38292 17280 38344 17289
rect 39212 17212 39264 17264
rect 20536 17144 20588 17196
rect 21916 17144 21968 17196
rect 24124 17144 24176 17196
rect 24860 17144 24912 17196
rect 20352 17076 20404 17128
rect 19248 17008 19300 17060
rect 21456 17076 21508 17128
rect 24768 17076 24820 17128
rect 27620 17144 27672 17196
rect 27988 17144 28040 17196
rect 28816 17144 28868 17196
rect 31392 17144 31444 17196
rect 32772 17187 32824 17196
rect 32772 17153 32781 17187
rect 32781 17153 32815 17187
rect 32815 17153 32824 17187
rect 32772 17144 32824 17153
rect 32864 17144 32916 17196
rect 2412 16983 2464 16992
rect 2412 16949 2421 16983
rect 2421 16949 2455 16983
rect 2455 16949 2464 16983
rect 2412 16940 2464 16949
rect 17132 16940 17184 16992
rect 17224 16940 17276 16992
rect 22284 17008 22336 17060
rect 29000 17076 29052 17128
rect 32220 17076 32272 17128
rect 32588 17119 32640 17128
rect 32588 17085 32597 17119
rect 32597 17085 32631 17119
rect 32631 17085 32640 17119
rect 32588 17076 32640 17085
rect 32680 17119 32732 17128
rect 32680 17085 32689 17119
rect 32689 17085 32723 17119
rect 32723 17085 32732 17119
rect 32680 17076 32732 17085
rect 33416 17076 33468 17128
rect 33508 17076 33560 17128
rect 40960 17187 41012 17196
rect 40960 17153 40969 17187
rect 40969 17153 41003 17187
rect 41003 17153 41012 17187
rect 40960 17144 41012 17153
rect 41144 17212 41196 17264
rect 51908 17280 51960 17332
rect 53932 17280 53984 17332
rect 55956 17280 56008 17332
rect 56324 17323 56376 17332
rect 56324 17289 56333 17323
rect 56333 17289 56367 17323
rect 56367 17289 56376 17323
rect 56324 17280 56376 17289
rect 47952 17144 48004 17196
rect 51448 17187 51500 17196
rect 51448 17153 51457 17187
rect 51457 17153 51491 17187
rect 51491 17153 51500 17187
rect 51448 17144 51500 17153
rect 27712 17008 27764 17060
rect 27896 17008 27948 17060
rect 19524 16983 19576 16992
rect 19524 16949 19533 16983
rect 19533 16949 19567 16983
rect 19567 16949 19576 16983
rect 19524 16940 19576 16949
rect 20352 16940 20404 16992
rect 23664 16940 23716 16992
rect 29184 16940 29236 16992
rect 33508 16940 33560 16992
rect 38844 17076 38896 17128
rect 39948 17076 40000 17128
rect 40868 17076 40920 17128
rect 41328 17076 41380 17128
rect 54576 17212 54628 17264
rect 51632 17187 51684 17196
rect 51632 17153 51641 17187
rect 51641 17153 51675 17187
rect 51675 17153 51684 17187
rect 51632 17144 51684 17153
rect 51816 17076 51868 17128
rect 53932 17119 53984 17128
rect 53932 17085 53941 17119
rect 53941 17085 53975 17119
rect 53975 17085 53984 17119
rect 53932 17076 53984 17085
rect 54116 17187 54168 17196
rect 54116 17153 54125 17187
rect 54125 17153 54159 17187
rect 54159 17153 54168 17187
rect 54116 17144 54168 17153
rect 58072 17212 58124 17264
rect 55128 17187 55180 17196
rect 55128 17153 55137 17187
rect 55137 17153 55171 17187
rect 55171 17153 55180 17187
rect 55128 17144 55180 17153
rect 34796 16940 34848 16992
rect 36912 16940 36964 16992
rect 40224 16940 40276 16992
rect 44180 16940 44232 16992
rect 54300 16983 54352 16992
rect 54300 16949 54309 16983
rect 54309 16949 54343 16983
rect 54343 16949 54352 16983
rect 54300 16940 54352 16949
rect 55312 17187 55364 17196
rect 55312 17153 55321 17187
rect 55321 17153 55355 17187
rect 55355 17153 55364 17187
rect 55312 17144 55364 17153
rect 56232 17144 56284 17196
rect 55956 17119 56008 17128
rect 55956 17085 55965 17119
rect 55965 17085 55999 17119
rect 55999 17085 56008 17119
rect 55956 17076 56008 17085
rect 58992 17076 59044 17128
rect 57152 16940 57204 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 16212 16779 16264 16788
rect 16212 16745 16221 16779
rect 16221 16745 16255 16779
rect 16255 16745 16264 16779
rect 16212 16736 16264 16745
rect 18788 16736 18840 16788
rect 12808 16668 12860 16720
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 18696 16711 18748 16720
rect 18696 16677 18705 16711
rect 18705 16677 18739 16711
rect 18739 16677 18748 16711
rect 18696 16668 18748 16677
rect 19524 16668 19576 16720
rect 22652 16779 22704 16788
rect 22652 16745 22661 16779
rect 22661 16745 22695 16779
rect 22695 16745 22704 16779
rect 22652 16736 22704 16745
rect 28908 16736 28960 16788
rect 29000 16736 29052 16788
rect 41144 16736 41196 16788
rect 52920 16736 52972 16788
rect 55312 16736 55364 16788
rect 56600 16736 56652 16788
rect 10416 16532 10468 16584
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 12256 16532 12308 16541
rect 13360 16575 13412 16584
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 940 16464 992 16516
rect 11152 16464 11204 16516
rect 16396 16575 16448 16584
rect 16396 16541 16405 16575
rect 16405 16541 16439 16575
rect 16439 16541 16448 16575
rect 16396 16532 16448 16541
rect 11704 16396 11756 16448
rect 13912 16464 13964 16516
rect 16948 16532 17000 16584
rect 17132 16575 17184 16584
rect 17132 16541 17166 16575
rect 17166 16541 17184 16575
rect 17132 16532 17184 16541
rect 19248 16600 19300 16652
rect 31760 16668 31812 16720
rect 32772 16668 32824 16720
rect 40684 16668 40736 16720
rect 41328 16668 41380 16720
rect 20812 16643 20864 16652
rect 20812 16609 20821 16643
rect 20821 16609 20855 16643
rect 20855 16609 20864 16643
rect 20812 16600 20864 16609
rect 18880 16575 18932 16584
rect 18880 16541 18889 16575
rect 18889 16541 18923 16575
rect 18923 16541 18932 16575
rect 18880 16532 18932 16541
rect 17224 16464 17276 16516
rect 19524 16532 19576 16584
rect 20352 16575 20404 16584
rect 20352 16541 20361 16575
rect 20361 16541 20395 16575
rect 20395 16541 20404 16575
rect 20352 16532 20404 16541
rect 21088 16575 21140 16584
rect 21088 16541 21122 16575
rect 21122 16541 21140 16575
rect 21088 16532 21140 16541
rect 22652 16575 22704 16584
rect 22652 16541 22661 16575
rect 22661 16541 22695 16575
rect 22695 16541 22704 16575
rect 22652 16532 22704 16541
rect 22836 16575 22888 16584
rect 22836 16541 22845 16575
rect 22845 16541 22879 16575
rect 22879 16541 22888 16575
rect 22836 16532 22888 16541
rect 24584 16532 24636 16584
rect 27528 16600 27580 16652
rect 28448 16643 28500 16652
rect 28448 16609 28457 16643
rect 28457 16609 28491 16643
rect 28491 16609 28500 16643
rect 28448 16600 28500 16609
rect 28632 16643 28684 16652
rect 28632 16609 28641 16643
rect 28641 16609 28675 16643
rect 28675 16609 28684 16643
rect 28632 16600 28684 16609
rect 29000 16600 29052 16652
rect 30012 16600 30064 16652
rect 26516 16532 26568 16584
rect 26608 16532 26660 16584
rect 18420 16396 18472 16448
rect 18788 16396 18840 16448
rect 26056 16464 26108 16516
rect 27160 16464 27212 16516
rect 21916 16396 21968 16448
rect 24492 16396 24544 16448
rect 26148 16396 26200 16448
rect 27252 16396 27304 16448
rect 27712 16396 27764 16448
rect 28356 16439 28408 16448
rect 28356 16405 28365 16439
rect 28365 16405 28399 16439
rect 28399 16405 28408 16439
rect 28356 16396 28408 16405
rect 32404 16464 32456 16516
rect 32864 16600 32916 16652
rect 36728 16643 36780 16652
rect 36728 16609 36737 16643
rect 36737 16609 36771 16643
rect 36771 16609 36780 16643
rect 36728 16600 36780 16609
rect 36912 16643 36964 16652
rect 36912 16609 36921 16643
rect 36921 16609 36955 16643
rect 36955 16609 36964 16643
rect 36912 16600 36964 16609
rect 37188 16600 37240 16652
rect 40040 16600 40092 16652
rect 51540 16668 51592 16720
rect 33232 16575 33284 16584
rect 33232 16541 33266 16575
rect 33266 16541 33284 16575
rect 33232 16532 33284 16541
rect 36544 16532 36596 16584
rect 38292 16532 38344 16584
rect 40684 16575 40736 16584
rect 40684 16541 40693 16575
rect 40693 16541 40727 16575
rect 40727 16541 40736 16575
rect 40684 16532 40736 16541
rect 35808 16464 35860 16516
rect 36176 16464 36228 16516
rect 32496 16396 32548 16448
rect 33968 16396 34020 16448
rect 36268 16439 36320 16448
rect 36268 16405 36277 16439
rect 36277 16405 36311 16439
rect 36311 16405 36320 16439
rect 36268 16396 36320 16405
rect 38844 16439 38896 16448
rect 38844 16405 38853 16439
rect 38853 16405 38887 16439
rect 38887 16405 38896 16439
rect 38844 16396 38896 16405
rect 40500 16439 40552 16448
rect 40500 16405 40509 16439
rect 40509 16405 40543 16439
rect 40543 16405 40552 16439
rect 40500 16396 40552 16405
rect 40960 16575 41012 16584
rect 40960 16541 40969 16575
rect 40969 16541 41003 16575
rect 41003 16541 41012 16575
rect 40960 16532 41012 16541
rect 41052 16575 41104 16584
rect 41052 16541 41061 16575
rect 41061 16541 41095 16575
rect 41095 16541 41104 16575
rect 41052 16532 41104 16541
rect 42800 16600 42852 16652
rect 44272 16600 44324 16652
rect 46756 16600 46808 16652
rect 51816 16600 51868 16652
rect 41972 16575 42024 16584
rect 41972 16541 41981 16575
rect 41981 16541 42015 16575
rect 42015 16541 42024 16575
rect 41972 16532 42024 16541
rect 42064 16575 42116 16584
rect 42064 16541 42073 16575
rect 42073 16541 42107 16575
rect 42107 16541 42116 16575
rect 42064 16532 42116 16541
rect 51632 16575 51684 16584
rect 51632 16541 51641 16575
rect 51641 16541 51675 16575
rect 51675 16541 51684 16575
rect 51632 16532 51684 16541
rect 54300 16532 54352 16584
rect 58808 16532 58860 16584
rect 43444 16464 43496 16516
rect 46388 16464 46440 16516
rect 47676 16464 47728 16516
rect 56784 16464 56836 16516
rect 58992 16464 59044 16516
rect 41696 16396 41748 16448
rect 42708 16396 42760 16448
rect 45560 16396 45612 16448
rect 46572 16439 46624 16448
rect 46572 16405 46581 16439
rect 46581 16405 46615 16439
rect 46615 16405 46624 16439
rect 46572 16396 46624 16405
rect 51816 16439 51868 16448
rect 51816 16405 51825 16439
rect 51825 16405 51859 16439
rect 51859 16405 51868 16439
rect 51816 16396 51868 16405
rect 52920 16396 52972 16448
rect 55312 16396 55364 16448
rect 56232 16396 56284 16448
rect 58072 16439 58124 16448
rect 58072 16405 58081 16439
rect 58081 16405 58115 16439
rect 58115 16405 58124 16439
rect 58072 16396 58124 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 13544 16235 13596 16244
rect 13544 16201 13553 16235
rect 13553 16201 13587 16235
rect 13587 16201 13596 16235
rect 13544 16192 13596 16201
rect 20352 16192 20404 16244
rect 18972 16124 19024 16176
rect 19248 16167 19300 16176
rect 19248 16133 19257 16167
rect 19257 16133 19291 16167
rect 19291 16133 19300 16167
rect 19248 16124 19300 16133
rect 20536 16124 20588 16176
rect 22928 16192 22980 16244
rect 23296 16192 23348 16244
rect 24124 16235 24176 16244
rect 24124 16201 24133 16235
rect 24133 16201 24167 16235
rect 24167 16201 24176 16235
rect 24124 16192 24176 16201
rect 24676 16192 24728 16244
rect 26608 16192 26660 16244
rect 27160 16235 27212 16244
rect 27160 16201 27169 16235
rect 27169 16201 27203 16235
rect 27203 16201 27212 16235
rect 27160 16192 27212 16201
rect 27528 16235 27580 16244
rect 27528 16201 27537 16235
rect 27537 16201 27571 16235
rect 27571 16201 27580 16235
rect 27528 16192 27580 16201
rect 31116 16192 31168 16244
rect 31300 16192 31352 16244
rect 36728 16192 36780 16244
rect 1860 16056 1912 16108
rect 10324 16056 10376 16108
rect 11704 16099 11756 16108
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 940 15988 992 16040
rect 13360 16056 13412 16108
rect 13820 16099 13872 16108
rect 13820 16065 13829 16099
rect 13829 16065 13863 16099
rect 13863 16065 13872 16099
rect 13820 16056 13872 16065
rect 13912 16099 13964 16108
rect 13912 16065 13921 16099
rect 13921 16065 13955 16099
rect 13955 16065 13964 16099
rect 13912 16056 13964 16065
rect 15752 16099 15804 16108
rect 15752 16065 15761 16099
rect 15761 16065 15795 16099
rect 15795 16065 15804 16099
rect 15752 16056 15804 16065
rect 17040 16099 17092 16108
rect 17040 16065 17049 16099
rect 17049 16065 17083 16099
rect 17083 16065 17092 16099
rect 17040 16056 17092 16065
rect 17776 16056 17828 16108
rect 18696 16056 18748 16108
rect 19156 16099 19208 16108
rect 19156 16065 19165 16099
rect 19165 16065 19199 16099
rect 19199 16065 19208 16099
rect 19156 16056 19208 16065
rect 23572 16124 23624 16176
rect 14096 15988 14148 16040
rect 21916 16056 21968 16108
rect 23204 16056 23256 16108
rect 23848 16056 23900 16108
rect 9680 15852 9732 15904
rect 12624 15895 12676 15904
rect 12624 15861 12633 15895
rect 12633 15861 12667 15895
rect 12667 15861 12676 15895
rect 12624 15852 12676 15861
rect 15200 15852 15252 15904
rect 19892 15852 19944 15904
rect 23848 15920 23900 15972
rect 24308 16056 24360 16108
rect 25136 16056 25188 16108
rect 25596 16124 25648 16176
rect 26056 16056 26108 16108
rect 28356 16056 28408 16108
rect 29552 16167 29604 16176
rect 29552 16133 29561 16167
rect 29561 16133 29595 16167
rect 29595 16133 29604 16167
rect 29552 16124 29604 16133
rect 31208 16167 31260 16176
rect 31208 16133 31217 16167
rect 31217 16133 31251 16167
rect 31251 16133 31260 16167
rect 31208 16124 31260 16133
rect 32312 16124 32364 16176
rect 40040 16192 40092 16244
rect 40132 16192 40184 16244
rect 40960 16192 41012 16244
rect 41052 16192 41104 16244
rect 45468 16235 45520 16244
rect 45468 16201 45477 16235
rect 45477 16201 45511 16235
rect 45511 16201 45520 16235
rect 45468 16192 45520 16201
rect 46388 16235 46440 16244
rect 46388 16201 46397 16235
rect 46397 16201 46431 16235
rect 46431 16201 46440 16235
rect 46388 16192 46440 16201
rect 46572 16192 46624 16244
rect 51080 16192 51132 16244
rect 25688 15988 25740 16040
rect 27252 15988 27304 16040
rect 27896 15988 27948 16040
rect 28172 15988 28224 16040
rect 29736 16031 29788 16040
rect 29736 15997 29745 16031
rect 29745 15997 29779 16031
rect 29779 15997 29788 16031
rect 29736 15988 29788 15997
rect 26608 15920 26660 15972
rect 31300 15920 31352 15972
rect 31760 16056 31812 16108
rect 31852 16056 31904 16108
rect 40500 16124 40552 16176
rect 41788 16124 41840 16176
rect 42708 16124 42760 16176
rect 43076 16124 43128 16176
rect 51172 16124 51224 16176
rect 51632 16235 51684 16244
rect 51632 16201 51641 16235
rect 51641 16201 51675 16235
rect 51675 16201 51684 16235
rect 51632 16192 51684 16201
rect 51540 16124 51592 16176
rect 53840 16192 53892 16244
rect 54116 16192 54168 16244
rect 35808 16056 35860 16108
rect 41696 16056 41748 16108
rect 42064 16056 42116 16108
rect 42432 16056 42484 16108
rect 37556 15988 37608 16040
rect 41604 16031 41656 16040
rect 41604 15997 41613 16031
rect 41613 15997 41647 16031
rect 41647 15997 41656 16031
rect 41604 15988 41656 15997
rect 42984 16099 43036 16108
rect 42984 16065 42993 16099
rect 42993 16065 43027 16099
rect 43027 16065 43036 16099
rect 42984 16056 43036 16065
rect 44180 16099 44232 16108
rect 44180 16065 44189 16099
rect 44189 16065 44223 16099
rect 44223 16065 44232 16099
rect 44180 16056 44232 16065
rect 47860 16056 47912 16108
rect 50712 16056 50764 16108
rect 51356 16099 51408 16108
rect 51356 16065 51365 16099
rect 51365 16065 51399 16099
rect 51399 16065 51408 16099
rect 51356 16056 51408 16065
rect 55312 16124 55364 16176
rect 21916 15852 21968 15904
rect 23112 15852 23164 15904
rect 23664 15852 23716 15904
rect 23940 15852 23992 15904
rect 24676 15852 24728 15904
rect 28724 15852 28776 15904
rect 32220 15852 32272 15904
rect 32956 15920 33008 15972
rect 40868 15920 40920 15972
rect 41512 15920 41564 15972
rect 42892 15988 42944 16040
rect 47768 16031 47820 16040
rect 47768 15997 47777 16031
rect 47777 15997 47811 16031
rect 47811 15997 47820 16031
rect 47768 15988 47820 15997
rect 50988 15988 51040 16040
rect 52920 16099 52972 16108
rect 52920 16065 52929 16099
rect 52929 16065 52963 16099
rect 52963 16065 52972 16099
rect 52920 16056 52972 16065
rect 53104 16099 53156 16108
rect 53104 16065 53113 16099
rect 53113 16065 53147 16099
rect 53147 16065 53156 16099
rect 53104 16056 53156 16065
rect 53196 16056 53248 16108
rect 53840 16099 53892 16108
rect 53840 16065 53849 16099
rect 53849 16065 53883 16099
rect 53883 16065 53892 16099
rect 53840 16056 53892 16065
rect 54944 16056 54996 16108
rect 36452 15852 36504 15904
rect 37096 15852 37148 15904
rect 38200 15852 38252 15904
rect 46848 15852 46900 15904
rect 48136 15852 48188 15904
rect 50712 15895 50764 15904
rect 50712 15861 50721 15895
rect 50721 15861 50755 15895
rect 50755 15861 50764 15895
rect 50712 15852 50764 15861
rect 51540 15852 51592 15904
rect 53840 15852 53892 15904
rect 55128 15852 55180 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 10324 15691 10376 15700
rect 10324 15657 10333 15691
rect 10333 15657 10367 15691
rect 10367 15657 10376 15691
rect 10324 15648 10376 15657
rect 10416 15648 10468 15700
rect 17776 15691 17828 15700
rect 17776 15657 17785 15691
rect 17785 15657 17819 15691
rect 17819 15657 17828 15691
rect 17776 15648 17828 15657
rect 17132 15580 17184 15632
rect 11060 15555 11112 15564
rect 11060 15521 11069 15555
rect 11069 15521 11103 15555
rect 11103 15521 11112 15555
rect 11060 15512 11112 15521
rect 12072 15512 12124 15564
rect 13820 15512 13872 15564
rect 22836 15580 22888 15632
rect 23388 15580 23440 15632
rect 24032 15580 24084 15632
rect 24308 15580 24360 15632
rect 28540 15580 28592 15632
rect 36452 15580 36504 15632
rect 41696 15691 41748 15700
rect 41696 15657 41705 15691
rect 41705 15657 41739 15691
rect 41739 15657 41748 15691
rect 41696 15648 41748 15657
rect 42064 15648 42116 15700
rect 45284 15648 45336 15700
rect 48228 15648 48280 15700
rect 51356 15648 51408 15700
rect 53104 15648 53156 15700
rect 58532 15648 58584 15700
rect 9772 15444 9824 15496
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 13268 15487 13320 15496
rect 13268 15453 13277 15487
rect 13277 15453 13311 15487
rect 13311 15453 13320 15487
rect 13268 15444 13320 15453
rect 12624 15376 12676 15428
rect 13912 15444 13964 15496
rect 14280 15487 14332 15496
rect 14280 15453 14289 15487
rect 14289 15453 14323 15487
rect 14323 15453 14332 15487
rect 14280 15444 14332 15453
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 16488 15376 16540 15428
rect 19156 15512 19208 15564
rect 19892 15555 19944 15564
rect 19892 15521 19901 15555
rect 19901 15521 19935 15555
rect 19935 15521 19944 15555
rect 19892 15512 19944 15521
rect 18880 15444 18932 15496
rect 20260 15444 20312 15496
rect 20444 15487 20496 15496
rect 20444 15453 20453 15487
rect 20453 15453 20487 15487
rect 20487 15453 20496 15487
rect 20444 15444 20496 15453
rect 24124 15512 24176 15564
rect 14464 15351 14516 15360
rect 14464 15317 14473 15351
rect 14473 15317 14507 15351
rect 14507 15317 14516 15351
rect 14464 15308 14516 15317
rect 15476 15351 15528 15360
rect 15476 15317 15485 15351
rect 15485 15317 15519 15351
rect 15519 15317 15528 15351
rect 15476 15308 15528 15317
rect 16764 15308 16816 15360
rect 17132 15376 17184 15428
rect 17960 15308 18012 15360
rect 19248 15376 19300 15428
rect 19432 15351 19484 15360
rect 19432 15317 19441 15351
rect 19441 15317 19475 15351
rect 19475 15317 19484 15351
rect 19432 15308 19484 15317
rect 21732 15376 21784 15428
rect 23020 15419 23072 15428
rect 23020 15385 23029 15419
rect 23029 15385 23063 15419
rect 23063 15385 23072 15419
rect 23020 15376 23072 15385
rect 23848 15487 23900 15496
rect 23848 15453 23857 15487
rect 23857 15453 23891 15487
rect 23891 15453 23900 15487
rect 23848 15444 23900 15453
rect 24584 15487 24636 15496
rect 24584 15453 24593 15487
rect 24593 15453 24627 15487
rect 24627 15453 24636 15487
rect 24584 15444 24636 15453
rect 24676 15444 24728 15496
rect 25688 15444 25740 15496
rect 26700 15487 26752 15496
rect 26700 15453 26709 15487
rect 26709 15453 26743 15487
rect 26743 15453 26752 15487
rect 26700 15444 26752 15453
rect 27528 15487 27580 15496
rect 27528 15453 27537 15487
rect 27537 15453 27571 15487
rect 27571 15453 27580 15487
rect 27528 15444 27580 15453
rect 31208 15512 31260 15564
rect 34060 15512 34112 15564
rect 35348 15512 35400 15564
rect 36268 15512 36320 15564
rect 24216 15376 24268 15428
rect 27896 15376 27948 15428
rect 31760 15444 31812 15496
rect 32680 15444 32732 15496
rect 35624 15444 35676 15496
rect 36544 15487 36596 15496
rect 36544 15453 36553 15487
rect 36553 15453 36587 15487
rect 36587 15453 36596 15487
rect 36544 15444 36596 15453
rect 37556 15512 37608 15564
rect 42064 15512 42116 15564
rect 41052 15487 41104 15496
rect 41052 15453 41061 15487
rect 41061 15453 41095 15487
rect 41095 15453 41104 15487
rect 41052 15444 41104 15453
rect 41236 15487 41288 15496
rect 41236 15453 41243 15487
rect 41243 15453 41288 15487
rect 41236 15444 41288 15453
rect 41328 15487 41380 15496
rect 41328 15453 41337 15487
rect 41337 15453 41371 15487
rect 41371 15453 41380 15487
rect 41328 15444 41380 15453
rect 41420 15487 41472 15496
rect 41420 15453 41429 15487
rect 41429 15453 41463 15487
rect 41463 15453 41472 15487
rect 41420 15444 41472 15453
rect 41604 15444 41656 15496
rect 42984 15444 43036 15496
rect 48228 15444 48280 15496
rect 51448 15444 51500 15496
rect 53196 15444 53248 15496
rect 24952 15308 25004 15360
rect 28356 15308 28408 15360
rect 34704 15308 34756 15360
rect 35624 15308 35676 15360
rect 36728 15308 36780 15360
rect 44180 15376 44232 15428
rect 51816 15419 51868 15428
rect 51816 15385 51850 15419
rect 51850 15385 51868 15419
rect 51816 15376 51868 15385
rect 58164 15419 58216 15428
rect 58164 15385 58173 15419
rect 58173 15385 58207 15419
rect 58207 15385 58216 15419
rect 58164 15376 58216 15385
rect 50712 15308 50764 15360
rect 51172 15308 51224 15360
rect 58624 15308 58676 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 940 14900 992 14952
rect 9312 14968 9364 15020
rect 11060 14968 11112 15020
rect 15476 15104 15528 15156
rect 16488 15104 16540 15156
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 12624 14968 12676 15020
rect 12716 15011 12768 15020
rect 12716 14977 12725 15011
rect 12725 14977 12759 15011
rect 12759 14977 12768 15011
rect 12716 14968 12768 14977
rect 14188 14968 14240 15020
rect 14372 14968 14424 15020
rect 11428 14832 11480 14884
rect 14464 14900 14516 14952
rect 12256 14875 12308 14884
rect 12256 14841 12265 14875
rect 12265 14841 12299 14875
rect 12299 14841 12308 14875
rect 12256 14832 12308 14841
rect 10876 14764 10928 14816
rect 12992 14832 13044 14884
rect 13452 14764 13504 14816
rect 13728 14764 13780 14816
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 18972 15104 19024 15156
rect 19248 15147 19300 15156
rect 19248 15113 19257 15147
rect 19257 15113 19291 15147
rect 19291 15113 19300 15147
rect 19248 15104 19300 15113
rect 20444 15104 20496 15156
rect 18144 15079 18196 15088
rect 18144 15045 18153 15079
rect 18153 15045 18187 15079
rect 18187 15045 18196 15079
rect 18144 15036 18196 15045
rect 18696 15036 18748 15088
rect 18880 15079 18932 15088
rect 18880 15045 18889 15079
rect 18889 15045 18923 15079
rect 18923 15045 18932 15079
rect 18880 15036 18932 15045
rect 22560 15104 22612 15156
rect 22744 15104 22796 15156
rect 23664 15104 23716 15156
rect 17040 14900 17092 14952
rect 19432 14968 19484 15020
rect 20260 14968 20312 15020
rect 22652 14968 22704 15020
rect 22744 15011 22796 15020
rect 22744 14977 22786 15011
rect 22786 14977 22796 15011
rect 22744 14968 22796 14977
rect 23480 14968 23532 15020
rect 25136 15104 25188 15156
rect 26700 15104 26752 15156
rect 27896 15147 27948 15156
rect 27896 15113 27905 15147
rect 27905 15113 27939 15147
rect 27939 15113 27948 15147
rect 27896 15104 27948 15113
rect 24308 15079 24360 15088
rect 24308 15045 24317 15079
rect 24317 15045 24351 15079
rect 24351 15045 24360 15079
rect 24308 15036 24360 15045
rect 24952 15036 25004 15088
rect 26332 15036 26384 15088
rect 27436 15036 27488 15088
rect 29460 15104 29512 15156
rect 29552 15104 29604 15156
rect 30840 15104 30892 15156
rect 32956 15104 33008 15156
rect 34428 15104 34480 15156
rect 28724 15079 28776 15088
rect 28724 15045 28758 15079
rect 28758 15045 28776 15079
rect 28724 15036 28776 15045
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 24216 14968 24268 15020
rect 25136 14968 25188 15020
rect 25504 14968 25556 15020
rect 19984 14900 20036 14952
rect 25780 15011 25832 15020
rect 25780 14977 25789 15011
rect 25789 14977 25823 15011
rect 25823 14977 25832 15011
rect 25780 14968 25832 14977
rect 27712 15011 27764 15020
rect 27712 14977 27721 15011
rect 27721 14977 27755 15011
rect 27755 14977 27764 15011
rect 27712 14968 27764 14977
rect 29092 15036 29144 15088
rect 30196 15036 30248 15088
rect 30932 15079 30984 15088
rect 30932 15045 30941 15079
rect 30941 15045 30975 15079
rect 30975 15045 30984 15079
rect 30932 15036 30984 15045
rect 31484 15036 31536 15088
rect 27436 14900 27488 14952
rect 29000 14968 29052 15020
rect 30564 14968 30616 15020
rect 32128 14968 32180 15020
rect 32312 15011 32364 15020
rect 32312 14977 32321 15011
rect 32321 14977 32355 15011
rect 32355 14977 32364 15011
rect 32312 14968 32364 14977
rect 32864 14968 32916 15020
rect 36544 15036 36596 15088
rect 37924 15104 37976 15156
rect 39304 15104 39356 15156
rect 40868 15036 40920 15088
rect 41512 15104 41564 15156
rect 41972 15104 42024 15156
rect 42248 15104 42300 15156
rect 47860 15104 47912 15156
rect 42708 15036 42760 15088
rect 48412 15036 48464 15088
rect 34704 15011 34756 15020
rect 34704 14977 34738 15011
rect 34738 14977 34756 15011
rect 34704 14968 34756 14977
rect 40040 14968 40092 15020
rect 21824 14832 21876 14884
rect 15016 14807 15068 14816
rect 15016 14773 15025 14807
rect 15025 14773 15059 14807
rect 15059 14773 15068 14807
rect 15016 14764 15068 14773
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 16856 14764 16908 14816
rect 19156 14764 19208 14816
rect 23296 14764 23348 14816
rect 24308 14764 24360 14816
rect 24676 14875 24728 14884
rect 24676 14841 24685 14875
rect 24685 14841 24719 14875
rect 24719 14841 24728 14875
rect 24676 14832 24728 14841
rect 25504 14832 25556 14884
rect 25780 14832 25832 14884
rect 26056 14764 26108 14816
rect 31760 14900 31812 14952
rect 38752 14900 38804 14952
rect 41512 15011 41564 15020
rect 41512 14977 41521 15011
rect 41521 14977 41555 15011
rect 41555 14977 41564 15011
rect 41512 14968 41564 14977
rect 41604 15011 41656 15020
rect 41604 14977 41613 15011
rect 41613 14977 41647 15011
rect 41647 14977 41656 15011
rect 41604 14968 41656 14977
rect 42800 14968 42852 15020
rect 58440 14968 58492 15020
rect 29460 14832 29512 14884
rect 29736 14764 29788 14816
rect 31944 14764 31996 14816
rect 32680 14764 32732 14816
rect 46204 14832 46256 14884
rect 35624 14764 35676 14816
rect 38936 14764 38988 14816
rect 39120 14764 39172 14816
rect 40868 14764 40920 14816
rect 42708 14764 42760 14816
rect 42984 14764 43036 14816
rect 44272 14764 44324 14816
rect 48228 14943 48280 14952
rect 48228 14909 48237 14943
rect 48237 14909 48271 14943
rect 48271 14909 48280 14943
rect 48228 14900 48280 14909
rect 46848 14832 46900 14884
rect 50160 14764 50212 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 9312 14467 9364 14476
rect 9312 14433 9321 14467
rect 9321 14433 9355 14467
rect 9355 14433 9364 14467
rect 9312 14424 9364 14433
rect 11428 14467 11480 14476
rect 11428 14433 11437 14467
rect 11437 14433 11471 14467
rect 11471 14433 11480 14467
rect 11428 14424 11480 14433
rect 1584 14399 1636 14408
rect 1584 14365 1593 14399
rect 1593 14365 1627 14399
rect 1627 14365 1636 14399
rect 1584 14356 1636 14365
rect 8852 14356 8904 14408
rect 9864 14356 9916 14408
rect 14004 14424 14056 14476
rect 14188 14424 14240 14476
rect 940 14288 992 14340
rect 11888 14288 11940 14340
rect 9680 14220 9732 14272
rect 10232 14220 10284 14272
rect 15568 14220 15620 14272
rect 17040 14560 17092 14612
rect 18696 14560 18748 14612
rect 19156 14560 19208 14612
rect 21824 14603 21876 14612
rect 21824 14569 21833 14603
rect 21833 14569 21867 14603
rect 21867 14569 21876 14603
rect 21824 14560 21876 14569
rect 17960 14492 18012 14544
rect 26700 14560 26752 14612
rect 31668 14560 31720 14612
rect 31760 14603 31812 14612
rect 31760 14569 31769 14603
rect 31769 14569 31803 14603
rect 31803 14569 31812 14603
rect 31760 14560 31812 14569
rect 32128 14560 32180 14612
rect 33600 14560 33652 14612
rect 38016 14560 38068 14612
rect 52368 14560 52420 14612
rect 58072 14603 58124 14612
rect 58072 14569 58081 14603
rect 58081 14569 58115 14603
rect 58115 14569 58124 14603
rect 58072 14560 58124 14569
rect 16764 14467 16816 14476
rect 16764 14433 16773 14467
rect 16773 14433 16807 14467
rect 16807 14433 16816 14467
rect 16764 14424 16816 14433
rect 17776 14424 17828 14476
rect 16856 14356 16908 14408
rect 18696 14399 18748 14408
rect 18696 14365 18705 14399
rect 18705 14365 18739 14399
rect 18739 14365 18748 14399
rect 18696 14356 18748 14365
rect 18880 14399 18932 14408
rect 18880 14365 18889 14399
rect 18889 14365 18923 14399
rect 18923 14365 18932 14399
rect 18880 14356 18932 14365
rect 19340 14356 19392 14408
rect 20260 14399 20312 14408
rect 20260 14365 20269 14399
rect 20269 14365 20303 14399
rect 20303 14365 20312 14399
rect 20260 14356 20312 14365
rect 25320 14492 25372 14544
rect 25964 14492 26016 14544
rect 23480 14424 23532 14476
rect 23664 14424 23716 14476
rect 29092 14424 29144 14476
rect 22100 14356 22152 14408
rect 22928 14356 22980 14408
rect 23112 14399 23164 14408
rect 23112 14365 23121 14399
rect 23121 14365 23155 14399
rect 23155 14365 23164 14399
rect 23112 14356 23164 14365
rect 23388 14399 23440 14408
rect 23388 14365 23397 14399
rect 23397 14365 23431 14399
rect 23431 14365 23440 14399
rect 23388 14356 23440 14365
rect 22560 14288 22612 14340
rect 22652 14288 22704 14340
rect 23204 14288 23256 14340
rect 24216 14356 24268 14408
rect 24952 14399 25004 14408
rect 24952 14365 24961 14399
rect 24961 14365 24995 14399
rect 24995 14365 25004 14399
rect 24952 14356 25004 14365
rect 25504 14356 25556 14408
rect 25688 14356 25740 14408
rect 25964 14356 26016 14408
rect 29368 14356 29420 14408
rect 29736 14467 29788 14476
rect 29736 14433 29745 14467
rect 29745 14433 29779 14467
rect 29779 14433 29788 14467
rect 29736 14424 29788 14433
rect 32956 14492 33008 14544
rect 37924 14492 37976 14544
rect 42984 14467 43036 14476
rect 24676 14288 24728 14340
rect 16764 14220 16816 14272
rect 20168 14220 20220 14272
rect 20628 14220 20680 14272
rect 25320 14220 25372 14272
rect 25504 14263 25556 14272
rect 25504 14229 25513 14263
rect 25513 14229 25547 14263
rect 25547 14229 25556 14263
rect 25504 14220 25556 14229
rect 27436 14220 27488 14272
rect 29460 14220 29512 14272
rect 31024 14220 31076 14272
rect 31300 14288 31352 14340
rect 32680 14399 32732 14408
rect 32680 14365 32689 14399
rect 32689 14365 32723 14399
rect 32723 14365 32732 14399
rect 32680 14356 32732 14365
rect 32956 14399 33008 14408
rect 32956 14365 32965 14399
rect 32965 14365 32999 14399
rect 32999 14365 33008 14399
rect 32956 14356 33008 14365
rect 32588 14288 32640 14340
rect 32864 14288 32916 14340
rect 33600 14399 33652 14408
rect 33600 14365 33609 14399
rect 33609 14365 33643 14399
rect 33643 14365 33652 14399
rect 33600 14356 33652 14365
rect 37372 14399 37424 14408
rect 37372 14365 37381 14399
rect 37381 14365 37415 14399
rect 37415 14365 37424 14399
rect 37372 14356 37424 14365
rect 37556 14399 37608 14408
rect 37556 14365 37565 14399
rect 37565 14365 37599 14399
rect 37599 14365 37608 14399
rect 37556 14356 37608 14365
rect 40684 14356 40736 14408
rect 42984 14433 42993 14467
rect 42993 14433 43027 14467
rect 43027 14433 43036 14467
rect 42984 14424 43036 14433
rect 43260 14467 43312 14476
rect 43260 14433 43269 14467
rect 43269 14433 43303 14467
rect 43303 14433 43312 14467
rect 43260 14424 43312 14433
rect 41972 14356 42024 14408
rect 42248 14356 42300 14408
rect 42340 14399 42392 14408
rect 42340 14365 42349 14399
rect 42349 14365 42383 14399
rect 42383 14365 42392 14399
rect 42340 14356 42392 14365
rect 42708 14356 42760 14408
rect 36084 14288 36136 14340
rect 39028 14288 39080 14340
rect 49056 14356 49108 14408
rect 57980 14399 58032 14408
rect 57980 14365 57989 14399
rect 57989 14365 58023 14399
rect 58023 14365 58032 14399
rect 57980 14356 58032 14365
rect 39120 14220 39172 14272
rect 40040 14220 40092 14272
rect 41512 14220 41564 14272
rect 43996 14220 44048 14272
rect 44548 14263 44600 14272
rect 44548 14229 44557 14263
rect 44557 14229 44591 14263
rect 44591 14229 44600 14263
rect 44548 14220 44600 14229
rect 56876 14220 56928 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 8852 14059 8904 14068
rect 8852 14025 8861 14059
rect 8861 14025 8895 14059
rect 8895 14025 8904 14059
rect 8852 14016 8904 14025
rect 12440 14016 12492 14068
rect 12716 14016 12768 14068
rect 940 13812 992 13864
rect 11796 13948 11848 14000
rect 11980 13948 12032 14000
rect 16212 14016 16264 14068
rect 16856 14016 16908 14068
rect 17592 14016 17644 14068
rect 18144 14016 18196 14068
rect 20812 14016 20864 14068
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 2504 13812 2556 13864
rect 9772 13812 9824 13864
rect 3424 13744 3476 13796
rect 10048 13744 10100 13796
rect 11612 13744 11664 13796
rect 11152 13719 11204 13728
rect 11152 13685 11161 13719
rect 11161 13685 11195 13719
rect 11195 13685 11204 13719
rect 11152 13676 11204 13685
rect 12256 13812 12308 13864
rect 14556 13880 14608 13932
rect 16764 13880 16816 13932
rect 17408 13880 17460 13932
rect 20352 13948 20404 14000
rect 22376 14059 22428 14068
rect 22376 14025 22385 14059
rect 22385 14025 22419 14059
rect 22419 14025 22428 14059
rect 22376 14016 22428 14025
rect 22468 14059 22520 14068
rect 22468 14025 22477 14059
rect 22477 14025 22511 14059
rect 22511 14025 22520 14059
rect 22468 14016 22520 14025
rect 22560 14016 22612 14068
rect 25964 14016 26016 14068
rect 26148 14059 26200 14068
rect 26148 14025 26157 14059
rect 26157 14025 26191 14059
rect 26191 14025 26200 14059
rect 26148 14016 26200 14025
rect 29092 14016 29144 14068
rect 29368 14059 29420 14068
rect 29368 14025 29377 14059
rect 29377 14025 29411 14059
rect 29411 14025 29420 14059
rect 29368 14016 29420 14025
rect 29920 14016 29972 14068
rect 30840 14016 30892 14068
rect 32864 14016 32916 14068
rect 36360 14016 36412 14068
rect 37372 14016 37424 14068
rect 37924 14016 37976 14068
rect 14832 13812 14884 13864
rect 16028 13812 16080 13864
rect 12348 13744 12400 13796
rect 12624 13676 12676 13728
rect 16580 13744 16632 13796
rect 19432 13812 19484 13864
rect 20168 13880 20220 13932
rect 31300 13948 31352 14000
rect 19524 13744 19576 13796
rect 19708 13744 19760 13796
rect 20628 13744 20680 13796
rect 20996 13855 21048 13864
rect 20996 13821 21005 13855
rect 21005 13821 21039 13855
rect 21039 13821 21048 13855
rect 20996 13812 21048 13821
rect 23940 13880 23992 13932
rect 24216 13880 24268 13932
rect 24768 13923 24820 13932
rect 24768 13889 24777 13923
rect 24777 13889 24811 13923
rect 24811 13889 24820 13923
rect 24768 13880 24820 13889
rect 24952 13923 25004 13932
rect 24952 13889 24961 13923
rect 24961 13889 24995 13923
rect 24995 13889 25004 13923
rect 24952 13880 25004 13889
rect 25044 13923 25096 13932
rect 25044 13889 25053 13923
rect 25053 13889 25087 13923
rect 25087 13889 25096 13923
rect 25044 13880 25096 13889
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 25504 13880 25556 13932
rect 25964 13880 26016 13932
rect 25872 13812 25924 13864
rect 26148 13812 26200 13864
rect 28172 13812 28224 13864
rect 28816 13880 28868 13932
rect 29552 13880 29604 13932
rect 31024 13880 31076 13932
rect 34704 13948 34756 14000
rect 37556 13948 37608 14000
rect 39028 14059 39080 14068
rect 39028 14025 39037 14059
rect 39037 14025 39071 14059
rect 39071 14025 39080 14059
rect 39028 14016 39080 14025
rect 42984 14016 43036 14068
rect 43996 14016 44048 14068
rect 56692 14016 56744 14068
rect 31576 13923 31628 13932
rect 31576 13889 31585 13923
rect 31585 13889 31619 13923
rect 31619 13889 31628 13923
rect 31576 13880 31628 13889
rect 31760 13923 31812 13932
rect 31760 13889 31769 13923
rect 31769 13889 31803 13923
rect 31803 13889 31812 13923
rect 31760 13880 31812 13889
rect 31944 13880 31996 13932
rect 32496 13880 32548 13932
rect 29828 13855 29880 13864
rect 29828 13821 29837 13855
rect 29837 13821 29871 13855
rect 29871 13821 29880 13855
rect 29828 13812 29880 13821
rect 15476 13676 15528 13728
rect 18420 13676 18472 13728
rect 19616 13676 19668 13728
rect 21272 13676 21324 13728
rect 21456 13676 21508 13728
rect 25136 13744 25188 13796
rect 29460 13744 29512 13796
rect 30380 13812 30432 13864
rect 30564 13855 30616 13864
rect 30564 13821 30573 13855
rect 30573 13821 30607 13855
rect 30607 13821 30616 13855
rect 30564 13812 30616 13821
rect 30840 13812 30892 13864
rect 36728 13880 36780 13932
rect 38016 13923 38068 13932
rect 38016 13889 38022 13923
rect 38022 13889 38056 13923
rect 38056 13889 38068 13923
rect 38016 13880 38068 13889
rect 41328 13948 41380 14000
rect 46204 13948 46256 14000
rect 57796 13948 57848 14000
rect 38660 13880 38712 13932
rect 38936 13923 38988 13932
rect 38936 13889 38945 13923
rect 38945 13889 38979 13923
rect 38979 13889 38988 13923
rect 38936 13880 38988 13889
rect 34796 13812 34848 13864
rect 35348 13812 35400 13864
rect 35716 13812 35768 13864
rect 38752 13812 38804 13864
rect 40500 13880 40552 13932
rect 41696 13923 41748 13932
rect 41696 13889 41705 13923
rect 41705 13889 41739 13923
rect 41739 13889 41748 13923
rect 41696 13880 41748 13889
rect 41788 13923 41840 13932
rect 41788 13889 41797 13923
rect 41797 13889 41831 13923
rect 41831 13889 41840 13923
rect 41788 13880 41840 13889
rect 41420 13812 41472 13864
rect 43076 13923 43128 13932
rect 43076 13889 43085 13923
rect 43085 13889 43119 13923
rect 43119 13889 43128 13923
rect 43076 13880 43128 13889
rect 30932 13744 30984 13796
rect 25780 13719 25832 13728
rect 25780 13685 25789 13719
rect 25789 13685 25823 13719
rect 25823 13685 25832 13719
rect 25780 13676 25832 13685
rect 26056 13676 26108 13728
rect 43352 13855 43404 13864
rect 43352 13821 43361 13855
rect 43361 13821 43395 13855
rect 43395 13821 43404 13855
rect 43352 13812 43404 13821
rect 43536 13812 43588 13864
rect 57520 13812 57572 13864
rect 31852 13676 31904 13728
rect 33508 13676 33560 13728
rect 34520 13719 34572 13728
rect 34520 13685 34529 13719
rect 34529 13685 34563 13719
rect 34563 13685 34572 13719
rect 34520 13676 34572 13685
rect 37280 13676 37332 13728
rect 41328 13676 41380 13728
rect 42524 13676 42576 13728
rect 44456 13676 44508 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 9864 13515 9916 13524
rect 9864 13481 9873 13515
rect 9873 13481 9907 13515
rect 9907 13481 9916 13515
rect 9864 13472 9916 13481
rect 10140 13472 10192 13524
rect 14280 13472 14332 13524
rect 15752 13472 15804 13524
rect 13728 13336 13780 13388
rect 16580 13404 16632 13456
rect 18512 13404 18564 13456
rect 18880 13404 18932 13456
rect 20260 13404 20312 13456
rect 17316 13379 17368 13388
rect 17316 13345 17325 13379
rect 17325 13345 17359 13379
rect 17359 13345 17368 13379
rect 17316 13336 17368 13345
rect 17776 13336 17828 13388
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 9680 13311 9732 13320
rect 9680 13277 9689 13311
rect 9689 13277 9723 13311
rect 9723 13277 9732 13311
rect 9680 13268 9732 13277
rect 940 13200 992 13252
rect 10600 13200 10652 13252
rect 10692 13243 10744 13252
rect 10692 13209 10701 13243
rect 10701 13209 10735 13243
rect 10735 13209 10744 13243
rect 10692 13200 10744 13209
rect 12624 13311 12676 13320
rect 12624 13277 12633 13311
rect 12633 13277 12667 13311
rect 12667 13277 12676 13311
rect 12624 13268 12676 13277
rect 13452 13311 13504 13320
rect 13452 13277 13461 13311
rect 13461 13277 13495 13311
rect 13495 13277 13504 13311
rect 13452 13268 13504 13277
rect 15108 13268 15160 13320
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 15384 13311 15436 13320
rect 15384 13277 15393 13311
rect 15393 13277 15427 13311
rect 15427 13277 15436 13311
rect 15384 13268 15436 13277
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 19340 13336 19392 13388
rect 20904 13404 20956 13456
rect 22376 13515 22428 13524
rect 22376 13481 22385 13515
rect 22385 13481 22419 13515
rect 22419 13481 22428 13515
rect 22376 13472 22428 13481
rect 24584 13472 24636 13524
rect 27528 13472 27580 13524
rect 27712 13472 27764 13524
rect 30840 13472 30892 13524
rect 24032 13404 24084 13456
rect 28816 13404 28868 13456
rect 20812 13336 20864 13388
rect 20996 13379 21048 13388
rect 20996 13345 21005 13379
rect 21005 13345 21039 13379
rect 21039 13345 21048 13379
rect 20996 13336 21048 13345
rect 24676 13336 24728 13388
rect 26332 13336 26384 13388
rect 12348 13200 12400 13252
rect 11980 13132 12032 13184
rect 12164 13175 12216 13184
rect 12164 13141 12173 13175
rect 12173 13141 12207 13175
rect 12207 13141 12216 13175
rect 12164 13132 12216 13141
rect 15200 13132 15252 13184
rect 18420 13311 18472 13320
rect 18420 13277 18429 13311
rect 18429 13277 18463 13311
rect 18463 13277 18472 13311
rect 18420 13268 18472 13277
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 19616 13268 19668 13320
rect 20260 13268 20312 13320
rect 20720 13268 20772 13320
rect 21272 13311 21324 13320
rect 21272 13277 21306 13311
rect 21306 13277 21324 13311
rect 21272 13268 21324 13277
rect 24860 13268 24912 13320
rect 19708 13200 19760 13252
rect 20904 13200 20956 13252
rect 23572 13200 23624 13252
rect 28540 13268 28592 13320
rect 30104 13268 30156 13320
rect 15844 13132 15896 13184
rect 16948 13132 17000 13184
rect 18144 13132 18196 13184
rect 21088 13132 21140 13184
rect 21916 13132 21968 13184
rect 28632 13200 28684 13252
rect 31392 13200 31444 13252
rect 31944 13404 31996 13456
rect 31852 13336 31904 13388
rect 32588 13472 32640 13524
rect 38016 13472 38068 13524
rect 33600 13404 33652 13456
rect 38844 13404 38896 13456
rect 43260 13472 43312 13524
rect 57336 13404 57388 13456
rect 32404 13268 32456 13320
rect 35992 13336 36044 13388
rect 36084 13336 36136 13388
rect 41696 13336 41748 13388
rect 33048 13311 33100 13320
rect 33048 13277 33057 13311
rect 33057 13277 33091 13311
rect 33091 13277 33100 13311
rect 33048 13268 33100 13277
rect 24952 13132 25004 13184
rect 31852 13243 31904 13252
rect 31852 13209 31861 13243
rect 31861 13209 31895 13243
rect 31895 13209 31904 13243
rect 31852 13200 31904 13209
rect 35808 13200 35860 13252
rect 36452 13311 36504 13320
rect 36452 13277 36461 13311
rect 36461 13277 36495 13311
rect 36495 13277 36504 13311
rect 36452 13268 36504 13277
rect 38292 13311 38344 13320
rect 38292 13277 38301 13311
rect 38301 13277 38335 13311
rect 38335 13277 38344 13311
rect 38292 13268 38344 13277
rect 38752 13311 38804 13320
rect 38752 13277 38761 13311
rect 38761 13277 38795 13311
rect 38795 13277 38804 13311
rect 38752 13268 38804 13277
rect 39120 13268 39172 13320
rect 44548 13336 44600 13388
rect 58164 13379 58216 13388
rect 58164 13345 58173 13379
rect 58173 13345 58207 13379
rect 58207 13345 58216 13379
rect 58164 13336 58216 13345
rect 41972 13200 42024 13252
rect 31944 13132 31996 13184
rect 32588 13132 32640 13184
rect 36636 13175 36688 13184
rect 36636 13141 36645 13175
rect 36645 13141 36679 13175
rect 36679 13141 36688 13175
rect 36636 13132 36688 13141
rect 42524 13311 42576 13320
rect 42524 13277 42533 13311
rect 42533 13277 42567 13311
rect 42567 13277 42576 13311
rect 42524 13268 42576 13277
rect 42708 13268 42760 13320
rect 46572 13268 46624 13320
rect 42524 13132 42576 13184
rect 58992 13200 59044 13252
rect 57152 13175 57204 13184
rect 57152 13141 57161 13175
rect 57161 13141 57195 13175
rect 57195 13141 57204 13175
rect 57152 13132 57204 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 9772 12928 9824 12980
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 14004 12971 14056 12980
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 15200 12971 15252 12980
rect 15200 12937 15209 12971
rect 15209 12937 15243 12971
rect 15243 12937 15252 12971
rect 15200 12928 15252 12937
rect 15476 12928 15528 12980
rect 14556 12903 14608 12912
rect 14556 12869 14565 12903
rect 14565 12869 14599 12903
rect 14599 12869 14608 12903
rect 14556 12860 14608 12869
rect 15384 12860 15436 12912
rect 10508 12835 10560 12844
rect 10508 12801 10517 12835
rect 10517 12801 10551 12835
rect 10551 12801 10560 12835
rect 10508 12792 10560 12801
rect 11152 12792 11204 12844
rect 12440 12835 12492 12844
rect 12440 12801 12449 12835
rect 12449 12801 12483 12835
rect 12483 12801 12492 12835
rect 12440 12792 12492 12801
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 15108 12792 15160 12844
rect 17316 12835 17368 12844
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 18052 12792 18104 12844
rect 18144 12835 18196 12844
rect 18144 12801 18153 12835
rect 18153 12801 18187 12835
rect 18187 12801 18196 12835
rect 18144 12792 18196 12801
rect 19340 12928 19392 12980
rect 20720 12971 20772 12980
rect 20720 12937 20729 12971
rect 20729 12937 20763 12971
rect 20763 12937 20772 12971
rect 20720 12928 20772 12937
rect 23388 12928 23440 12980
rect 20996 12860 21048 12912
rect 24584 12860 24636 12912
rect 21640 12792 21692 12844
rect 15384 12656 15436 12708
rect 18236 12656 18288 12708
rect 19156 12656 19208 12708
rect 21180 12767 21232 12776
rect 21180 12733 21189 12767
rect 21189 12733 21223 12767
rect 21223 12733 21232 12767
rect 21180 12724 21232 12733
rect 21456 12724 21508 12776
rect 20812 12656 20864 12708
rect 22192 12792 22244 12844
rect 23020 12792 23072 12844
rect 25780 12860 25832 12912
rect 27804 12928 27856 12980
rect 28632 12903 28684 12912
rect 28632 12869 28641 12903
rect 28641 12869 28675 12903
rect 28675 12869 28684 12903
rect 28632 12860 28684 12869
rect 29736 12928 29788 12980
rect 31484 12928 31536 12980
rect 34796 12928 34848 12980
rect 35256 12928 35308 12980
rect 39672 12928 39724 12980
rect 42800 12928 42852 12980
rect 43352 12928 43404 12980
rect 24768 12724 24820 12776
rect 26148 12792 26200 12844
rect 26884 12792 26936 12844
rect 27804 12792 27856 12844
rect 29736 12724 29788 12776
rect 32312 12860 32364 12912
rect 34520 12860 34572 12912
rect 36084 12903 36136 12912
rect 36084 12869 36093 12903
rect 36093 12869 36127 12903
rect 36127 12869 36136 12903
rect 36084 12860 36136 12869
rect 38016 12860 38068 12912
rect 30748 12792 30800 12844
rect 31116 12724 31168 12776
rect 32588 12835 32640 12844
rect 32588 12801 32597 12835
rect 32597 12801 32631 12835
rect 32631 12801 32640 12835
rect 32588 12792 32640 12801
rect 32772 12792 32824 12844
rect 33784 12835 33836 12844
rect 33784 12801 33793 12835
rect 33793 12801 33827 12835
rect 33827 12801 33836 12835
rect 33784 12792 33836 12801
rect 34796 12792 34848 12844
rect 37280 12792 37332 12844
rect 38660 12792 38712 12844
rect 39672 12792 39724 12844
rect 42708 12792 42760 12844
rect 42984 12835 43036 12844
rect 42984 12801 42993 12835
rect 42993 12801 43027 12835
rect 43027 12801 43036 12835
rect 42984 12792 43036 12801
rect 56140 12792 56192 12844
rect 32404 12724 32456 12776
rect 33048 12724 33100 12776
rect 33232 12767 33284 12776
rect 33232 12733 33241 12767
rect 33241 12733 33275 12767
rect 33275 12733 33284 12767
rect 33232 12724 33284 12733
rect 35992 12724 36044 12776
rect 42156 12724 42208 12776
rect 11980 12588 12032 12640
rect 17224 12588 17276 12640
rect 18420 12588 18472 12640
rect 18512 12588 18564 12640
rect 27988 12656 28040 12708
rect 32496 12656 32548 12708
rect 26424 12588 26476 12640
rect 31024 12588 31076 12640
rect 36452 12699 36504 12708
rect 36452 12665 36461 12699
rect 36461 12665 36495 12699
rect 36495 12665 36504 12699
rect 36452 12656 36504 12665
rect 40868 12656 40920 12708
rect 41144 12656 41196 12708
rect 41420 12656 41472 12708
rect 41972 12656 42024 12708
rect 35900 12588 35952 12640
rect 36176 12588 36228 12640
rect 42800 12588 42852 12640
rect 43076 12588 43128 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 10508 12384 10560 12436
rect 11612 12427 11664 12436
rect 11612 12393 11621 12427
rect 11621 12393 11655 12427
rect 11655 12393 11664 12427
rect 11612 12384 11664 12393
rect 2320 12359 2372 12368
rect 2320 12325 2329 12359
rect 2329 12325 2363 12359
rect 2363 12325 2372 12359
rect 2320 12316 2372 12325
rect 6184 12316 6236 12368
rect 14188 12384 14240 12436
rect 14832 12384 14884 12436
rect 16120 12384 16172 12436
rect 18052 12384 18104 12436
rect 19248 12384 19300 12436
rect 21824 12384 21876 12436
rect 22192 12427 22244 12436
rect 22192 12393 22201 12427
rect 22201 12393 22235 12427
rect 22235 12393 22244 12427
rect 22192 12384 22244 12393
rect 9956 12248 10008 12300
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 10600 12180 10652 12232
rect 10692 12223 10744 12232
rect 10692 12189 10701 12223
rect 10701 12189 10735 12223
rect 10735 12189 10744 12223
rect 10692 12180 10744 12189
rect 11980 12180 12032 12232
rect 20260 12316 20312 12368
rect 24860 12316 24912 12368
rect 15016 12248 15068 12300
rect 17960 12248 18012 12300
rect 13176 12112 13228 12164
rect 13360 12112 13412 12164
rect 15752 12180 15804 12232
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 18512 12248 18564 12300
rect 20076 12248 20128 12300
rect 20536 12248 20588 12300
rect 27068 12384 27120 12436
rect 27620 12427 27672 12436
rect 27620 12393 27629 12427
rect 27629 12393 27663 12427
rect 27663 12393 27672 12427
rect 27620 12384 27672 12393
rect 30012 12427 30064 12436
rect 30012 12393 30021 12427
rect 30021 12393 30055 12427
rect 30055 12393 30064 12427
rect 30012 12384 30064 12393
rect 26516 12316 26568 12368
rect 29920 12316 29972 12368
rect 26240 12248 26292 12300
rect 29092 12248 29144 12300
rect 31024 12359 31076 12368
rect 31024 12325 31033 12359
rect 31033 12325 31067 12359
rect 31067 12325 31076 12359
rect 31024 12316 31076 12325
rect 31116 12316 31168 12368
rect 31576 12316 31628 12368
rect 17684 12180 17736 12189
rect 18420 12223 18472 12232
rect 18420 12189 18429 12223
rect 18429 12189 18463 12223
rect 18463 12189 18472 12223
rect 18420 12180 18472 12189
rect 20260 12180 20312 12232
rect 20628 12180 20680 12232
rect 20904 12180 20956 12232
rect 21088 12223 21140 12232
rect 21088 12189 21122 12223
rect 21122 12189 21140 12223
rect 21088 12180 21140 12189
rect 24676 12180 24728 12232
rect 14464 12044 14516 12096
rect 15200 12112 15252 12164
rect 24768 12112 24820 12164
rect 25320 12112 25372 12164
rect 25964 12180 26016 12232
rect 17960 12044 18012 12096
rect 25136 12044 25188 12096
rect 25228 12044 25280 12096
rect 26056 12087 26108 12096
rect 26056 12053 26065 12087
rect 26065 12053 26099 12087
rect 26099 12053 26108 12087
rect 26056 12044 26108 12053
rect 26516 12087 26568 12096
rect 26516 12053 26525 12087
rect 26525 12053 26559 12087
rect 26559 12053 26568 12087
rect 26516 12044 26568 12053
rect 26700 12112 26752 12164
rect 27804 12223 27856 12232
rect 27804 12189 27813 12223
rect 27813 12189 27847 12223
rect 27847 12189 27856 12223
rect 27804 12180 27856 12189
rect 28264 12180 28316 12232
rect 30104 12180 30156 12232
rect 28448 12112 28500 12164
rect 31116 12180 31168 12232
rect 31208 12223 31260 12232
rect 31208 12189 31217 12223
rect 31217 12189 31251 12223
rect 31251 12189 31260 12223
rect 31208 12180 31260 12189
rect 31392 12180 31444 12232
rect 35808 12427 35860 12436
rect 35808 12393 35817 12427
rect 35817 12393 35851 12427
rect 35851 12393 35860 12427
rect 35808 12384 35860 12393
rect 32772 12316 32824 12368
rect 33784 12248 33836 12300
rect 36636 12248 36688 12300
rect 35348 12180 35400 12232
rect 35532 12223 35584 12232
rect 35532 12189 35541 12223
rect 35541 12189 35575 12223
rect 35575 12189 35584 12223
rect 35532 12180 35584 12189
rect 31576 12112 31628 12164
rect 34336 12112 34388 12164
rect 26884 12044 26936 12096
rect 30288 12044 30340 12096
rect 31300 12044 31352 12096
rect 32864 12044 32916 12096
rect 38016 12384 38068 12436
rect 38384 12384 38436 12436
rect 40040 12223 40092 12232
rect 40040 12189 40049 12223
rect 40049 12189 40083 12223
rect 40083 12189 40092 12223
rect 40040 12180 40092 12189
rect 41604 12316 41656 12368
rect 41696 12316 41748 12368
rect 46296 12384 46348 12436
rect 53196 12384 53248 12436
rect 54392 12384 54444 12436
rect 53472 12316 53524 12368
rect 40408 12223 40460 12232
rect 40408 12189 40417 12223
rect 40417 12189 40451 12223
rect 40451 12189 40460 12223
rect 40408 12180 40460 12189
rect 41144 12223 41196 12232
rect 41144 12189 41153 12223
rect 41153 12189 41187 12223
rect 41187 12189 41196 12223
rect 41144 12180 41196 12189
rect 41328 12180 41380 12232
rect 41420 12223 41472 12232
rect 41420 12189 41429 12223
rect 41429 12189 41463 12223
rect 41463 12189 41472 12223
rect 41420 12180 41472 12189
rect 41512 12223 41564 12232
rect 41512 12189 41521 12223
rect 41521 12189 41555 12223
rect 41555 12189 41564 12223
rect 41512 12180 41564 12189
rect 43444 12248 43496 12300
rect 53564 12248 53616 12300
rect 57888 12223 57940 12232
rect 57888 12189 57897 12223
rect 57897 12189 57931 12223
rect 57931 12189 57940 12223
rect 57888 12180 57940 12189
rect 40868 12112 40920 12164
rect 58164 12155 58216 12164
rect 58164 12121 58173 12155
rect 58173 12121 58207 12155
rect 58207 12121 58216 12155
rect 58164 12112 58216 12121
rect 37924 12044 37976 12096
rect 38384 12044 38436 12096
rect 41144 12044 41196 12096
rect 41788 12087 41840 12096
rect 41788 12053 41797 12087
rect 41797 12053 41831 12087
rect 41831 12053 41840 12087
rect 41788 12044 41840 12053
rect 46388 12044 46440 12096
rect 46848 12044 46900 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 2596 11840 2648 11892
rect 11060 11840 11112 11892
rect 13820 11840 13872 11892
rect 14924 11840 14976 11892
rect 940 11772 992 11824
rect 10692 11772 10744 11824
rect 17408 11883 17460 11892
rect 17408 11849 17417 11883
rect 17417 11849 17451 11883
rect 17451 11849 17460 11883
rect 17408 11840 17460 11849
rect 14372 11704 14424 11756
rect 14464 11747 14516 11756
rect 14464 11713 14473 11747
rect 14473 11713 14507 11747
rect 14507 11713 14516 11747
rect 14464 11704 14516 11713
rect 15568 11772 15620 11824
rect 17224 11747 17276 11756
rect 17224 11713 17233 11747
rect 17233 11713 17267 11747
rect 17267 11713 17276 11747
rect 17224 11704 17276 11713
rect 24032 11840 24084 11892
rect 24492 11840 24544 11892
rect 24768 11840 24820 11892
rect 25320 11883 25372 11892
rect 25320 11849 25329 11883
rect 25329 11849 25363 11883
rect 25363 11849 25372 11883
rect 25320 11840 25372 11849
rect 25412 11840 25464 11892
rect 25688 11840 25740 11892
rect 26148 11840 26200 11892
rect 26516 11840 26568 11892
rect 29828 11840 29880 11892
rect 31116 11840 31168 11892
rect 31852 11840 31904 11892
rect 31944 11840 31996 11892
rect 32312 11840 32364 11892
rect 18328 11772 18380 11824
rect 21088 11772 21140 11824
rect 21364 11772 21416 11824
rect 26056 11772 26108 11824
rect 27528 11772 27580 11824
rect 11152 11568 11204 11620
rect 12072 11679 12124 11688
rect 12072 11645 12081 11679
rect 12081 11645 12115 11679
rect 12115 11645 12124 11679
rect 12072 11636 12124 11645
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 12256 11636 12308 11688
rect 20352 11747 20404 11756
rect 20352 11713 20361 11747
rect 20361 11713 20395 11747
rect 20395 11713 20404 11747
rect 20352 11704 20404 11713
rect 19616 11636 19668 11688
rect 20076 11636 20128 11688
rect 20260 11636 20312 11688
rect 20904 11636 20956 11688
rect 25228 11704 25280 11756
rect 25688 11747 25740 11756
rect 25688 11713 25697 11747
rect 25697 11713 25731 11747
rect 25731 11713 25740 11747
rect 25688 11704 25740 11713
rect 26792 11704 26844 11756
rect 24952 11636 25004 11688
rect 26056 11636 26108 11688
rect 29276 11704 29328 11756
rect 29552 11747 29604 11756
rect 29552 11713 29561 11747
rect 29561 11713 29595 11747
rect 29595 11713 29604 11747
rect 29552 11704 29604 11713
rect 29644 11747 29696 11756
rect 29644 11713 29653 11747
rect 29653 11713 29687 11747
rect 29687 11713 29696 11747
rect 29644 11704 29696 11713
rect 29828 11747 29880 11756
rect 29828 11713 29837 11747
rect 29837 11713 29871 11747
rect 29871 11713 29880 11747
rect 29828 11704 29880 11713
rect 31576 11772 31628 11824
rect 31668 11772 31720 11824
rect 35348 11840 35400 11892
rect 35624 11840 35676 11892
rect 42248 11840 42300 11892
rect 56416 11840 56468 11892
rect 33600 11772 33652 11824
rect 41052 11772 41104 11824
rect 41972 11772 42024 11824
rect 30748 11704 30800 11756
rect 32864 11704 32916 11756
rect 32956 11747 33008 11756
rect 32956 11713 32965 11747
rect 32965 11713 32999 11747
rect 32999 11713 33008 11747
rect 32956 11704 33008 11713
rect 33140 11704 33192 11756
rect 33784 11704 33836 11756
rect 35348 11704 35400 11756
rect 38752 11747 38804 11756
rect 38752 11713 38761 11747
rect 38761 11713 38795 11747
rect 38795 11713 38804 11747
rect 38752 11704 38804 11713
rect 41144 11704 41196 11756
rect 42248 11704 42300 11756
rect 42340 11704 42392 11756
rect 46296 11704 46348 11756
rect 59452 11772 59504 11824
rect 48320 11704 48372 11756
rect 58992 11704 59044 11756
rect 11336 11500 11388 11552
rect 12072 11500 12124 11552
rect 15384 11500 15436 11552
rect 16304 11500 16356 11552
rect 16488 11500 16540 11552
rect 19524 11500 19576 11552
rect 19892 11500 19944 11552
rect 20076 11500 20128 11552
rect 24400 11568 24452 11620
rect 32036 11636 32088 11688
rect 41328 11636 41380 11688
rect 43444 11636 43496 11688
rect 43996 11636 44048 11688
rect 46756 11679 46808 11688
rect 46756 11645 46765 11679
rect 46765 11645 46799 11679
rect 46799 11645 46808 11679
rect 46756 11636 46808 11645
rect 46940 11636 46992 11688
rect 28632 11568 28684 11620
rect 25688 11500 25740 11552
rect 29276 11500 29328 11552
rect 29368 11543 29420 11552
rect 29368 11509 29377 11543
rect 29377 11509 29411 11543
rect 29411 11509 29420 11543
rect 29368 11500 29420 11509
rect 30748 11543 30800 11552
rect 30748 11509 30757 11543
rect 30757 11509 30791 11543
rect 30791 11509 30800 11543
rect 30748 11500 30800 11509
rect 44180 11568 44232 11620
rect 45468 11568 45520 11620
rect 35992 11543 36044 11552
rect 35992 11509 36001 11543
rect 36001 11509 36035 11543
rect 36035 11509 36044 11543
rect 35992 11500 36044 11509
rect 36636 11500 36688 11552
rect 46204 11500 46256 11552
rect 46296 11543 46348 11552
rect 46296 11509 46305 11543
rect 46305 11509 46339 11543
rect 46339 11509 46348 11543
rect 46296 11500 46348 11509
rect 52092 11500 52144 11552
rect 57244 11543 57296 11552
rect 57244 11509 57253 11543
rect 57253 11509 57287 11543
rect 57287 11509 57296 11543
rect 57244 11500 57296 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 940 11160 992 11212
rect 11152 11203 11204 11212
rect 11152 11169 11161 11203
rect 11161 11169 11195 11203
rect 11195 11169 11204 11203
rect 11152 11160 11204 11169
rect 15200 11296 15252 11348
rect 15752 11296 15804 11348
rect 19156 11296 19208 11348
rect 11796 11228 11848 11280
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 11888 11160 11940 11212
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 8944 11024 8996 11076
rect 13176 11203 13228 11212
rect 13176 11169 13185 11203
rect 13185 11169 13219 11203
rect 13219 11169 13228 11203
rect 13176 11160 13228 11169
rect 13820 11160 13872 11212
rect 16488 11228 16540 11280
rect 17500 11228 17552 11280
rect 19432 11228 19484 11280
rect 19248 11160 19300 11212
rect 20996 11339 21048 11348
rect 20996 11305 21005 11339
rect 21005 11305 21039 11339
rect 21039 11305 21048 11339
rect 20996 11296 21048 11305
rect 21088 11296 21140 11348
rect 25688 11296 25740 11348
rect 26424 11339 26476 11348
rect 26424 11305 26433 11339
rect 26433 11305 26467 11339
rect 26467 11305 26476 11339
rect 26424 11296 26476 11305
rect 20812 11228 20864 11280
rect 23940 11228 23992 11280
rect 24768 11228 24820 11280
rect 24952 11228 25004 11280
rect 29644 11296 29696 11348
rect 31208 11296 31260 11348
rect 31668 11296 31720 11348
rect 33416 11296 33468 11348
rect 34152 11296 34204 11348
rect 35348 11296 35400 11348
rect 35532 11296 35584 11348
rect 41328 11296 41380 11348
rect 26976 11228 27028 11280
rect 15660 11067 15712 11076
rect 15660 11033 15669 11067
rect 15669 11033 15703 11067
rect 15703 11033 15712 11067
rect 15660 11024 15712 11033
rect 16304 11135 16356 11144
rect 16304 11101 16313 11135
rect 16313 11101 16347 11135
rect 16347 11101 16356 11135
rect 16304 11092 16356 11101
rect 16672 11135 16724 11144
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 16856 11135 16908 11144
rect 16856 11101 16865 11135
rect 16865 11101 16899 11135
rect 16899 11101 16908 11135
rect 16856 11092 16908 11101
rect 17500 11067 17552 11076
rect 17500 11033 17509 11067
rect 17509 11033 17543 11067
rect 17543 11033 17552 11067
rect 17500 11024 17552 11033
rect 18236 11092 18288 11144
rect 19432 11092 19484 11144
rect 25320 11160 25372 11212
rect 26792 11160 26844 11212
rect 29552 11160 29604 11212
rect 32404 11228 32456 11280
rect 32496 11228 32548 11280
rect 33140 11228 33192 11280
rect 19892 11067 19944 11076
rect 12808 10956 12860 11008
rect 13084 10956 13136 11008
rect 17408 10956 17460 11008
rect 17684 10956 17736 11008
rect 19616 10956 19668 11008
rect 19892 11033 19915 11067
rect 19915 11033 19944 11067
rect 19892 11024 19944 11033
rect 21640 11092 21692 11144
rect 22008 11092 22060 11144
rect 25136 11092 25188 11144
rect 27160 11092 27212 11144
rect 27344 11135 27396 11144
rect 27344 11101 27353 11135
rect 27353 11101 27387 11135
rect 27387 11101 27396 11135
rect 27344 11092 27396 11101
rect 27436 11092 27488 11144
rect 24400 11024 24452 11076
rect 24676 11024 24728 11076
rect 27528 11024 27580 11076
rect 28080 11024 28132 11076
rect 28264 11024 28316 11076
rect 30656 11092 30708 11144
rect 31668 11092 31720 11144
rect 31852 11092 31904 11144
rect 32496 11092 32548 11144
rect 35808 11203 35860 11212
rect 35808 11169 35817 11203
rect 35817 11169 35851 11203
rect 35851 11169 35860 11203
rect 35808 11160 35860 11169
rect 35900 11160 35952 11212
rect 36820 11160 36872 11212
rect 33048 11092 33100 11144
rect 33508 11092 33560 11144
rect 39212 11228 39264 11280
rect 38108 11160 38160 11212
rect 38844 11160 38896 11212
rect 42616 11296 42668 11348
rect 46204 11296 46256 11348
rect 57244 11296 57296 11348
rect 46756 11228 46808 11280
rect 53564 11228 53616 11280
rect 38476 11135 38528 11144
rect 38476 11101 38485 11135
rect 38485 11101 38519 11135
rect 38519 11101 38528 11135
rect 38476 11092 38528 11101
rect 41788 11160 41840 11212
rect 42248 11160 42300 11212
rect 30196 11024 30248 11076
rect 20720 10956 20772 11008
rect 25504 10956 25556 11008
rect 26056 10956 26108 11008
rect 30656 10956 30708 11008
rect 31300 11067 31352 11076
rect 31300 11033 31309 11067
rect 31309 11033 31343 11067
rect 31343 11033 31352 11067
rect 31300 11024 31352 11033
rect 32864 11024 32916 11076
rect 33324 11024 33376 11076
rect 33784 11024 33836 11076
rect 34428 11024 34480 11076
rect 35992 11024 36044 11076
rect 37372 11024 37424 11076
rect 38384 11024 38436 11076
rect 41972 11092 42024 11144
rect 42984 11092 43036 11144
rect 43260 11203 43312 11212
rect 43260 11169 43269 11203
rect 43269 11169 43303 11203
rect 43303 11169 43312 11203
rect 43260 11160 43312 11169
rect 45468 11160 45520 11212
rect 39028 11024 39080 11076
rect 39396 11024 39448 11076
rect 40224 11024 40276 11076
rect 40500 11024 40552 11076
rect 40960 11024 41012 11076
rect 41052 11024 41104 11076
rect 42340 11024 42392 11076
rect 42524 11067 42576 11076
rect 42524 11033 42533 11067
rect 42533 11033 42567 11067
rect 42567 11033 42576 11067
rect 42524 11024 42576 11033
rect 44456 11067 44508 11076
rect 44456 11033 44465 11067
rect 44465 11033 44499 11067
rect 44499 11033 44508 11067
rect 44456 11024 44508 11033
rect 46940 11092 46992 11144
rect 47768 11092 47820 11144
rect 54208 11160 54260 11212
rect 57888 11228 57940 11280
rect 53196 11092 53248 11144
rect 53472 11135 53524 11144
rect 53472 11101 53481 11135
rect 53481 11101 53515 11135
rect 53515 11101 53524 11135
rect 53472 11092 53524 11101
rect 56140 11135 56192 11144
rect 56140 11101 56149 11135
rect 56149 11101 56183 11135
rect 56183 11101 56192 11135
rect 56140 11092 56192 11101
rect 56416 11135 56468 11144
rect 56416 11101 56425 11135
rect 56425 11101 56459 11135
rect 56459 11101 56468 11135
rect 56416 11092 56468 11101
rect 56876 11135 56928 11144
rect 56876 11101 56885 11135
rect 56885 11101 56919 11135
rect 56919 11101 56928 11135
rect 56876 11092 56928 11101
rect 35900 10956 35952 11008
rect 39948 10956 40000 11008
rect 46296 11024 46348 11076
rect 46664 11024 46716 11076
rect 56048 11024 56100 11076
rect 56968 11024 57020 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 3516 10752 3568 10804
rect 940 10684 992 10736
rect 9680 10684 9732 10736
rect 12164 10795 12216 10804
rect 12164 10761 12173 10795
rect 12173 10761 12207 10795
rect 12207 10761 12216 10795
rect 12164 10752 12216 10761
rect 17684 10752 17736 10804
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 9588 10659 9640 10668
rect 9588 10625 9598 10659
rect 9598 10625 9632 10659
rect 9632 10625 9640 10659
rect 9588 10616 9640 10625
rect 11336 10616 11388 10668
rect 12808 10616 12860 10668
rect 14004 10616 14056 10668
rect 1676 10548 1728 10600
rect 9588 10412 9640 10464
rect 10968 10412 11020 10464
rect 11152 10412 11204 10464
rect 13176 10480 13228 10532
rect 19340 10752 19392 10804
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 17224 10616 17276 10668
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 17500 10659 17552 10668
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 20536 10684 20588 10736
rect 22284 10752 22336 10804
rect 32956 10752 33008 10804
rect 34336 10752 34388 10804
rect 21456 10684 21508 10736
rect 15476 10548 15528 10600
rect 15936 10591 15988 10600
rect 15936 10557 15945 10591
rect 15945 10557 15979 10591
rect 15979 10557 15988 10591
rect 15936 10548 15988 10557
rect 16948 10591 17000 10600
rect 16948 10557 16957 10591
rect 16957 10557 16991 10591
rect 16991 10557 17000 10591
rect 16948 10548 17000 10557
rect 16120 10480 16172 10532
rect 18420 10548 18472 10600
rect 18604 10548 18656 10600
rect 17224 10480 17276 10532
rect 18512 10480 18564 10532
rect 19432 10616 19484 10668
rect 20904 10616 20956 10668
rect 21088 10548 21140 10600
rect 23756 10616 23808 10668
rect 27804 10684 27856 10736
rect 19708 10480 19760 10532
rect 21824 10480 21876 10532
rect 23848 10548 23900 10600
rect 24124 10548 24176 10600
rect 24952 10591 25004 10600
rect 24952 10557 24961 10591
rect 24961 10557 24995 10591
rect 24995 10557 25004 10591
rect 24952 10548 25004 10557
rect 25780 10548 25832 10600
rect 24308 10523 24360 10532
rect 24308 10489 24317 10523
rect 24317 10489 24351 10523
rect 24351 10489 24360 10523
rect 24308 10480 24360 10489
rect 24492 10480 24544 10532
rect 27068 10616 27120 10668
rect 27620 10616 27672 10668
rect 27896 10659 27948 10668
rect 27896 10625 27905 10659
rect 27905 10625 27939 10659
rect 27939 10625 27948 10659
rect 27896 10616 27948 10625
rect 28264 10616 28316 10668
rect 28540 10659 28592 10668
rect 28540 10625 28556 10659
rect 28556 10625 28590 10659
rect 28590 10625 28592 10659
rect 28540 10616 28592 10625
rect 28816 10659 28868 10668
rect 28816 10625 28825 10659
rect 28825 10625 28859 10659
rect 28859 10625 28868 10659
rect 28816 10616 28868 10625
rect 31760 10684 31812 10736
rect 34612 10752 34664 10804
rect 27804 10548 27856 10600
rect 31024 10616 31076 10668
rect 33140 10659 33192 10668
rect 33140 10625 33149 10659
rect 33149 10625 33183 10659
rect 33183 10625 33192 10659
rect 33140 10616 33192 10625
rect 33324 10659 33376 10668
rect 33324 10625 33331 10659
rect 33331 10625 33376 10659
rect 33324 10616 33376 10625
rect 33416 10659 33468 10668
rect 33416 10625 33425 10659
rect 33425 10625 33459 10659
rect 33459 10625 33468 10659
rect 33416 10616 33468 10625
rect 33508 10659 33560 10668
rect 33508 10625 33517 10659
rect 33517 10625 33551 10659
rect 33551 10625 33560 10659
rect 33508 10616 33560 10625
rect 33876 10616 33928 10668
rect 34244 10659 34296 10668
rect 34244 10625 34253 10659
rect 34253 10625 34287 10659
rect 34287 10625 34296 10659
rect 34244 10616 34296 10625
rect 35348 10752 35400 10804
rect 36176 10752 36228 10804
rect 40684 10752 40736 10804
rect 45192 10752 45244 10804
rect 56968 10752 57020 10804
rect 35164 10616 35216 10668
rect 37556 10684 37608 10736
rect 55772 10684 55824 10736
rect 35440 10659 35492 10668
rect 35440 10625 35449 10659
rect 35449 10625 35483 10659
rect 35483 10625 35492 10659
rect 35440 10616 35492 10625
rect 27160 10480 27212 10532
rect 29276 10548 29328 10600
rect 32588 10548 32640 10600
rect 32680 10548 32732 10600
rect 38384 10659 38436 10668
rect 38384 10625 38393 10659
rect 38393 10625 38427 10659
rect 38427 10625 38436 10659
rect 38384 10616 38436 10625
rect 41328 10616 41380 10668
rect 44180 10659 44232 10668
rect 44180 10625 44189 10659
rect 44189 10625 44223 10659
rect 44223 10625 44232 10659
rect 44180 10616 44232 10625
rect 44824 10616 44876 10668
rect 56784 10616 56836 10668
rect 57888 10616 57940 10668
rect 14832 10455 14884 10464
rect 14832 10421 14841 10455
rect 14841 10421 14875 10455
rect 14875 10421 14884 10455
rect 14832 10412 14884 10421
rect 16856 10412 16908 10464
rect 17316 10412 17368 10464
rect 24124 10412 24176 10464
rect 24584 10412 24636 10464
rect 25136 10412 25188 10464
rect 25412 10412 25464 10464
rect 27988 10412 28040 10464
rect 36544 10480 36596 10532
rect 29552 10412 29604 10464
rect 31760 10412 31812 10464
rect 32312 10412 32364 10464
rect 35164 10412 35216 10464
rect 35532 10455 35584 10464
rect 35532 10421 35541 10455
rect 35541 10421 35575 10455
rect 35575 10421 35584 10455
rect 35532 10412 35584 10421
rect 35716 10455 35768 10464
rect 35716 10421 35725 10455
rect 35725 10421 35759 10455
rect 35759 10421 35768 10455
rect 35716 10412 35768 10421
rect 38016 10412 38068 10464
rect 40040 10548 40092 10600
rect 40684 10591 40736 10600
rect 40684 10557 40693 10591
rect 40693 10557 40727 10591
rect 40727 10557 40736 10591
rect 40684 10548 40736 10557
rect 41604 10412 41656 10464
rect 41788 10412 41840 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 11428 10208 11480 10260
rect 14004 10208 14056 10260
rect 15384 10208 15436 10260
rect 16396 10208 16448 10260
rect 16488 10208 16540 10260
rect 8484 10140 8536 10192
rect 13176 10140 13228 10192
rect 14740 10140 14792 10192
rect 16672 10140 16724 10192
rect 17040 10140 17092 10192
rect 18788 10208 18840 10260
rect 19156 10208 19208 10260
rect 24492 10208 24544 10260
rect 19064 10140 19116 10192
rect 940 10072 992 10124
rect 17224 10072 17276 10124
rect 18512 10072 18564 10124
rect 19432 10072 19484 10124
rect 11336 10004 11388 10056
rect 11704 10004 11756 10056
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 13452 10004 13504 10056
rect 1952 9868 2004 9920
rect 14832 10004 14884 10056
rect 16120 10004 16172 10056
rect 14464 9936 14516 9988
rect 15200 9868 15252 9920
rect 15476 9936 15528 9988
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 16672 10004 16724 10056
rect 17684 10047 17736 10056
rect 17684 10013 17693 10047
rect 17693 10013 17727 10047
rect 17727 10013 17736 10047
rect 17684 10004 17736 10013
rect 20536 10004 20588 10056
rect 17408 9936 17460 9988
rect 18972 9936 19024 9988
rect 21088 10140 21140 10192
rect 21272 10140 21324 10192
rect 21824 10140 21876 10192
rect 24768 10183 24820 10192
rect 24768 10149 24792 10183
rect 24792 10149 24820 10183
rect 24768 10140 24820 10149
rect 24860 10183 24912 10192
rect 24860 10149 24869 10183
rect 24869 10149 24903 10183
rect 24903 10149 24912 10183
rect 24860 10140 24912 10149
rect 27712 10183 27764 10192
rect 27712 10149 27721 10183
rect 27721 10149 27755 10183
rect 27755 10149 27764 10183
rect 27712 10140 27764 10149
rect 23572 10072 23624 10124
rect 25044 10072 25096 10124
rect 25136 10072 25188 10124
rect 21088 10004 21140 10056
rect 20904 9936 20956 9988
rect 16488 9868 16540 9920
rect 16580 9868 16632 9920
rect 16856 9868 16908 9920
rect 19064 9868 19116 9920
rect 21456 9868 21508 9920
rect 21640 9911 21692 9920
rect 21640 9877 21649 9911
rect 21649 9877 21683 9911
rect 21683 9877 21692 9911
rect 21640 9868 21692 9877
rect 22468 9868 22520 9920
rect 24860 10004 24912 10056
rect 25412 10004 25464 10056
rect 26056 10047 26108 10056
rect 26056 10013 26065 10047
rect 26065 10013 26099 10047
rect 26099 10013 26108 10047
rect 26056 10004 26108 10013
rect 26148 10004 26200 10056
rect 26516 10047 26568 10056
rect 26516 10013 26525 10047
rect 26525 10013 26559 10047
rect 26559 10013 26568 10047
rect 26516 10004 26568 10013
rect 27344 10004 27396 10056
rect 27528 9936 27580 9988
rect 31852 10208 31904 10260
rect 33600 10208 33652 10260
rect 34244 10208 34296 10260
rect 36084 10208 36136 10260
rect 34428 10140 34480 10192
rect 28264 10072 28316 10124
rect 29736 10115 29788 10124
rect 29736 10081 29745 10115
rect 29745 10081 29779 10115
rect 29779 10081 29788 10115
rect 29736 10072 29788 10081
rect 29460 10004 29512 10056
rect 30748 10072 30800 10124
rect 38200 10140 38252 10192
rect 29000 9979 29052 9988
rect 29000 9945 29009 9979
rect 29009 9945 29043 9979
rect 29043 9945 29052 9979
rect 29000 9936 29052 9945
rect 29920 9979 29972 9988
rect 29920 9945 29929 9979
rect 29929 9945 29963 9979
rect 29963 9945 29972 9979
rect 29920 9936 29972 9945
rect 25504 9868 25556 9920
rect 26884 9868 26936 9920
rect 27068 9868 27120 9920
rect 28356 9868 28408 9920
rect 28908 9868 28960 9920
rect 32128 10047 32180 10056
rect 32128 10013 32137 10047
rect 32137 10013 32171 10047
rect 32171 10013 32180 10047
rect 32128 10004 32180 10013
rect 32404 10047 32456 10056
rect 32404 10013 32413 10047
rect 32413 10013 32447 10047
rect 32447 10013 32456 10047
rect 32404 10004 32456 10013
rect 33600 10004 33652 10056
rect 33876 10004 33928 10056
rect 35716 10004 35768 10056
rect 35900 10004 35952 10056
rect 30288 9979 30340 9988
rect 30288 9945 30297 9979
rect 30297 9945 30331 9979
rect 30331 9945 30340 9979
rect 30288 9936 30340 9945
rect 31852 9936 31904 9988
rect 32496 9936 32548 9988
rect 30104 9911 30156 9920
rect 30104 9877 30113 9911
rect 30113 9877 30147 9911
rect 30147 9877 30156 9911
rect 30104 9868 30156 9877
rect 30380 9868 30432 9920
rect 30564 9868 30616 9920
rect 32312 9911 32364 9920
rect 32312 9877 32321 9911
rect 32321 9877 32355 9911
rect 32355 9877 32364 9911
rect 32312 9868 32364 9877
rect 35256 9979 35308 9988
rect 35256 9945 35265 9979
rect 35265 9945 35299 9979
rect 35299 9945 35308 9979
rect 35256 9936 35308 9945
rect 35440 9979 35492 9988
rect 35440 9945 35449 9979
rect 35449 9945 35483 9979
rect 35483 9945 35492 9979
rect 35440 9936 35492 9945
rect 37280 9868 37332 9920
rect 38292 10047 38344 10056
rect 38292 10013 38301 10047
rect 38301 10013 38335 10047
rect 38335 10013 38344 10047
rect 38292 10004 38344 10013
rect 39304 10072 39356 10124
rect 41328 10251 41380 10260
rect 41328 10217 41337 10251
rect 41337 10217 41371 10251
rect 41371 10217 41380 10251
rect 41328 10208 41380 10217
rect 39948 10140 40000 10192
rect 41788 10115 41840 10124
rect 41788 10081 41797 10115
rect 41797 10081 41831 10115
rect 41831 10081 41840 10115
rect 41788 10072 41840 10081
rect 46388 10140 46440 10192
rect 42340 10072 42392 10124
rect 42708 10072 42760 10124
rect 38660 9979 38712 9988
rect 38660 9945 38669 9979
rect 38669 9945 38703 9979
rect 38703 9945 38712 9979
rect 38660 9936 38712 9945
rect 39120 9936 39172 9988
rect 41880 9936 41932 9988
rect 44180 10047 44232 10056
rect 44180 10013 44189 10047
rect 44189 10013 44223 10047
rect 44223 10013 44232 10047
rect 44180 10004 44232 10013
rect 44272 10047 44324 10056
rect 44272 10013 44281 10047
rect 44281 10013 44315 10047
rect 44315 10013 44324 10047
rect 44272 10004 44324 10013
rect 46572 10072 46624 10124
rect 58164 10115 58216 10124
rect 58164 10081 58173 10115
rect 58173 10081 58207 10115
rect 58207 10081 58216 10115
rect 58164 10072 58216 10081
rect 46112 10047 46164 10056
rect 46112 10013 46121 10047
rect 46121 10013 46155 10047
rect 46155 10013 46164 10047
rect 46112 10004 46164 10013
rect 52368 10004 52420 10056
rect 44824 9936 44876 9988
rect 55312 9936 55364 9988
rect 38292 9868 38344 9920
rect 38384 9868 38436 9920
rect 45468 9868 45520 9920
rect 46296 9868 46348 9920
rect 46940 9868 46992 9920
rect 56876 9868 56928 9920
rect 58992 9936 59044 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 4068 9528 4120 9580
rect 12808 9528 12860 9580
rect 13452 9571 13504 9580
rect 13452 9537 13461 9571
rect 13461 9537 13495 9571
rect 13495 9537 13504 9571
rect 13452 9528 13504 9537
rect 940 9460 992 9512
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 9680 9460 9732 9512
rect 11060 9460 11112 9512
rect 12348 9460 12400 9512
rect 14464 9528 14516 9580
rect 7196 9392 7248 9444
rect 10784 9392 10836 9444
rect 10968 9324 11020 9376
rect 14372 9324 14424 9376
rect 14924 9392 14976 9444
rect 15476 9571 15528 9580
rect 15476 9537 15485 9571
rect 15485 9537 15519 9571
rect 15519 9537 15528 9571
rect 15476 9528 15528 9537
rect 15936 9596 15988 9648
rect 22008 9664 22060 9716
rect 22836 9664 22888 9716
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 16212 9528 16264 9580
rect 18328 9528 18380 9580
rect 21640 9596 21692 9648
rect 20444 9528 20496 9580
rect 17316 9460 17368 9512
rect 17776 9503 17828 9512
rect 17776 9469 17785 9503
rect 17785 9469 17819 9503
rect 17819 9469 17828 9503
rect 17776 9460 17828 9469
rect 19432 9460 19484 9512
rect 15568 9392 15620 9444
rect 21824 9528 21876 9580
rect 23388 9528 23440 9580
rect 24216 9596 24268 9648
rect 24584 9528 24636 9580
rect 25504 9596 25556 9648
rect 25964 9596 26016 9648
rect 26056 9596 26108 9648
rect 27528 9707 27580 9716
rect 27528 9673 27537 9707
rect 27537 9673 27571 9707
rect 27571 9673 27580 9707
rect 27528 9664 27580 9673
rect 28172 9664 28224 9716
rect 30104 9664 30156 9716
rect 30380 9664 30432 9716
rect 32036 9664 32088 9716
rect 32128 9664 32180 9716
rect 33140 9664 33192 9716
rect 26700 9528 26752 9580
rect 27712 9596 27764 9648
rect 28448 9596 28500 9648
rect 28172 9528 28224 9580
rect 18512 9324 18564 9376
rect 18880 9324 18932 9376
rect 24032 9392 24084 9444
rect 25412 9460 25464 9512
rect 25780 9503 25832 9512
rect 25780 9469 25789 9503
rect 25789 9469 25823 9503
rect 25823 9469 25832 9503
rect 25780 9460 25832 9469
rect 26056 9503 26108 9512
rect 26056 9469 26065 9503
rect 26065 9469 26099 9503
rect 26099 9469 26108 9503
rect 26056 9460 26108 9469
rect 26792 9460 26844 9512
rect 21088 9324 21140 9376
rect 23664 9324 23716 9376
rect 24860 9324 24912 9376
rect 25044 9324 25096 9376
rect 26240 9324 26292 9376
rect 28448 9435 28500 9444
rect 28448 9401 28457 9435
rect 28457 9401 28491 9435
rect 28491 9401 28500 9435
rect 28448 9392 28500 9401
rect 28908 9528 28960 9580
rect 29184 9596 29236 9648
rect 33324 9664 33376 9716
rect 36452 9664 36504 9716
rect 36544 9664 36596 9716
rect 44272 9664 44324 9716
rect 46572 9707 46624 9716
rect 46572 9673 46581 9707
rect 46581 9673 46615 9707
rect 46615 9673 46624 9707
rect 46572 9664 46624 9673
rect 29184 9460 29236 9512
rect 29092 9392 29144 9444
rect 29276 9324 29328 9376
rect 30012 9571 30064 9580
rect 30012 9537 30021 9571
rect 30021 9537 30055 9571
rect 30055 9537 30064 9571
rect 30012 9528 30064 9537
rect 30288 9528 30340 9580
rect 31668 9528 31720 9580
rect 31944 9460 31996 9512
rect 32588 9571 32640 9580
rect 32588 9537 32597 9571
rect 32597 9537 32631 9571
rect 32631 9537 32640 9571
rect 32588 9528 32640 9537
rect 32772 9571 32824 9580
rect 32772 9537 32781 9571
rect 32781 9537 32815 9571
rect 32815 9537 32824 9571
rect 32772 9528 32824 9537
rect 34336 9596 34388 9648
rect 38108 9596 38160 9648
rect 38384 9596 38436 9648
rect 44456 9596 44508 9648
rect 45468 9639 45520 9648
rect 45468 9605 45502 9639
rect 45502 9605 45520 9639
rect 45468 9596 45520 9605
rect 33416 9528 33468 9580
rect 35992 9571 36044 9580
rect 35992 9537 36001 9571
rect 36001 9537 36035 9571
rect 36035 9537 36044 9571
rect 35992 9528 36044 9537
rect 36176 9571 36228 9580
rect 36176 9537 36185 9571
rect 36185 9537 36219 9571
rect 36219 9537 36228 9571
rect 36176 9528 36228 9537
rect 37648 9571 37700 9580
rect 37648 9537 37655 9571
rect 37655 9537 37700 9571
rect 34244 9460 34296 9512
rect 36544 9392 36596 9444
rect 37648 9528 37700 9537
rect 37740 9571 37792 9580
rect 37740 9537 37749 9571
rect 37749 9537 37783 9571
rect 37783 9537 37792 9571
rect 37740 9528 37792 9537
rect 37924 9571 37976 9580
rect 37924 9537 37938 9571
rect 37938 9537 37972 9571
rect 37972 9537 37976 9571
rect 37924 9528 37976 9537
rect 41420 9528 41472 9580
rect 43904 9571 43956 9580
rect 43904 9537 43913 9571
rect 43913 9537 43947 9571
rect 43947 9537 43956 9571
rect 43904 9528 43956 9537
rect 43996 9571 44048 9580
rect 43996 9537 44005 9571
rect 44005 9537 44039 9571
rect 44039 9537 44048 9571
rect 43996 9528 44048 9537
rect 45100 9528 45152 9580
rect 45192 9571 45244 9580
rect 45192 9537 45201 9571
rect 45201 9537 45235 9571
rect 45235 9537 45244 9571
rect 45192 9528 45244 9537
rect 56784 9528 56836 9580
rect 57244 9571 57296 9580
rect 57244 9537 57253 9571
rect 57253 9537 57287 9571
rect 57287 9537 57296 9571
rect 57244 9528 57296 9537
rect 37740 9392 37792 9444
rect 39396 9392 39448 9444
rect 30288 9324 30340 9376
rect 31484 9324 31536 9376
rect 32956 9324 33008 9376
rect 35900 9324 35952 9376
rect 36268 9324 36320 9376
rect 37556 9324 37608 9376
rect 40592 9367 40644 9376
rect 40592 9333 40601 9367
rect 40601 9333 40635 9367
rect 40635 9333 40644 9367
rect 40592 9324 40644 9333
rect 46204 9324 46256 9376
rect 46480 9324 46532 9376
rect 47124 9324 47176 9376
rect 56324 9324 56376 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 25964 9120 26016 9172
rect 27896 9120 27948 9172
rect 12992 9052 13044 9104
rect 13268 9095 13320 9104
rect 13268 9061 13277 9095
rect 13277 9061 13311 9095
rect 13311 9061 13320 9095
rect 13268 9052 13320 9061
rect 12348 8984 12400 9036
rect 15476 9052 15528 9104
rect 16304 9052 16356 9104
rect 17132 9052 17184 9104
rect 18880 9052 18932 9104
rect 20720 9052 20772 9104
rect 21640 9052 21692 9104
rect 13452 8916 13504 8968
rect 940 8848 992 8900
rect 12624 8848 12676 8900
rect 14924 8891 14976 8900
rect 14924 8857 14933 8891
rect 14933 8857 14967 8891
rect 14967 8857 14976 8891
rect 14924 8848 14976 8857
rect 14832 8823 14884 8832
rect 14832 8789 14841 8823
rect 14841 8789 14875 8823
rect 14875 8789 14884 8823
rect 14832 8780 14884 8789
rect 18512 8984 18564 9036
rect 19432 8984 19484 9036
rect 16304 8916 16356 8968
rect 16672 8959 16724 8968
rect 16672 8925 16681 8959
rect 16681 8925 16715 8959
rect 16715 8925 16724 8959
rect 16672 8916 16724 8925
rect 17408 8959 17460 8968
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 16948 8848 17000 8900
rect 17316 8848 17368 8900
rect 18420 8959 18472 8968
rect 18420 8925 18429 8959
rect 18429 8925 18463 8959
rect 18463 8925 18472 8959
rect 18420 8916 18472 8925
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 15108 8780 15160 8789
rect 16672 8780 16724 8832
rect 18328 8780 18380 8832
rect 18420 8780 18472 8832
rect 20260 8848 20312 8900
rect 23940 8916 23992 8968
rect 25136 9052 25188 9104
rect 25504 9052 25556 9104
rect 26332 9052 26384 9104
rect 33876 9120 33928 9172
rect 37740 9163 37792 9172
rect 37740 9129 37749 9163
rect 37749 9129 37783 9163
rect 37783 9129 37792 9163
rect 37740 9120 37792 9129
rect 38016 9120 38068 9172
rect 24952 8984 25004 9036
rect 25044 8916 25096 8968
rect 25136 8959 25188 8968
rect 25136 8925 25145 8959
rect 25145 8925 25179 8959
rect 25179 8925 25188 8959
rect 25136 8916 25188 8925
rect 22652 8848 22704 8900
rect 23480 8891 23532 8900
rect 23480 8857 23489 8891
rect 23489 8857 23523 8891
rect 23523 8857 23532 8891
rect 23480 8848 23532 8857
rect 23664 8891 23716 8900
rect 23664 8857 23673 8891
rect 23673 8857 23707 8891
rect 23707 8857 23716 8891
rect 23664 8848 23716 8857
rect 20904 8823 20956 8832
rect 20904 8789 20913 8823
rect 20913 8789 20947 8823
rect 20947 8789 20956 8823
rect 20904 8780 20956 8789
rect 25412 8848 25464 8900
rect 25780 8916 25832 8968
rect 26056 8984 26108 9036
rect 26976 8984 27028 9036
rect 28816 8984 28868 9036
rect 29000 9027 29052 9036
rect 29000 8993 29009 9027
rect 29009 8993 29043 9027
rect 29043 8993 29052 9027
rect 29000 8984 29052 8993
rect 29092 8984 29144 9036
rect 31852 9052 31904 9104
rect 32956 9052 33008 9104
rect 33140 9052 33192 9104
rect 35808 9052 35860 9104
rect 38292 9052 38344 9104
rect 38660 9095 38712 9104
rect 38660 9061 38669 9095
rect 38669 9061 38703 9095
rect 38703 9061 38712 9095
rect 38660 9052 38712 9061
rect 41420 9163 41472 9172
rect 41420 9129 41429 9163
rect 41429 9129 41463 9163
rect 41463 9129 41472 9163
rect 41420 9120 41472 9129
rect 52368 9120 52420 9172
rect 42708 9052 42760 9104
rect 43904 9052 43956 9104
rect 44916 9052 44968 9104
rect 58348 9120 58400 9172
rect 31392 8984 31444 9036
rect 36268 9027 36320 9036
rect 36268 8993 36277 9027
rect 36277 8993 36311 9027
rect 36311 8993 36320 9027
rect 36268 8984 36320 8993
rect 36728 8984 36780 9036
rect 26608 8916 26660 8968
rect 27896 8916 27948 8968
rect 29184 8916 29236 8968
rect 30840 8916 30892 8968
rect 31484 8916 31536 8968
rect 31852 8916 31904 8968
rect 32128 8959 32180 8968
rect 32128 8925 32137 8959
rect 32137 8925 32171 8959
rect 32171 8925 32180 8959
rect 32128 8916 32180 8925
rect 32588 8916 32640 8968
rect 33416 8916 33468 8968
rect 26240 8848 26292 8900
rect 27712 8848 27764 8900
rect 24032 8780 24084 8832
rect 24952 8780 25004 8832
rect 26700 8780 26752 8832
rect 27528 8780 27580 8832
rect 29736 8891 29788 8900
rect 29736 8857 29745 8891
rect 29745 8857 29779 8891
rect 29779 8857 29788 8891
rect 29736 8848 29788 8857
rect 29828 8848 29880 8900
rect 31668 8891 31720 8900
rect 31668 8857 31677 8891
rect 31677 8857 31711 8891
rect 31711 8857 31720 8891
rect 31668 8848 31720 8857
rect 32404 8891 32456 8900
rect 32404 8857 32413 8891
rect 32413 8857 32447 8891
rect 32447 8857 32456 8891
rect 32404 8848 32456 8857
rect 32680 8848 32732 8900
rect 34152 8959 34204 8968
rect 34152 8925 34161 8959
rect 34161 8925 34195 8959
rect 34195 8925 34204 8959
rect 34152 8916 34204 8925
rect 34244 8959 34296 8968
rect 34244 8925 34253 8959
rect 34253 8925 34287 8959
rect 34287 8925 34296 8959
rect 34244 8916 34296 8925
rect 35808 8959 35860 8968
rect 35808 8925 35817 8959
rect 35817 8925 35851 8959
rect 35851 8925 35860 8959
rect 35808 8916 35860 8925
rect 35900 8916 35952 8968
rect 36360 8959 36412 8968
rect 36360 8925 36369 8959
rect 36369 8925 36403 8959
rect 36403 8925 36412 8959
rect 36360 8916 36412 8925
rect 37188 8959 37240 8968
rect 37188 8925 37197 8959
rect 37197 8925 37231 8959
rect 37231 8925 37240 8959
rect 37188 8916 37240 8925
rect 37464 8959 37516 8968
rect 37464 8925 37473 8959
rect 37473 8925 37507 8959
rect 37507 8925 37516 8959
rect 37464 8916 37516 8925
rect 37832 8984 37884 9036
rect 38108 8984 38160 9036
rect 40040 9027 40092 9036
rect 40040 8993 40049 9027
rect 40049 8993 40083 9027
rect 40083 8993 40092 9027
rect 40040 8984 40092 8993
rect 38568 8916 38620 8968
rect 40132 8916 40184 8968
rect 29552 8780 29604 8832
rect 30656 8780 30708 8832
rect 31392 8823 31444 8832
rect 31392 8789 31401 8823
rect 31401 8789 31435 8823
rect 31435 8789 31444 8823
rect 31392 8780 31444 8789
rect 31484 8823 31536 8832
rect 31484 8789 31493 8823
rect 31493 8789 31527 8823
rect 31527 8789 31536 8823
rect 33968 8891 34020 8900
rect 33968 8857 33977 8891
rect 33977 8857 34011 8891
rect 34011 8857 34020 8891
rect 33968 8848 34020 8857
rect 38200 8848 38252 8900
rect 44456 8959 44508 8968
rect 44456 8925 44465 8959
rect 44465 8925 44499 8959
rect 44499 8925 44508 8959
rect 44456 8916 44508 8925
rect 44548 8916 44600 8968
rect 46112 8959 46164 8968
rect 46112 8925 46121 8959
rect 46121 8925 46155 8959
rect 46155 8925 46164 8959
rect 46112 8916 46164 8925
rect 46296 8959 46348 8968
rect 46296 8925 46305 8959
rect 46305 8925 46339 8959
rect 46339 8925 46348 8959
rect 46296 8916 46348 8925
rect 31484 8780 31536 8789
rect 33232 8823 33284 8832
rect 33232 8789 33241 8823
rect 33241 8789 33275 8823
rect 33275 8789 33284 8823
rect 33232 8780 33284 8789
rect 38936 8780 38988 8832
rect 43720 8891 43772 8900
rect 43720 8857 43729 8891
rect 43729 8857 43763 8891
rect 43763 8857 43772 8891
rect 43720 8848 43772 8857
rect 44180 8848 44232 8900
rect 56140 8959 56192 8968
rect 56140 8925 56149 8959
rect 56149 8925 56183 8959
rect 56183 8925 56192 8959
rect 56140 8916 56192 8925
rect 56324 8959 56376 8968
rect 56324 8925 56333 8959
rect 56333 8925 56367 8959
rect 56367 8925 56376 8959
rect 56324 8916 56376 8925
rect 56876 9027 56928 9036
rect 56876 8993 56885 9027
rect 56885 8993 56919 9027
rect 56919 8993 56928 9027
rect 56876 8984 56928 8993
rect 43904 8780 43956 8832
rect 52276 8848 52328 8900
rect 46664 8780 46716 8832
rect 52368 8780 52420 8832
rect 57244 8780 57296 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 13452 8576 13504 8628
rect 15108 8576 15160 8628
rect 15292 8576 15344 8628
rect 10600 8440 10652 8492
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 16304 8508 16356 8560
rect 16948 8551 17000 8560
rect 16948 8517 16957 8551
rect 16957 8517 16991 8551
rect 16991 8517 17000 8551
rect 16948 8508 17000 8517
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 17500 8619 17552 8628
rect 17500 8585 17509 8619
rect 17509 8585 17543 8619
rect 17543 8585 17552 8619
rect 17500 8576 17552 8585
rect 18052 8576 18104 8628
rect 18420 8508 18472 8560
rect 17868 8440 17920 8492
rect 19156 8576 19208 8628
rect 20260 8619 20312 8628
rect 20260 8585 20269 8619
rect 20269 8585 20303 8619
rect 20303 8585 20312 8619
rect 20260 8576 20312 8585
rect 21180 8576 21232 8628
rect 23388 8576 23440 8628
rect 19248 8508 19300 8560
rect 20904 8508 20956 8560
rect 23296 8551 23348 8560
rect 23296 8517 23305 8551
rect 23305 8517 23339 8551
rect 23339 8517 23348 8551
rect 23296 8508 23348 8517
rect 25320 8619 25372 8628
rect 25320 8585 25329 8619
rect 25329 8585 25363 8619
rect 25363 8585 25372 8619
rect 25320 8576 25372 8585
rect 25964 8619 26016 8628
rect 25964 8585 25973 8619
rect 25973 8585 26007 8619
rect 26007 8585 26016 8619
rect 25964 8576 26016 8585
rect 24032 8508 24084 8560
rect 940 8372 992 8424
rect 15292 8372 15344 8424
rect 16212 8415 16264 8424
rect 16212 8381 16221 8415
rect 16221 8381 16255 8415
rect 16255 8381 16264 8415
rect 16212 8372 16264 8381
rect 16304 8372 16356 8424
rect 17408 8304 17460 8356
rect 21272 8372 21324 8424
rect 23572 8440 23624 8492
rect 23664 8440 23716 8492
rect 24308 8483 24360 8492
rect 24308 8449 24317 8483
rect 24317 8449 24351 8483
rect 24351 8449 24360 8483
rect 24308 8440 24360 8449
rect 24492 8483 24544 8492
rect 24492 8449 24501 8483
rect 24501 8449 24535 8483
rect 24535 8449 24544 8483
rect 24492 8440 24544 8449
rect 24952 8372 25004 8424
rect 26056 8483 26108 8492
rect 26056 8449 26065 8483
rect 26065 8449 26099 8483
rect 26099 8449 26108 8483
rect 26056 8440 26108 8449
rect 25872 8372 25924 8424
rect 26516 8576 26568 8628
rect 27712 8576 27764 8628
rect 28724 8576 28776 8628
rect 31300 8619 31352 8628
rect 31300 8585 31309 8619
rect 31309 8585 31343 8619
rect 31343 8585 31352 8619
rect 31300 8576 31352 8585
rect 31484 8576 31536 8628
rect 31944 8576 31996 8628
rect 32864 8576 32916 8628
rect 29092 8508 29144 8560
rect 30932 8508 30984 8560
rect 31852 8508 31904 8560
rect 33324 8576 33376 8628
rect 35808 8576 35860 8628
rect 36544 8576 36596 8628
rect 27252 8440 27304 8492
rect 27344 8483 27396 8492
rect 27344 8449 27353 8483
rect 27353 8449 27387 8483
rect 27387 8449 27396 8483
rect 27344 8440 27396 8449
rect 27620 8483 27672 8492
rect 27620 8449 27629 8483
rect 27629 8449 27663 8483
rect 27663 8449 27672 8483
rect 27620 8440 27672 8449
rect 27712 8483 27764 8492
rect 27712 8449 27721 8483
rect 27721 8449 27755 8483
rect 27755 8449 27764 8483
rect 27712 8440 27764 8449
rect 27988 8440 28040 8492
rect 28172 8440 28224 8492
rect 29184 8440 29236 8492
rect 29552 8483 29604 8492
rect 29552 8449 29561 8483
rect 29561 8449 29595 8483
rect 29595 8449 29604 8483
rect 29552 8440 29604 8449
rect 31576 8483 31628 8492
rect 31576 8449 31585 8483
rect 31585 8449 31619 8483
rect 31619 8449 31628 8483
rect 31576 8440 31628 8449
rect 35440 8508 35492 8560
rect 32864 8483 32916 8492
rect 32864 8449 32874 8483
rect 32874 8449 32908 8483
rect 32908 8449 32916 8483
rect 32864 8440 32916 8449
rect 33048 8483 33100 8492
rect 33048 8449 33057 8483
rect 33057 8449 33091 8483
rect 33091 8449 33100 8483
rect 33048 8440 33100 8449
rect 28264 8372 28316 8424
rect 28724 8372 28776 8424
rect 29920 8415 29972 8424
rect 29920 8381 29929 8415
rect 29929 8381 29963 8415
rect 29963 8381 29972 8415
rect 29920 8372 29972 8381
rect 33876 8483 33928 8492
rect 33876 8449 33885 8483
rect 33885 8449 33919 8483
rect 33919 8449 33928 8483
rect 33876 8440 33928 8449
rect 33968 8483 34020 8492
rect 33968 8449 33978 8483
rect 33978 8449 34012 8483
rect 34012 8449 34020 8483
rect 33968 8440 34020 8449
rect 34152 8483 34204 8492
rect 34152 8449 34161 8483
rect 34161 8449 34195 8483
rect 34195 8449 34204 8483
rect 34152 8440 34204 8449
rect 34336 8483 34388 8492
rect 36360 8508 36412 8560
rect 37372 8508 37424 8560
rect 38936 8576 38988 8628
rect 40592 8576 40644 8628
rect 34336 8449 34350 8483
rect 34350 8449 34384 8483
rect 34384 8449 34388 8483
rect 34336 8440 34388 8449
rect 36728 8483 36780 8492
rect 36728 8449 36737 8483
rect 36737 8449 36771 8483
rect 36771 8449 36780 8483
rect 36728 8440 36780 8449
rect 37556 8483 37608 8492
rect 37556 8449 37565 8483
rect 37565 8449 37599 8483
rect 37599 8449 37608 8483
rect 37556 8440 37608 8449
rect 23848 8304 23900 8356
rect 29828 8304 29880 8356
rect 30012 8304 30064 8356
rect 30840 8304 30892 8356
rect 31760 8304 31812 8356
rect 34336 8304 34388 8356
rect 35716 8415 35768 8424
rect 35716 8381 35725 8415
rect 35725 8381 35759 8415
rect 35759 8381 35768 8415
rect 35716 8372 35768 8381
rect 35808 8415 35860 8424
rect 35808 8381 35817 8415
rect 35817 8381 35851 8415
rect 35851 8381 35860 8415
rect 35808 8372 35860 8381
rect 36636 8372 36688 8424
rect 38108 8440 38160 8492
rect 38292 8440 38344 8492
rect 38936 8483 38988 8492
rect 38936 8449 38945 8483
rect 38945 8449 38979 8483
rect 38979 8449 38988 8483
rect 38936 8440 38988 8449
rect 39212 8483 39264 8492
rect 39212 8449 39221 8483
rect 39221 8449 39255 8483
rect 39255 8449 39264 8483
rect 39212 8440 39264 8449
rect 39672 8508 39724 8560
rect 37740 8304 37792 8356
rect 39304 8372 39356 8424
rect 39948 8440 40000 8492
rect 44180 8576 44232 8628
rect 46112 8576 46164 8628
rect 46204 8576 46256 8628
rect 58900 8576 58952 8628
rect 42708 8508 42760 8560
rect 43628 8508 43680 8560
rect 38660 8304 38712 8356
rect 43812 8440 43864 8492
rect 44916 8508 44968 8560
rect 44548 8483 44600 8492
rect 44548 8449 44557 8483
rect 44557 8449 44591 8483
rect 44591 8449 44600 8483
rect 44548 8440 44600 8449
rect 44732 8483 44784 8492
rect 44732 8449 44741 8483
rect 44741 8449 44775 8483
rect 44775 8449 44784 8483
rect 44732 8440 44784 8449
rect 46388 8483 46440 8492
rect 46388 8449 46397 8483
rect 46397 8449 46431 8483
rect 46431 8449 46440 8483
rect 46388 8440 46440 8449
rect 45376 8372 45428 8424
rect 46112 8372 46164 8424
rect 58992 8508 59044 8560
rect 53104 8372 53156 8424
rect 57244 8440 57296 8492
rect 58992 8372 59044 8424
rect 12900 8236 12952 8288
rect 22928 8236 22980 8288
rect 27436 8236 27488 8288
rect 27620 8236 27672 8288
rect 27896 8279 27948 8288
rect 27896 8245 27905 8279
rect 27905 8245 27939 8279
rect 27939 8245 27948 8279
rect 27896 8236 27948 8245
rect 28264 8236 28316 8288
rect 32312 8236 32364 8288
rect 36268 8236 36320 8288
rect 36544 8236 36596 8288
rect 36912 8279 36964 8288
rect 36912 8245 36921 8279
rect 36921 8245 36955 8279
rect 36955 8245 36964 8279
rect 36912 8236 36964 8245
rect 37372 8236 37424 8288
rect 40132 8304 40184 8356
rect 43628 8304 43680 8356
rect 56416 8347 56468 8356
rect 56416 8313 56425 8347
rect 56425 8313 56459 8347
rect 56459 8313 56468 8347
rect 56416 8304 56468 8313
rect 40040 8236 40092 8288
rect 46296 8236 46348 8288
rect 54852 8236 54904 8288
rect 58716 8236 58768 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19340 8032 19392 8084
rect 25044 8075 25096 8084
rect 25044 8041 25053 8075
rect 25053 8041 25087 8075
rect 25087 8041 25096 8075
rect 25044 8032 25096 8041
rect 12808 7964 12860 8016
rect 13820 7964 13872 8016
rect 16856 7964 16908 8016
rect 17960 7964 18012 8016
rect 25688 8032 25740 8084
rect 29368 8032 29420 8084
rect 27804 7964 27856 8016
rect 28356 7964 28408 8016
rect 31668 8032 31720 8084
rect 32864 8032 32916 8084
rect 33968 8032 34020 8084
rect 35808 8032 35860 8084
rect 39212 8032 39264 8084
rect 43720 8032 43772 8084
rect 8944 7896 8996 7948
rect 12624 7939 12676 7948
rect 12624 7905 12633 7939
rect 12633 7905 12667 7939
rect 12667 7905 12676 7939
rect 12624 7896 12676 7905
rect 14740 7896 14792 7948
rect 15108 7896 15160 7948
rect 19064 7896 19116 7948
rect 20444 7896 20496 7948
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 7104 7828 7156 7880
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 8760 7828 8812 7880
rect 10140 7828 10192 7880
rect 940 7760 992 7812
rect 2688 7760 2740 7812
rect 9864 7803 9916 7812
rect 9864 7769 9873 7803
rect 9873 7769 9907 7803
rect 9907 7769 9916 7803
rect 9864 7760 9916 7769
rect 12532 7760 12584 7812
rect 10048 7692 10100 7744
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 15844 7828 15896 7880
rect 16120 7828 16172 7880
rect 16948 7828 17000 7880
rect 15568 7760 15620 7812
rect 17500 7871 17552 7880
rect 17500 7837 17509 7871
rect 17509 7837 17543 7871
rect 17543 7837 17552 7871
rect 17500 7828 17552 7837
rect 18052 7871 18104 7880
rect 18052 7837 18061 7871
rect 18061 7837 18095 7871
rect 18095 7837 18104 7871
rect 18052 7828 18104 7837
rect 18512 7828 18564 7880
rect 22928 7828 22980 7880
rect 23480 7896 23532 7948
rect 24308 7896 24360 7948
rect 17868 7760 17920 7812
rect 18420 7760 18472 7812
rect 16488 7692 16540 7744
rect 17040 7692 17092 7744
rect 24124 7760 24176 7812
rect 25044 7896 25096 7948
rect 27436 7896 27488 7948
rect 26424 7828 26476 7880
rect 26700 7871 26752 7880
rect 26700 7837 26709 7871
rect 26709 7837 26743 7871
rect 26743 7837 26752 7871
rect 26700 7828 26752 7837
rect 29184 7896 29236 7948
rect 29276 7896 29328 7948
rect 26608 7760 26660 7812
rect 22652 7735 22704 7744
rect 22652 7701 22661 7735
rect 22661 7701 22695 7735
rect 22695 7701 22704 7735
rect 22652 7692 22704 7701
rect 22928 7692 22980 7744
rect 23112 7735 23164 7744
rect 23112 7701 23121 7735
rect 23121 7701 23155 7735
rect 23155 7701 23164 7735
rect 23112 7692 23164 7701
rect 24768 7735 24820 7744
rect 24768 7701 24777 7735
rect 24777 7701 24811 7735
rect 24811 7701 24820 7735
rect 24768 7692 24820 7701
rect 27160 7692 27212 7744
rect 27896 7760 27948 7812
rect 29276 7760 29328 7812
rect 29092 7735 29144 7744
rect 29092 7701 29101 7735
rect 29101 7701 29135 7735
rect 29135 7701 29144 7735
rect 29092 7692 29144 7701
rect 30012 7871 30064 7880
rect 30012 7837 30021 7871
rect 30021 7837 30055 7871
rect 30055 7837 30064 7871
rect 30012 7828 30064 7837
rect 39948 7964 40000 8016
rect 40040 7964 40092 8016
rect 46388 8032 46440 8084
rect 30288 7896 30340 7948
rect 30472 7896 30524 7948
rect 30472 7803 30524 7812
rect 30472 7769 30481 7803
rect 30481 7769 30515 7803
rect 30515 7769 30524 7803
rect 30472 7760 30524 7769
rect 31668 7871 31720 7880
rect 31668 7837 31677 7871
rect 31677 7837 31711 7871
rect 31711 7837 31720 7871
rect 31668 7828 31720 7837
rect 33232 7828 33284 7880
rect 33416 7828 33468 7880
rect 33140 7803 33192 7812
rect 33140 7769 33149 7803
rect 33149 7769 33183 7803
rect 33183 7769 33192 7803
rect 33140 7760 33192 7769
rect 35348 7828 35400 7880
rect 36084 7871 36136 7880
rect 36084 7837 36093 7871
rect 36093 7837 36127 7871
rect 36127 7837 36136 7871
rect 36084 7828 36136 7837
rect 36912 7828 36964 7880
rect 39028 7896 39080 7948
rect 43904 7896 43956 7948
rect 38108 7871 38160 7880
rect 38108 7837 38118 7871
rect 38118 7837 38152 7871
rect 38152 7837 38160 7871
rect 38108 7828 38160 7837
rect 38200 7828 38252 7880
rect 31668 7692 31720 7744
rect 33048 7735 33100 7744
rect 33048 7701 33057 7735
rect 33057 7701 33091 7735
rect 33091 7701 33100 7735
rect 33048 7692 33100 7701
rect 34520 7692 34572 7744
rect 37004 7760 37056 7812
rect 37556 7760 37608 7812
rect 38292 7803 38344 7812
rect 38292 7769 38301 7803
rect 38301 7769 38335 7803
rect 38335 7769 38344 7803
rect 38292 7760 38344 7769
rect 42708 7828 42760 7880
rect 43628 7828 43680 7880
rect 43996 7871 44048 7880
rect 43996 7837 44005 7871
rect 44005 7837 44039 7871
rect 44039 7837 44048 7871
rect 43996 7828 44048 7837
rect 46480 7896 46532 7948
rect 44732 7828 44784 7880
rect 46112 7828 46164 7880
rect 56784 8032 56836 8084
rect 45100 7760 45152 7812
rect 46572 7760 46624 7812
rect 52276 7760 52328 7812
rect 55772 7760 55824 7812
rect 56140 7803 56192 7812
rect 56140 7769 56149 7803
rect 56149 7769 56183 7803
rect 56183 7769 56192 7803
rect 56140 7760 56192 7769
rect 56876 7939 56928 7948
rect 56876 7905 56885 7939
rect 56885 7905 56919 7939
rect 56919 7905 56928 7939
rect 56876 7896 56928 7905
rect 57888 7760 57940 7812
rect 36360 7692 36412 7744
rect 36544 7692 36596 7744
rect 38384 7692 38436 7744
rect 40776 7692 40828 7744
rect 49424 7692 49476 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 10600 7531 10652 7540
rect 10600 7497 10609 7531
rect 10609 7497 10643 7531
rect 10643 7497 10652 7531
rect 10600 7488 10652 7497
rect 10968 7488 11020 7540
rect 8760 7420 8812 7472
rect 1584 7352 1636 7404
rect 10692 7352 10744 7404
rect 10784 7395 10836 7404
rect 10784 7361 10793 7395
rect 10793 7361 10827 7395
rect 10827 7361 10836 7395
rect 10784 7352 10836 7361
rect 12532 7488 12584 7540
rect 17040 7488 17092 7540
rect 17500 7488 17552 7540
rect 20352 7488 20404 7540
rect 24400 7488 24452 7540
rect 24860 7488 24912 7540
rect 25136 7488 25188 7540
rect 28540 7488 28592 7540
rect 11336 7352 11388 7404
rect 12624 7352 12676 7404
rect 10876 7327 10928 7336
rect 10876 7293 10885 7327
rect 10885 7293 10919 7327
rect 10919 7293 10928 7327
rect 10876 7284 10928 7293
rect 11060 7327 11112 7336
rect 11060 7293 11069 7327
rect 11069 7293 11103 7327
rect 11103 7293 11112 7327
rect 11060 7284 11112 7293
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 9864 7216 9916 7268
rect 10968 7216 11020 7268
rect 7380 7148 7432 7200
rect 15108 7463 15160 7472
rect 15108 7429 15117 7463
rect 15117 7429 15151 7463
rect 15151 7429 15160 7463
rect 15108 7420 15160 7429
rect 15200 7463 15252 7472
rect 15200 7429 15209 7463
rect 15209 7429 15243 7463
rect 15243 7429 15252 7463
rect 15200 7420 15252 7429
rect 15844 7420 15896 7472
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 16672 7420 16724 7472
rect 16856 7420 16908 7472
rect 16948 7463 17000 7472
rect 16948 7429 16957 7463
rect 16957 7429 16991 7463
rect 16991 7429 17000 7463
rect 16948 7420 17000 7429
rect 18512 7463 18564 7472
rect 18512 7429 18521 7463
rect 18521 7429 18555 7463
rect 18555 7429 18564 7463
rect 18512 7420 18564 7429
rect 22928 7420 22980 7472
rect 23572 7420 23624 7472
rect 25504 7420 25556 7472
rect 28632 7463 28684 7472
rect 15292 7284 15344 7336
rect 15844 7284 15896 7336
rect 17316 7352 17368 7404
rect 17500 7395 17552 7404
rect 17500 7361 17509 7395
rect 17509 7361 17543 7395
rect 17543 7361 17552 7395
rect 17500 7352 17552 7361
rect 20628 7352 20680 7404
rect 22008 7395 22060 7404
rect 22008 7361 22023 7395
rect 22023 7361 22057 7395
rect 22057 7361 22060 7395
rect 22008 7352 22060 7361
rect 28632 7429 28641 7463
rect 28641 7429 28675 7463
rect 28675 7429 28684 7463
rect 28632 7420 28684 7429
rect 30012 7488 30064 7540
rect 35532 7531 35584 7540
rect 35532 7497 35541 7531
rect 35541 7497 35575 7531
rect 35575 7497 35584 7531
rect 35532 7488 35584 7497
rect 36728 7488 36780 7540
rect 38108 7488 38160 7540
rect 31300 7420 31352 7472
rect 29092 7352 29144 7404
rect 31024 7352 31076 7404
rect 17592 7284 17644 7336
rect 17868 7284 17920 7336
rect 19432 7284 19484 7336
rect 20076 7327 20128 7336
rect 20076 7293 20085 7327
rect 20085 7293 20119 7327
rect 20119 7293 20128 7327
rect 20076 7284 20128 7293
rect 27712 7327 27764 7336
rect 27712 7293 27721 7327
rect 27721 7293 27755 7327
rect 27755 7293 27764 7327
rect 27712 7284 27764 7293
rect 27988 7284 28040 7336
rect 30656 7284 30708 7336
rect 31484 7327 31536 7336
rect 31484 7293 31493 7327
rect 31493 7293 31527 7327
rect 31527 7293 31536 7327
rect 31484 7284 31536 7293
rect 36084 7420 36136 7472
rect 36544 7463 36596 7472
rect 36544 7429 36553 7463
rect 36553 7429 36587 7463
rect 36587 7429 36596 7463
rect 36544 7420 36596 7429
rect 37004 7420 37056 7472
rect 44548 7463 44600 7472
rect 44548 7429 44557 7463
rect 44557 7429 44591 7463
rect 44591 7429 44600 7463
rect 44548 7420 44600 7429
rect 34428 7395 34480 7404
rect 34428 7361 34462 7395
rect 34462 7361 34480 7395
rect 34428 7352 34480 7361
rect 34796 7352 34848 7404
rect 36728 7352 36780 7404
rect 36820 7327 36872 7336
rect 36820 7293 36829 7327
rect 36829 7293 36863 7327
rect 36863 7293 36872 7327
rect 36820 7284 36872 7293
rect 25044 7216 25096 7268
rect 25136 7216 25188 7268
rect 25412 7216 25464 7268
rect 21456 7191 21508 7200
rect 21456 7157 21465 7191
rect 21465 7157 21499 7191
rect 21499 7157 21508 7191
rect 21456 7148 21508 7157
rect 25504 7148 25556 7200
rect 26516 7148 26568 7200
rect 28264 7216 28316 7268
rect 29736 7216 29788 7268
rect 29920 7216 29972 7268
rect 38384 7352 38436 7404
rect 43996 7352 44048 7404
rect 54852 7420 54904 7472
rect 55772 7463 55824 7472
rect 55772 7429 55781 7463
rect 55781 7429 55815 7463
rect 55815 7429 55824 7463
rect 55772 7420 55824 7429
rect 27988 7191 28040 7200
rect 27988 7157 27997 7191
rect 27997 7157 28031 7191
rect 28031 7157 28040 7191
rect 27988 7148 28040 7157
rect 29644 7148 29696 7200
rect 30196 7148 30248 7200
rect 31116 7148 31168 7200
rect 45376 7395 45428 7404
rect 45376 7361 45385 7395
rect 45385 7361 45419 7395
rect 45419 7361 45428 7395
rect 45376 7352 45428 7361
rect 46296 7395 46348 7404
rect 46296 7361 46305 7395
rect 46305 7361 46339 7395
rect 46339 7361 46348 7395
rect 46296 7352 46348 7361
rect 56140 7420 56192 7472
rect 45100 7284 45152 7336
rect 46480 7327 46532 7336
rect 46480 7293 46489 7327
rect 46489 7293 46523 7327
rect 46523 7293 46532 7327
rect 46480 7284 46532 7293
rect 52276 7216 52328 7268
rect 56692 7352 56744 7404
rect 56784 7352 56836 7404
rect 58256 7395 58308 7404
rect 58256 7361 58265 7395
rect 58265 7361 58299 7395
rect 58299 7361 58308 7395
rect 58256 7352 58308 7361
rect 41512 7148 41564 7200
rect 45468 7148 45520 7200
rect 45836 7191 45888 7200
rect 45836 7157 45845 7191
rect 45845 7157 45879 7191
rect 45879 7157 45888 7191
rect 45836 7148 45888 7157
rect 56968 7148 57020 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 12624 6944 12676 6996
rect 10876 6876 10928 6928
rect 18972 6944 19024 6996
rect 20076 6944 20128 6996
rect 15108 6876 15160 6928
rect 940 6808 992 6860
rect 8760 6808 8812 6860
rect 9128 6740 9180 6792
rect 10692 6808 10744 6860
rect 15752 6808 15804 6860
rect 15936 6808 15988 6860
rect 16396 6808 16448 6860
rect 10876 6740 10928 6792
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 17500 6876 17552 6928
rect 20628 6944 20680 6996
rect 17316 6808 17368 6860
rect 16948 6740 17000 6792
rect 17408 6783 17460 6792
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 17592 6740 17644 6792
rect 19984 6808 20036 6860
rect 20260 6876 20312 6928
rect 23388 6944 23440 6996
rect 24400 6944 24452 6996
rect 24492 6944 24544 6996
rect 27896 6944 27948 6996
rect 28356 6944 28408 6996
rect 31668 6944 31720 6996
rect 34428 6944 34480 6996
rect 39028 6944 39080 6996
rect 46112 6944 46164 6996
rect 46296 6944 46348 6996
rect 21088 6808 21140 6860
rect 21272 6851 21324 6860
rect 21272 6817 21281 6851
rect 21281 6817 21315 6851
rect 21315 6817 21324 6851
rect 21272 6808 21324 6817
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 26056 6740 26108 6792
rect 27160 6808 27212 6860
rect 30012 6876 30064 6928
rect 30748 6876 30800 6928
rect 31484 6876 31536 6928
rect 27620 6808 27672 6860
rect 28080 6808 28132 6860
rect 28632 6808 28684 6860
rect 30932 6808 30984 6860
rect 33784 6808 33836 6860
rect 36820 6808 36872 6860
rect 40040 6808 40092 6860
rect 46848 6808 46900 6860
rect 49608 6808 49660 6860
rect 56876 6851 56928 6860
rect 56876 6817 56885 6851
rect 56885 6817 56919 6851
rect 56919 6817 56928 6851
rect 56876 6808 56928 6817
rect 26976 6783 27028 6792
rect 26976 6749 26985 6783
rect 26985 6749 27019 6783
rect 27019 6749 27028 6783
rect 26976 6740 27028 6749
rect 11336 6672 11388 6724
rect 9496 6604 9548 6656
rect 11704 6604 11756 6656
rect 16120 6672 16172 6724
rect 15752 6604 15804 6656
rect 17868 6672 17920 6724
rect 17960 6672 18012 6724
rect 18236 6672 18288 6724
rect 19432 6672 19484 6724
rect 20444 6672 20496 6724
rect 22376 6672 22428 6724
rect 22652 6672 22704 6724
rect 16580 6604 16632 6656
rect 21456 6604 21508 6656
rect 22192 6604 22244 6656
rect 23848 6647 23900 6656
rect 23848 6613 23857 6647
rect 23857 6613 23891 6647
rect 23891 6613 23900 6647
rect 23848 6604 23900 6613
rect 25044 6604 25096 6656
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 25780 6604 25832 6656
rect 26792 6672 26844 6724
rect 30380 6740 30432 6792
rect 27804 6672 27856 6724
rect 28540 6672 28592 6724
rect 30288 6672 30340 6724
rect 31208 6715 31260 6724
rect 31208 6681 31217 6715
rect 31217 6681 31251 6715
rect 31251 6681 31260 6715
rect 31208 6672 31260 6681
rect 28448 6604 28500 6656
rect 28724 6604 28776 6656
rect 30840 6604 30892 6656
rect 33692 6740 33744 6792
rect 31760 6715 31812 6724
rect 31760 6681 31769 6715
rect 31769 6681 31803 6715
rect 31803 6681 31812 6715
rect 31760 6672 31812 6681
rect 32588 6672 32640 6724
rect 34796 6672 34848 6724
rect 31944 6604 31996 6656
rect 33140 6604 33192 6656
rect 46940 6740 46992 6792
rect 56968 6740 57020 6792
rect 45836 6672 45888 6724
rect 35256 6647 35308 6656
rect 35256 6613 35265 6647
rect 35265 6613 35299 6647
rect 35299 6613 35308 6647
rect 35256 6604 35308 6613
rect 35348 6647 35400 6656
rect 35348 6613 35357 6647
rect 35357 6613 35391 6647
rect 35391 6613 35400 6647
rect 35348 6604 35400 6613
rect 43076 6604 43128 6656
rect 58256 6647 58308 6656
rect 58256 6613 58265 6647
rect 58265 6613 58299 6647
rect 58299 6613 58308 6647
rect 58256 6604 58308 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 13360 6400 13412 6452
rect 9128 6264 9180 6316
rect 940 6196 992 6248
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 9496 6239 9548 6248
rect 9496 6205 9505 6239
rect 9505 6205 9539 6239
rect 9539 6205 9548 6239
rect 9496 6196 9548 6205
rect 10416 6196 10468 6248
rect 12624 6264 12676 6316
rect 19248 6400 19300 6452
rect 19984 6400 20036 6452
rect 20996 6400 21048 6452
rect 23112 6400 23164 6452
rect 15200 6332 15252 6384
rect 18052 6332 18104 6384
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 15844 6307 15896 6316
rect 15844 6273 15853 6307
rect 15853 6273 15887 6307
rect 15887 6273 15896 6307
rect 15844 6264 15896 6273
rect 15936 6264 15988 6316
rect 17500 6264 17552 6316
rect 20260 6332 20312 6384
rect 23204 6332 23256 6384
rect 7932 6060 7984 6112
rect 17960 6128 18012 6180
rect 19984 6264 20036 6316
rect 23388 6307 23440 6316
rect 23388 6273 23397 6307
rect 23397 6273 23431 6307
rect 23431 6273 23440 6307
rect 23388 6264 23440 6273
rect 25136 6400 25188 6452
rect 33048 6400 33100 6452
rect 33140 6400 33192 6452
rect 35256 6400 35308 6452
rect 36452 6400 36504 6452
rect 38844 6400 38896 6452
rect 24584 6332 24636 6384
rect 25044 6375 25096 6384
rect 24400 6264 24452 6316
rect 25044 6341 25078 6375
rect 25078 6341 25096 6375
rect 25044 6332 25096 6341
rect 25228 6332 25280 6384
rect 24032 6196 24084 6248
rect 24308 6196 24360 6248
rect 21088 6128 21140 6180
rect 27344 6264 27396 6316
rect 27620 6264 27672 6316
rect 28540 6332 28592 6384
rect 29368 6332 29420 6384
rect 28632 6307 28684 6316
rect 26608 6196 26660 6248
rect 27804 6239 27856 6248
rect 27804 6205 27813 6239
rect 27813 6205 27847 6239
rect 27847 6205 27856 6239
rect 27804 6196 27856 6205
rect 28632 6273 28641 6307
rect 28641 6273 28675 6307
rect 28675 6273 28684 6307
rect 28632 6264 28684 6273
rect 29276 6264 29328 6316
rect 33784 6332 33836 6384
rect 35532 6375 35584 6384
rect 35532 6341 35541 6375
rect 35541 6341 35575 6375
rect 35575 6341 35584 6375
rect 35532 6332 35584 6341
rect 36912 6332 36964 6384
rect 43260 6332 43312 6384
rect 30932 6307 30984 6316
rect 30932 6273 30941 6307
rect 30941 6273 30975 6307
rect 30975 6273 30984 6307
rect 30932 6264 30984 6273
rect 31116 6307 31168 6316
rect 31116 6273 31125 6307
rect 31125 6273 31159 6307
rect 31159 6273 31168 6307
rect 31116 6264 31168 6273
rect 34520 6307 34572 6316
rect 34520 6273 34529 6307
rect 34529 6273 34563 6307
rect 34563 6273 34572 6307
rect 34520 6264 34572 6273
rect 36084 6264 36136 6316
rect 38476 6264 38528 6316
rect 46848 6332 46900 6384
rect 46388 6307 46440 6316
rect 46388 6273 46397 6307
rect 46397 6273 46431 6307
rect 46431 6273 46440 6307
rect 46388 6264 46440 6273
rect 58072 6307 58124 6316
rect 58072 6273 58081 6307
rect 58081 6273 58115 6307
rect 58115 6273 58124 6307
rect 58072 6264 58124 6273
rect 20996 6060 21048 6112
rect 24676 6060 24728 6112
rect 26056 6060 26108 6112
rect 26148 6103 26200 6112
rect 26148 6069 26157 6103
rect 26157 6069 26191 6103
rect 26191 6069 26200 6103
rect 26148 6060 26200 6069
rect 27988 6060 28040 6112
rect 28356 6128 28408 6180
rect 28908 6128 28960 6180
rect 29920 6128 29972 6180
rect 36728 6196 36780 6248
rect 43444 6196 43496 6248
rect 46572 6239 46624 6248
rect 46572 6205 46581 6239
rect 46581 6205 46615 6239
rect 46615 6205 46624 6239
rect 46572 6196 46624 6205
rect 30380 6128 30432 6180
rect 38200 6128 38252 6180
rect 30748 6060 30800 6112
rect 31392 6060 31444 6112
rect 32956 6060 33008 6112
rect 56416 6128 56468 6180
rect 43444 6060 43496 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 9128 5899 9180 5908
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 11060 5856 11112 5908
rect 7840 5788 7892 5840
rect 16580 5720 16632 5772
rect 940 5584 992 5636
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 9588 5695 9640 5704
rect 9588 5661 9597 5695
rect 9597 5661 9631 5695
rect 9631 5661 9640 5695
rect 9588 5652 9640 5661
rect 17684 5788 17736 5840
rect 23572 5899 23624 5908
rect 23572 5865 23581 5899
rect 23581 5865 23615 5899
rect 23615 5865 23624 5899
rect 23572 5856 23624 5865
rect 23940 5856 23992 5908
rect 25780 5899 25832 5908
rect 25780 5865 25789 5899
rect 25789 5865 25823 5899
rect 25823 5865 25832 5899
rect 25780 5856 25832 5865
rect 26056 5856 26108 5908
rect 30380 5856 30432 5908
rect 17316 5652 17368 5704
rect 10048 5584 10100 5636
rect 10600 5584 10652 5636
rect 12716 5584 12768 5636
rect 18052 5652 18104 5704
rect 18420 5695 18472 5704
rect 18420 5661 18429 5695
rect 18429 5661 18463 5695
rect 18463 5661 18472 5695
rect 18420 5652 18472 5661
rect 10232 5516 10284 5568
rect 10324 5516 10376 5568
rect 14464 5516 14516 5568
rect 17868 5584 17920 5636
rect 19432 5584 19484 5636
rect 24492 5788 24544 5840
rect 20260 5584 20312 5636
rect 21088 5584 21140 5636
rect 23940 5720 23992 5772
rect 27712 5788 27764 5840
rect 28908 5788 28960 5840
rect 20996 5516 21048 5568
rect 21272 5516 21324 5568
rect 23848 5652 23900 5704
rect 26056 5720 26108 5772
rect 26424 5720 26476 5772
rect 25320 5652 25372 5704
rect 26976 5652 27028 5704
rect 28632 5652 28684 5704
rect 29644 5695 29696 5704
rect 29644 5661 29653 5695
rect 29653 5661 29687 5695
rect 29687 5661 29696 5695
rect 29644 5652 29696 5661
rect 30380 5652 30432 5704
rect 24124 5584 24176 5636
rect 26792 5584 26844 5636
rect 28816 5627 28868 5636
rect 28816 5593 28825 5627
rect 28825 5593 28859 5627
rect 28859 5593 28868 5627
rect 28816 5584 28868 5593
rect 24308 5516 24360 5568
rect 26056 5516 26108 5568
rect 31024 5856 31076 5908
rect 32772 5856 32824 5908
rect 33048 5856 33100 5908
rect 35532 5856 35584 5908
rect 35624 5856 35676 5908
rect 37648 5856 37700 5908
rect 30748 5831 30800 5840
rect 30748 5797 30757 5831
rect 30757 5797 30791 5831
rect 30791 5797 30800 5831
rect 30748 5788 30800 5797
rect 31300 5763 31352 5772
rect 31300 5729 31309 5763
rect 31309 5729 31343 5763
rect 31343 5729 31352 5763
rect 31300 5720 31352 5729
rect 35900 5720 35952 5772
rect 35992 5720 36044 5772
rect 36268 5720 36320 5772
rect 36820 5720 36872 5772
rect 37096 5720 37148 5772
rect 38384 5763 38436 5772
rect 38384 5729 38393 5763
rect 38393 5729 38427 5763
rect 38427 5729 38436 5763
rect 38384 5720 38436 5729
rect 31392 5652 31444 5704
rect 34060 5652 34112 5704
rect 35440 5652 35492 5704
rect 40040 5720 40092 5772
rect 58256 5788 58308 5840
rect 58992 5720 59044 5772
rect 34244 5516 34296 5568
rect 35164 5627 35216 5636
rect 35164 5593 35173 5627
rect 35173 5593 35207 5627
rect 35207 5593 35216 5627
rect 35164 5584 35216 5593
rect 36268 5584 36320 5636
rect 36728 5584 36780 5636
rect 35808 5516 35860 5568
rect 35992 5559 36044 5568
rect 35992 5525 36001 5559
rect 36001 5525 36035 5559
rect 36035 5525 36044 5559
rect 35992 5516 36044 5525
rect 36360 5559 36412 5568
rect 36360 5525 36369 5559
rect 36369 5525 36403 5559
rect 36403 5525 36412 5559
rect 36360 5516 36412 5525
rect 36820 5516 36872 5568
rect 38844 5584 38896 5636
rect 41420 5627 41472 5636
rect 41420 5593 41429 5627
rect 41429 5593 41463 5627
rect 41463 5593 41472 5627
rect 41420 5584 41472 5593
rect 38936 5516 38988 5568
rect 57888 5695 57940 5704
rect 57888 5661 57897 5695
rect 57897 5661 57931 5695
rect 57931 5661 57940 5695
rect 57888 5652 57940 5661
rect 58900 5652 58952 5704
rect 57152 5516 57204 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 9588 5312 9640 5364
rect 10232 5355 10284 5364
rect 10232 5321 10241 5355
rect 10241 5321 10275 5355
rect 10275 5321 10284 5355
rect 10232 5312 10284 5321
rect 11980 5312 12032 5364
rect 13912 5312 13964 5364
rect 15568 5312 15620 5364
rect 16028 5312 16080 5364
rect 8116 5176 8168 5228
rect 940 5108 992 5160
rect 10140 5176 10192 5228
rect 9496 5108 9548 5160
rect 10048 5108 10100 5160
rect 6092 5040 6144 5092
rect 10600 5151 10652 5160
rect 10600 5117 10609 5151
rect 10609 5117 10643 5151
rect 10643 5117 10652 5151
rect 10600 5108 10652 5117
rect 10876 5108 10928 5160
rect 12256 5176 12308 5228
rect 13360 5219 13412 5228
rect 13360 5185 13369 5219
rect 13369 5185 13403 5219
rect 13403 5185 13412 5219
rect 13360 5176 13412 5185
rect 13912 5176 13964 5228
rect 19248 5176 19300 5228
rect 11980 5040 12032 5092
rect 12072 5040 12124 5092
rect 16580 5040 16632 5092
rect 8392 5015 8444 5024
rect 8392 4981 8401 5015
rect 8401 4981 8435 5015
rect 8435 4981 8444 5015
rect 8392 4972 8444 4981
rect 13452 4972 13504 5024
rect 13544 4972 13596 5024
rect 16672 4972 16724 5024
rect 16948 4972 17000 5024
rect 18604 5108 18656 5160
rect 19892 5312 19944 5364
rect 20444 5312 20496 5364
rect 25136 5312 25188 5364
rect 25872 5312 25924 5364
rect 32864 5312 32916 5364
rect 19524 5176 19576 5228
rect 20352 5244 20404 5296
rect 26884 5244 26936 5296
rect 21824 5176 21876 5228
rect 22560 5219 22612 5228
rect 22560 5185 22569 5219
rect 22569 5185 22603 5219
rect 22603 5185 22612 5219
rect 22560 5176 22612 5185
rect 24216 5176 24268 5228
rect 26148 5176 26200 5228
rect 20076 5108 20128 5160
rect 20904 5108 20956 5160
rect 21180 5151 21232 5160
rect 21180 5117 21189 5151
rect 21189 5117 21223 5151
rect 21223 5117 21232 5151
rect 21180 5108 21232 5117
rect 22468 5108 22520 5160
rect 23572 5108 23624 5160
rect 20996 5040 21048 5092
rect 21088 5040 21140 5092
rect 35348 5312 35400 5364
rect 27528 5176 27580 5228
rect 28540 5176 28592 5228
rect 29184 5219 29236 5228
rect 29184 5185 29193 5219
rect 29193 5185 29227 5219
rect 29227 5185 29236 5219
rect 29184 5176 29236 5185
rect 28724 5108 28776 5160
rect 29092 5108 29144 5160
rect 30840 5219 30892 5228
rect 30840 5185 30849 5219
rect 30849 5185 30883 5219
rect 30883 5185 30892 5219
rect 30840 5176 30892 5185
rect 31852 5176 31904 5228
rect 34244 5176 34296 5228
rect 34428 5176 34480 5228
rect 35992 5244 36044 5296
rect 39580 5312 39632 5364
rect 43168 5312 43220 5364
rect 43904 5312 43956 5364
rect 53104 5312 53156 5364
rect 33140 5040 33192 5092
rect 34336 5040 34388 5092
rect 34612 5040 34664 5092
rect 34980 5151 35032 5160
rect 34980 5117 34989 5151
rect 34989 5117 35023 5151
rect 35023 5117 35032 5151
rect 34980 5108 35032 5117
rect 36268 5176 36320 5228
rect 38016 5176 38068 5228
rect 39120 5176 39172 5228
rect 39212 5176 39264 5228
rect 40500 5176 40552 5228
rect 41880 5176 41932 5228
rect 42892 5176 42944 5228
rect 44180 5219 44232 5228
rect 44180 5185 44189 5219
rect 44189 5185 44223 5219
rect 44223 5185 44232 5219
rect 44180 5176 44232 5185
rect 44548 5176 44600 5228
rect 45652 5176 45704 5228
rect 46940 5176 46992 5228
rect 35348 5108 35400 5160
rect 35440 5040 35492 5092
rect 35716 5108 35768 5160
rect 37004 5108 37056 5160
rect 40592 5108 40644 5160
rect 46572 5108 46624 5160
rect 58072 5219 58124 5228
rect 58072 5185 58081 5219
rect 58081 5185 58115 5219
rect 58115 5185 58124 5219
rect 58072 5176 58124 5185
rect 37740 5040 37792 5092
rect 41236 5040 41288 5092
rect 20720 4972 20772 5024
rect 20904 4972 20956 5024
rect 23480 4972 23532 5024
rect 23848 4972 23900 5024
rect 26240 4972 26292 5024
rect 27528 4972 27580 5024
rect 28172 4972 28224 5024
rect 34796 4972 34848 5024
rect 35992 4972 36044 5024
rect 38660 4972 38712 5024
rect 38844 4972 38896 5024
rect 41144 4972 41196 5024
rect 43076 4972 43128 5024
rect 45008 5015 45060 5024
rect 45008 4981 45017 5015
rect 45017 4981 45051 5015
rect 45051 4981 45060 5015
rect 45008 4972 45060 4981
rect 51080 4972 51132 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 8116 4768 8168 4820
rect 11244 4768 11296 4820
rect 16120 4768 16172 4820
rect 19340 4768 19392 4820
rect 19524 4768 19576 4820
rect 7104 4743 7156 4752
rect 7104 4709 7113 4743
rect 7113 4709 7147 4743
rect 7147 4709 7156 4743
rect 7104 4700 7156 4709
rect 13452 4743 13504 4752
rect 13452 4709 13461 4743
rect 13461 4709 13495 4743
rect 13495 4709 13504 4743
rect 13452 4700 13504 4709
rect 9772 4632 9824 4684
rect 9864 4675 9916 4684
rect 9864 4641 9873 4675
rect 9873 4641 9907 4675
rect 9907 4641 9916 4675
rect 9864 4632 9916 4641
rect 7012 4564 7064 4616
rect 9680 4564 9732 4616
rect 10048 4607 10100 4616
rect 10048 4573 10057 4607
rect 10057 4573 10091 4607
rect 10091 4573 10100 4607
rect 10048 4564 10100 4573
rect 5908 4496 5960 4548
rect 8300 4496 8352 4548
rect 8576 4496 8628 4548
rect 10600 4564 10652 4616
rect 12716 4564 12768 4616
rect 13360 4632 13412 4684
rect 14556 4743 14608 4752
rect 14556 4709 14565 4743
rect 14565 4709 14599 4743
rect 14599 4709 14608 4743
rect 14556 4700 14608 4709
rect 15292 4632 15344 4684
rect 15200 4564 15252 4616
rect 15384 4607 15436 4616
rect 15384 4573 15393 4607
rect 15393 4573 15427 4607
rect 15427 4573 15436 4607
rect 15384 4564 15436 4573
rect 13084 4496 13136 4548
rect 7564 4428 7616 4480
rect 11980 4428 12032 4480
rect 14188 4496 14240 4548
rect 15292 4496 15344 4548
rect 17224 4564 17276 4616
rect 19616 4700 19668 4752
rect 20076 4700 20128 4752
rect 21088 4700 21140 4752
rect 19064 4564 19116 4616
rect 19340 4564 19392 4616
rect 21272 4675 21324 4684
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 33508 4768 33560 4820
rect 36360 4768 36412 4820
rect 37372 4768 37424 4820
rect 38844 4768 38896 4820
rect 39120 4811 39172 4820
rect 39120 4777 39129 4811
rect 39129 4777 39163 4811
rect 39163 4777 39172 4811
rect 39120 4768 39172 4777
rect 40224 4811 40276 4820
rect 40224 4777 40233 4811
rect 40233 4777 40267 4811
rect 40267 4777 40276 4811
rect 40224 4768 40276 4777
rect 40684 4768 40736 4820
rect 29644 4700 29696 4752
rect 23848 4675 23900 4684
rect 23848 4641 23857 4675
rect 23857 4641 23891 4675
rect 23891 4641 23900 4675
rect 23848 4632 23900 4641
rect 24952 4675 25004 4684
rect 20260 4564 20312 4616
rect 22376 4607 22428 4616
rect 22376 4573 22385 4607
rect 22385 4573 22419 4607
rect 22419 4573 22428 4607
rect 22376 4564 22428 4573
rect 24952 4641 24961 4675
rect 24961 4641 24995 4675
rect 24995 4641 25004 4675
rect 24952 4632 25004 4641
rect 27620 4675 27672 4684
rect 27620 4641 27629 4675
rect 27629 4641 27663 4675
rect 27663 4641 27672 4675
rect 27620 4632 27672 4641
rect 24676 4607 24728 4616
rect 24676 4573 24685 4607
rect 24685 4573 24719 4607
rect 24719 4573 24728 4607
rect 24676 4564 24728 4573
rect 26332 4564 26384 4616
rect 27804 4607 27856 4616
rect 27804 4573 27813 4607
rect 27813 4573 27847 4607
rect 27847 4573 27856 4607
rect 27804 4564 27856 4573
rect 18052 4496 18104 4548
rect 19156 4496 19208 4548
rect 19248 4496 19300 4548
rect 20352 4496 20404 4548
rect 22560 4496 22612 4548
rect 22744 4496 22796 4548
rect 23940 4496 23992 4548
rect 28724 4632 28776 4684
rect 29460 4632 29512 4684
rect 32864 4675 32916 4684
rect 32864 4641 32873 4675
rect 32873 4641 32907 4675
rect 32907 4641 32916 4675
rect 32864 4632 32916 4641
rect 36912 4700 36964 4752
rect 37832 4700 37884 4752
rect 38016 4700 38068 4752
rect 29000 4564 29052 4616
rect 29184 4564 29236 4616
rect 30012 4539 30064 4548
rect 30012 4505 30021 4539
rect 30021 4505 30055 4539
rect 30055 4505 30064 4539
rect 30012 4496 30064 4505
rect 30288 4496 30340 4548
rect 32956 4564 33008 4616
rect 39120 4632 39172 4684
rect 41052 4632 41104 4684
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 14832 4428 14884 4480
rect 20444 4428 20496 4480
rect 20628 4471 20680 4480
rect 20628 4437 20637 4471
rect 20637 4437 20671 4471
rect 20671 4437 20680 4471
rect 20628 4428 20680 4437
rect 21180 4428 21232 4480
rect 23480 4428 23532 4480
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 23756 4428 23808 4437
rect 26884 4428 26936 4480
rect 28540 4428 28592 4480
rect 28724 4428 28776 4480
rect 33140 4496 33192 4548
rect 34520 4564 34572 4616
rect 37004 4564 37056 4616
rect 37740 4607 37792 4616
rect 37740 4573 37749 4607
rect 37749 4573 37783 4607
rect 37783 4573 37792 4607
rect 37740 4564 37792 4573
rect 37832 4607 37884 4616
rect 37832 4573 37841 4607
rect 37841 4573 37875 4607
rect 37875 4573 37884 4607
rect 37832 4564 37884 4573
rect 38936 4607 38988 4616
rect 38936 4573 38945 4607
rect 38945 4573 38979 4607
rect 38979 4573 38988 4607
rect 38936 4564 38988 4573
rect 40040 4607 40092 4616
rect 40040 4573 40049 4607
rect 40049 4573 40083 4607
rect 40083 4573 40092 4607
rect 40040 4564 40092 4573
rect 40224 4564 40276 4616
rect 33784 4496 33836 4548
rect 34060 4496 34112 4548
rect 34428 4496 34480 4548
rect 35348 4496 35400 4548
rect 35992 4539 36044 4548
rect 35992 4505 36026 4539
rect 36026 4505 36044 4539
rect 35992 4496 36044 4505
rect 36360 4496 36412 4548
rect 39028 4496 39080 4548
rect 40868 4539 40920 4548
rect 40868 4505 40877 4539
rect 40877 4505 40911 4539
rect 40911 4505 40920 4539
rect 40868 4496 40920 4505
rect 33508 4428 33560 4480
rect 33600 4428 33652 4480
rect 36268 4428 36320 4480
rect 36728 4428 36780 4480
rect 38016 4471 38068 4480
rect 38016 4437 38025 4471
rect 38025 4437 38059 4471
rect 38059 4437 38068 4471
rect 38016 4428 38068 4437
rect 38844 4428 38896 4480
rect 42708 4607 42760 4616
rect 42708 4573 42717 4607
rect 42717 4573 42751 4607
rect 42751 4573 42760 4607
rect 42708 4564 42760 4573
rect 43260 4700 43312 4752
rect 45468 4743 45520 4752
rect 45468 4709 45477 4743
rect 45477 4709 45511 4743
rect 45511 4709 45520 4743
rect 45468 4700 45520 4709
rect 56692 4768 56744 4820
rect 51356 4700 51408 4752
rect 43076 4607 43128 4616
rect 43076 4573 43085 4607
rect 43085 4573 43119 4607
rect 43119 4573 43128 4607
rect 43076 4564 43128 4573
rect 43444 4564 43496 4616
rect 43904 4607 43956 4616
rect 43904 4573 43913 4607
rect 43913 4573 43947 4607
rect 43947 4573 43956 4607
rect 43904 4564 43956 4573
rect 43996 4564 44048 4616
rect 49608 4632 49660 4684
rect 42984 4539 43036 4548
rect 42984 4505 42993 4539
rect 42993 4505 43027 4539
rect 43027 4505 43036 4539
rect 42984 4496 43036 4505
rect 43352 4471 43404 4480
rect 43352 4437 43361 4471
rect 43361 4437 43395 4471
rect 43395 4437 43404 4471
rect 43352 4428 43404 4437
rect 51080 4607 51132 4616
rect 51080 4573 51089 4607
rect 51089 4573 51123 4607
rect 51123 4573 51132 4607
rect 51080 4564 51132 4573
rect 58808 4564 58860 4616
rect 44456 4496 44508 4548
rect 46020 4539 46072 4548
rect 46020 4505 46029 4539
rect 46029 4505 46063 4539
rect 46063 4505 46072 4539
rect 46020 4496 46072 4505
rect 53748 4428 53800 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 6460 4156 6512 4208
rect 5724 4088 5776 4140
rect 940 4020 992 4072
rect 8852 4224 8904 4276
rect 11152 4224 11204 4276
rect 14556 4224 14608 4276
rect 15200 4224 15252 4276
rect 21180 4267 21232 4276
rect 21180 4233 21189 4267
rect 21189 4233 21223 4267
rect 21223 4233 21232 4267
rect 21180 4224 21232 4233
rect 24676 4224 24728 4276
rect 9312 4156 9364 4208
rect 11704 4156 11756 4208
rect 12348 4156 12400 4208
rect 13360 4199 13412 4208
rect 13360 4165 13369 4199
rect 13369 4165 13403 4199
rect 13403 4165 13412 4199
rect 13360 4156 13412 4165
rect 8208 4088 8260 4140
rect 8392 4088 8444 4140
rect 8116 4020 8168 4072
rect 8944 4063 8996 4072
rect 8944 4029 8953 4063
rect 8953 4029 8987 4063
rect 8987 4029 8996 4063
rect 8944 4020 8996 4029
rect 9128 4063 9180 4072
rect 9128 4029 9137 4063
rect 9137 4029 9171 4063
rect 9171 4029 9180 4063
rect 9128 4020 9180 4029
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 9496 4020 9548 4072
rect 10416 4063 10468 4072
rect 10416 4029 10425 4063
rect 10425 4029 10459 4063
rect 10459 4029 10468 4063
rect 10416 4020 10468 4029
rect 6000 3995 6052 4004
rect 6000 3961 6009 3995
rect 6009 3961 6043 3995
rect 6043 3961 6052 3995
rect 6000 3952 6052 3961
rect 7472 3927 7524 3936
rect 7472 3893 7481 3927
rect 7481 3893 7515 3927
rect 7515 3893 7524 3927
rect 7472 3884 7524 3893
rect 8392 3995 8444 4004
rect 8392 3961 8401 3995
rect 8401 3961 8435 3995
rect 8435 3961 8444 3995
rect 8392 3952 8444 3961
rect 9772 3952 9824 4004
rect 8668 3884 8720 3936
rect 9404 3884 9456 3936
rect 11244 4088 11296 4140
rect 12900 4063 12952 4072
rect 12900 4029 12909 4063
rect 12909 4029 12943 4063
rect 12943 4029 12952 4063
rect 12900 4020 12952 4029
rect 12716 3995 12768 4004
rect 12716 3961 12725 3995
rect 12725 3961 12759 3995
rect 12759 3961 12768 3995
rect 12716 3952 12768 3961
rect 14924 4020 14976 4072
rect 15844 4020 15896 4072
rect 16120 4020 16172 4072
rect 17132 4088 17184 4140
rect 19892 4156 19944 4208
rect 20628 4156 20680 4208
rect 20720 4156 20772 4208
rect 28356 4224 28408 4276
rect 29552 4224 29604 4276
rect 27160 4156 27212 4208
rect 27436 4156 27488 4208
rect 18144 4088 18196 4140
rect 18972 4088 19024 4140
rect 13728 3952 13780 4004
rect 14832 3952 14884 4004
rect 17316 4063 17368 4072
rect 17316 4029 17325 4063
rect 17325 4029 17359 4063
rect 17359 4029 17368 4063
rect 17316 4020 17368 4029
rect 15936 3927 15988 3936
rect 15936 3893 15945 3927
rect 15945 3893 15979 3927
rect 15979 3893 15988 3927
rect 15936 3884 15988 3893
rect 17960 3952 18012 4004
rect 18972 3884 19024 3936
rect 19248 4020 19300 4072
rect 19708 4088 19760 4140
rect 20444 4088 20496 4140
rect 22652 4088 22704 4140
rect 23296 4088 23348 4140
rect 23480 4088 23532 4140
rect 25228 4131 25280 4140
rect 25228 4097 25237 4131
rect 25237 4097 25271 4131
rect 25271 4097 25280 4131
rect 25228 4088 25280 4097
rect 23112 4020 23164 4072
rect 24676 4020 24728 4072
rect 20076 3884 20128 3936
rect 20720 3884 20772 3936
rect 27344 4088 27396 4140
rect 27528 4131 27580 4140
rect 27528 4097 27562 4131
rect 27562 4097 27580 4131
rect 27528 4088 27580 4097
rect 27896 4088 27948 4140
rect 30748 4199 30800 4208
rect 30748 4165 30757 4199
rect 30757 4165 30791 4199
rect 30791 4165 30800 4199
rect 30748 4156 30800 4165
rect 31116 4156 31168 4208
rect 33324 4224 33376 4276
rect 34244 4224 34296 4276
rect 37372 4224 37424 4276
rect 37832 4224 37884 4276
rect 34612 4156 34664 4208
rect 37740 4156 37792 4208
rect 38108 4224 38160 4276
rect 38200 4156 38252 4208
rect 42064 4224 42116 4276
rect 43352 4224 43404 4276
rect 53104 4267 53156 4276
rect 53104 4233 53113 4267
rect 53113 4233 53147 4267
rect 53147 4233 53156 4267
rect 53104 4224 53156 4233
rect 35348 4131 35400 4140
rect 35348 4097 35357 4131
rect 35357 4097 35391 4131
rect 35391 4097 35400 4131
rect 35348 4088 35400 4097
rect 35900 4088 35952 4140
rect 37832 4131 37884 4140
rect 37832 4097 37841 4131
rect 37841 4097 37875 4131
rect 37875 4097 37884 4131
rect 37832 4088 37884 4097
rect 39396 4088 39448 4140
rect 44824 4156 44876 4208
rect 52000 4156 52052 4208
rect 52828 4156 52880 4208
rect 53380 4156 53432 4208
rect 58992 4156 59044 4208
rect 29644 4020 29696 4072
rect 32588 4020 32640 4072
rect 32864 4063 32916 4072
rect 32864 4029 32873 4063
rect 32873 4029 32907 4063
rect 32907 4029 32916 4063
rect 32864 4020 32916 4029
rect 33140 4020 33192 4072
rect 34612 4063 34664 4072
rect 34612 4029 34621 4063
rect 34621 4029 34655 4063
rect 34655 4029 34664 4063
rect 34612 4020 34664 4029
rect 34704 4020 34756 4072
rect 35624 4020 35676 4072
rect 32128 3952 32180 4004
rect 28448 3884 28500 3936
rect 28632 3927 28684 3936
rect 28632 3893 28641 3927
rect 28641 3893 28675 3927
rect 28675 3893 28684 3927
rect 28632 3884 28684 3893
rect 30840 3927 30892 3936
rect 30840 3893 30849 3927
rect 30849 3893 30883 3927
rect 30883 3893 30892 3927
rect 30840 3884 30892 3893
rect 31576 3884 31628 3936
rect 39856 4020 39908 4072
rect 38200 3952 38252 4004
rect 40132 4088 40184 4140
rect 41604 4131 41656 4140
rect 41604 4097 41613 4131
rect 41613 4097 41647 4131
rect 41647 4097 41656 4131
rect 41604 4088 41656 4097
rect 42064 4088 42116 4140
rect 42984 4088 43036 4140
rect 44272 4088 44324 4140
rect 44916 4088 44968 4140
rect 42616 4063 42668 4072
rect 42616 4029 42625 4063
rect 42625 4029 42659 4063
rect 42659 4029 42668 4063
rect 42616 4020 42668 4029
rect 43076 4063 43128 4072
rect 43076 4029 43085 4063
rect 43085 4029 43119 4063
rect 43119 4029 43128 4063
rect 43076 4020 43128 4029
rect 43444 4020 43496 4072
rect 43996 4020 44048 4072
rect 45928 4088 45980 4140
rect 46756 4131 46808 4140
rect 46756 4097 46765 4131
rect 46765 4097 46799 4131
rect 46799 4097 46808 4131
rect 46756 4088 46808 4097
rect 48136 4088 48188 4140
rect 52368 4088 52420 4140
rect 54484 4088 54536 4140
rect 46388 4020 46440 4072
rect 40408 3952 40460 4004
rect 41696 3952 41748 4004
rect 47952 3952 48004 4004
rect 48412 3995 48464 4004
rect 48412 3961 48421 3995
rect 48421 3961 48455 3995
rect 48455 3961 48464 3995
rect 48412 3952 48464 3961
rect 52276 4020 52328 4072
rect 43628 3884 43680 3936
rect 45192 3927 45244 3936
rect 45192 3893 45201 3927
rect 45201 3893 45235 3927
rect 45235 3893 45244 3927
rect 45192 3884 45244 3893
rect 52276 3927 52328 3936
rect 52276 3893 52285 3927
rect 52285 3893 52319 3927
rect 52319 3893 52328 3927
rect 52276 3884 52328 3893
rect 53656 3952 53708 4004
rect 57428 3884 57480 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 7472 3680 7524 3732
rect 5264 3655 5316 3664
rect 5264 3621 5273 3655
rect 5273 3621 5307 3655
rect 5307 3621 5316 3655
rect 5264 3612 5316 3621
rect 6184 3612 6236 3664
rect 7564 3655 7616 3664
rect 7564 3621 7573 3655
rect 7573 3621 7607 3655
rect 7607 3621 7616 3655
rect 7564 3612 7616 3621
rect 8576 3655 8628 3664
rect 8576 3621 8585 3655
rect 8585 3621 8619 3655
rect 8619 3621 8628 3655
rect 8576 3612 8628 3621
rect 10876 3723 10928 3732
rect 10876 3689 10885 3723
rect 10885 3689 10919 3723
rect 10919 3689 10928 3723
rect 10876 3680 10928 3689
rect 11060 3680 11112 3732
rect 13728 3680 13780 3732
rect 12072 3655 12124 3664
rect 12072 3621 12081 3655
rect 12081 3621 12115 3655
rect 12115 3621 12124 3655
rect 12072 3612 12124 3621
rect 12532 3612 12584 3664
rect 14188 3612 14240 3664
rect 14648 3612 14700 3664
rect 14096 3544 14148 3596
rect 15200 3544 15252 3596
rect 15844 3544 15896 3596
rect 23756 3680 23808 3732
rect 24952 3680 25004 3732
rect 25320 3680 25372 3732
rect 27252 3680 27304 3732
rect 27804 3723 27856 3732
rect 27804 3689 27813 3723
rect 27813 3689 27847 3723
rect 27847 3689 27856 3723
rect 27804 3680 27856 3689
rect 28448 3680 28500 3732
rect 31300 3680 31352 3732
rect 33324 3680 33376 3732
rect 36636 3680 36688 3732
rect 9588 3519 9640 3528
rect 9588 3485 9597 3519
rect 9597 3485 9631 3519
rect 9631 3485 9640 3519
rect 9588 3476 9640 3485
rect 940 3408 992 3460
rect 5080 3451 5132 3460
rect 5080 3417 5089 3451
rect 5089 3417 5123 3451
rect 5123 3417 5132 3451
rect 5080 3408 5132 3417
rect 7104 3408 7156 3460
rect 8208 3408 8260 3460
rect 7288 3340 7340 3392
rect 9496 3408 9548 3460
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 14832 3476 14884 3528
rect 16764 3476 16816 3528
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 18512 3476 18564 3485
rect 19064 3544 19116 3596
rect 19432 3544 19484 3596
rect 19708 3587 19760 3596
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 30472 3612 30524 3664
rect 25136 3587 25188 3596
rect 25136 3553 25145 3587
rect 25145 3553 25179 3587
rect 25179 3553 25188 3587
rect 25136 3544 25188 3553
rect 21916 3476 21968 3528
rect 22652 3519 22704 3528
rect 22652 3485 22661 3519
rect 22661 3485 22695 3519
rect 22695 3485 22704 3519
rect 22652 3476 22704 3485
rect 23296 3476 23348 3528
rect 23848 3476 23900 3528
rect 25780 3519 25832 3528
rect 25780 3485 25789 3519
rect 25789 3485 25823 3519
rect 25823 3485 25832 3519
rect 25780 3476 25832 3485
rect 27988 3544 28040 3596
rect 28264 3587 28316 3596
rect 28264 3553 28273 3587
rect 28273 3553 28307 3587
rect 28307 3553 28316 3587
rect 28264 3544 28316 3553
rect 28816 3544 28868 3596
rect 31300 3544 31352 3596
rect 33416 3544 33468 3596
rect 34612 3544 34664 3596
rect 9312 3340 9364 3392
rect 12624 3451 12676 3460
rect 12624 3417 12633 3451
rect 12633 3417 12667 3451
rect 12667 3417 12676 3451
rect 12624 3408 12676 3417
rect 13268 3451 13320 3460
rect 13268 3417 13277 3451
rect 13277 3417 13311 3451
rect 13311 3417 13320 3451
rect 13268 3408 13320 3417
rect 17500 3451 17552 3460
rect 17500 3417 17509 3451
rect 17509 3417 17543 3451
rect 17543 3417 17552 3451
rect 17500 3408 17552 3417
rect 13360 3340 13412 3392
rect 19340 3340 19392 3392
rect 22008 3451 22060 3460
rect 22008 3417 22017 3451
rect 22017 3417 22051 3451
rect 22051 3417 22060 3451
rect 22008 3408 22060 3417
rect 23204 3408 23256 3460
rect 26792 3451 26844 3460
rect 26792 3417 26801 3451
rect 26801 3417 26835 3451
rect 26835 3417 26844 3451
rect 26792 3408 26844 3417
rect 26976 3451 27028 3460
rect 26976 3417 26985 3451
rect 26985 3417 27019 3451
rect 27019 3417 27028 3451
rect 26976 3408 27028 3417
rect 27344 3519 27396 3528
rect 27344 3485 27353 3519
rect 27353 3485 27387 3519
rect 27387 3485 27396 3519
rect 27344 3476 27396 3485
rect 28632 3476 28684 3528
rect 30288 3519 30340 3528
rect 30288 3485 30297 3519
rect 30297 3485 30331 3519
rect 30331 3485 30340 3519
rect 30288 3476 30340 3485
rect 30932 3476 30984 3528
rect 31576 3519 31628 3528
rect 31576 3485 31585 3519
rect 31585 3485 31619 3519
rect 31619 3485 31628 3519
rect 31576 3476 31628 3485
rect 34796 3476 34848 3528
rect 35900 3519 35952 3528
rect 35900 3485 35909 3519
rect 35909 3485 35943 3519
rect 35943 3485 35952 3519
rect 35900 3476 35952 3485
rect 37004 3587 37056 3596
rect 37004 3553 37013 3587
rect 37013 3553 37047 3587
rect 37047 3553 37056 3587
rect 37004 3544 37056 3553
rect 38016 3544 38068 3596
rect 38200 3680 38252 3732
rect 40868 3680 40920 3732
rect 41052 3680 41104 3732
rect 41696 3680 41748 3732
rect 38292 3612 38344 3664
rect 39028 3612 39080 3664
rect 40224 3612 40276 3664
rect 40408 3655 40460 3664
rect 40408 3621 40417 3655
rect 40417 3621 40451 3655
rect 40451 3621 40460 3655
rect 40408 3612 40460 3621
rect 42708 3680 42760 3732
rect 44272 3680 44324 3732
rect 45560 3680 45612 3732
rect 47032 3723 47084 3732
rect 47032 3689 47041 3723
rect 47041 3689 47075 3723
rect 47075 3689 47084 3723
rect 47032 3680 47084 3689
rect 47952 3723 48004 3732
rect 47952 3689 47961 3723
rect 47961 3689 47995 3723
rect 47995 3689 48004 3723
rect 47952 3680 48004 3689
rect 48596 3680 48648 3732
rect 49424 3723 49476 3732
rect 49424 3689 49433 3723
rect 49433 3689 49467 3723
rect 49467 3689 49476 3723
rect 49424 3680 49476 3689
rect 50160 3680 50212 3732
rect 51356 3680 51408 3732
rect 54208 3723 54260 3732
rect 54208 3689 54217 3723
rect 54217 3689 54251 3723
rect 54251 3689 54260 3723
rect 54208 3680 54260 3689
rect 40592 3544 40644 3596
rect 42156 3612 42208 3664
rect 41328 3544 41380 3596
rect 36912 3476 36964 3528
rect 27988 3408 28040 3460
rect 30196 3408 30248 3460
rect 33232 3408 33284 3460
rect 38844 3476 38896 3528
rect 40776 3519 40828 3528
rect 40776 3485 40785 3519
rect 40785 3485 40819 3519
rect 40819 3485 40828 3519
rect 40776 3476 40828 3485
rect 41144 3519 41196 3528
rect 41144 3485 41153 3519
rect 41153 3485 41187 3519
rect 41187 3485 41196 3519
rect 41144 3476 41196 3485
rect 41236 3519 41288 3528
rect 41236 3485 41245 3519
rect 41245 3485 41279 3519
rect 41279 3485 41288 3519
rect 41236 3476 41288 3485
rect 43444 3476 43496 3528
rect 45008 3612 45060 3664
rect 45100 3612 45152 3664
rect 46020 3612 46072 3664
rect 48320 3612 48372 3664
rect 53840 3612 53892 3664
rect 43720 3519 43772 3528
rect 43720 3485 43729 3519
rect 43729 3485 43763 3519
rect 43763 3485 43772 3519
rect 43720 3476 43772 3485
rect 52276 3544 52328 3596
rect 56876 3587 56928 3596
rect 56876 3553 56885 3587
rect 56885 3553 56919 3587
rect 56919 3553 56928 3587
rect 56876 3544 56928 3553
rect 24032 3383 24084 3392
rect 24032 3349 24041 3383
rect 24041 3349 24075 3383
rect 24075 3349 24084 3383
rect 24032 3340 24084 3349
rect 25044 3383 25096 3392
rect 25044 3349 25053 3383
rect 25053 3349 25087 3383
rect 25087 3349 25096 3383
rect 25044 3340 25096 3349
rect 25136 3340 25188 3392
rect 26056 3340 26108 3392
rect 27252 3340 27304 3392
rect 29736 3340 29788 3392
rect 31024 3340 31076 3392
rect 32588 3340 32640 3392
rect 34796 3340 34848 3392
rect 35624 3340 35676 3392
rect 39120 3408 39172 3460
rect 39396 3408 39448 3460
rect 37924 3340 37976 3392
rect 38844 3340 38896 3392
rect 42984 3340 43036 3392
rect 43904 3408 43956 3460
rect 46112 3476 46164 3528
rect 47584 3476 47636 3528
rect 48688 3476 48740 3528
rect 51264 3476 51316 3528
rect 53104 3476 53156 3528
rect 54760 3476 54812 3528
rect 44732 3408 44784 3460
rect 45376 3408 45428 3460
rect 43720 3340 43772 3392
rect 44180 3340 44232 3392
rect 46756 3408 46808 3460
rect 49792 3408 49844 3460
rect 50620 3408 50672 3460
rect 51724 3408 51776 3460
rect 51080 3340 51132 3392
rect 52368 3340 52420 3392
rect 53748 3408 53800 3460
rect 53472 3383 53524 3392
rect 53472 3349 53481 3383
rect 53481 3349 53515 3383
rect 53515 3349 53524 3383
rect 53472 3340 53524 3349
rect 57244 3340 57296 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 5816 3136 5868 3188
rect 5172 3068 5224 3120
rect 6092 3136 6144 3188
rect 7104 3136 7156 3188
rect 8576 3136 8628 3188
rect 9864 3136 9916 3188
rect 12532 3179 12584 3188
rect 12532 3145 12541 3179
rect 12541 3145 12575 3179
rect 12575 3145 12584 3179
rect 12532 3136 12584 3145
rect 13176 3136 13228 3188
rect 940 2932 992 2984
rect 7656 3000 7708 3052
rect 8024 3000 8076 3052
rect 7564 2932 7616 2984
rect 8208 3068 8260 3120
rect 9220 3000 9272 3052
rect 8668 2907 8720 2916
rect 8668 2873 8677 2907
rect 8677 2873 8711 2907
rect 8711 2873 8720 2907
rect 8668 2864 8720 2873
rect 9312 2975 9364 2984
rect 9312 2941 9321 2975
rect 9321 2941 9355 2975
rect 9355 2941 9364 2975
rect 9312 2932 9364 2941
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 13728 3000 13780 3052
rect 13268 2932 13320 2984
rect 13544 2932 13596 2984
rect 15568 3136 15620 3188
rect 19064 3136 19116 3188
rect 20352 3136 20404 3188
rect 20444 3136 20496 3188
rect 23204 3136 23256 3188
rect 23664 3179 23716 3188
rect 23664 3145 23673 3179
rect 23673 3145 23707 3179
rect 23707 3145 23716 3179
rect 23664 3136 23716 3145
rect 25044 3136 25096 3188
rect 34244 3136 34296 3188
rect 34336 3136 34388 3188
rect 37648 3136 37700 3188
rect 39396 3136 39448 3188
rect 39764 3179 39816 3188
rect 39764 3145 39773 3179
rect 39773 3145 39807 3179
rect 39807 3145 39816 3179
rect 39764 3136 39816 3145
rect 40316 3136 40368 3188
rect 41788 3179 41840 3188
rect 41788 3145 41797 3179
rect 41797 3145 41831 3179
rect 41831 3145 41840 3179
rect 41788 3136 41840 3145
rect 44364 3136 44416 3188
rect 44640 3136 44692 3188
rect 47492 3136 47544 3188
rect 48780 3136 48832 3188
rect 49884 3136 49936 3188
rect 52184 3179 52236 3188
rect 52184 3145 52193 3179
rect 52193 3145 52227 3179
rect 52227 3145 52236 3179
rect 52184 3136 52236 3145
rect 54024 3136 54076 3188
rect 55220 3136 55272 3188
rect 57428 3179 57480 3188
rect 57428 3145 57437 3179
rect 57437 3145 57471 3179
rect 57471 3145 57480 3179
rect 57428 3136 57480 3145
rect 24032 3068 24084 3120
rect 28540 3068 28592 3120
rect 31300 3068 31352 3120
rect 14464 3000 14516 3052
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 15844 3043 15896 3052
rect 15844 3009 15853 3043
rect 15853 3009 15887 3043
rect 15887 3009 15896 3043
rect 15844 3000 15896 3009
rect 6920 2796 6972 2848
rect 7380 2796 7432 2848
rect 7932 2796 7984 2848
rect 8024 2796 8076 2848
rect 10876 2796 10928 2848
rect 14832 2796 14884 2848
rect 16028 2932 16080 2984
rect 16304 2932 16356 2984
rect 17592 2932 17644 2984
rect 17868 3043 17920 3052
rect 17868 3009 17877 3043
rect 17877 3009 17911 3043
rect 17911 3009 17920 3043
rect 17868 3000 17920 3009
rect 18696 3000 18748 3052
rect 19432 3000 19484 3052
rect 19984 3043 20036 3052
rect 19984 3009 20018 3043
rect 20018 3009 20036 3043
rect 19984 3000 20036 3009
rect 20352 3000 20404 3052
rect 21272 3000 21324 3052
rect 22836 3000 22888 3052
rect 17960 2932 18012 2984
rect 18144 2975 18196 2984
rect 18144 2941 18153 2975
rect 18153 2941 18187 2975
rect 18187 2941 18196 2975
rect 18144 2932 18196 2941
rect 18972 2975 19024 2984
rect 18972 2941 18981 2975
rect 18981 2941 19015 2975
rect 19015 2941 19024 2975
rect 18972 2932 19024 2941
rect 23388 2932 23440 2984
rect 23940 2975 23992 2984
rect 23940 2941 23949 2975
rect 23949 2941 23983 2975
rect 23983 2941 23992 2975
rect 23940 2932 23992 2941
rect 17500 2864 17552 2916
rect 19432 2864 19484 2916
rect 24952 2864 25004 2916
rect 25228 2864 25280 2916
rect 26976 3000 27028 3052
rect 27528 3043 27580 3052
rect 27528 3009 27537 3043
rect 27537 3009 27571 3043
rect 27571 3009 27580 3043
rect 27528 3000 27580 3009
rect 28448 3043 28500 3052
rect 28448 3009 28457 3043
rect 28457 3009 28491 3043
rect 28491 3009 28500 3043
rect 28448 3000 28500 3009
rect 30840 3043 30892 3052
rect 30840 3009 30849 3043
rect 30849 3009 30883 3043
rect 30883 3009 30892 3043
rect 30840 3000 30892 3009
rect 37924 3111 37976 3120
rect 37924 3077 37933 3111
rect 37933 3077 37967 3111
rect 37967 3077 37976 3111
rect 37924 3068 37976 3077
rect 38568 3068 38620 3120
rect 41052 3068 41104 3120
rect 42616 3111 42668 3120
rect 42616 3077 42625 3111
rect 42625 3077 42659 3111
rect 42659 3077 42668 3111
rect 42616 3068 42668 3077
rect 43168 3068 43220 3120
rect 44916 3068 44968 3120
rect 47124 3068 47176 3120
rect 49516 3068 49568 3120
rect 50896 3068 50948 3120
rect 53288 3068 53340 3120
rect 58164 3111 58216 3120
rect 58164 3077 58173 3111
rect 58173 3077 58207 3111
rect 58207 3077 58216 3111
rect 58164 3068 58216 3077
rect 27344 2932 27396 2984
rect 27804 2975 27856 2984
rect 27804 2941 27813 2975
rect 27813 2941 27847 2975
rect 27847 2941 27856 2975
rect 27804 2932 27856 2941
rect 30564 2932 30616 2984
rect 30748 2932 30800 2984
rect 29736 2864 29788 2916
rect 30104 2864 30156 2916
rect 34520 3000 34572 3052
rect 35440 3043 35492 3052
rect 35440 3009 35449 3043
rect 35449 3009 35483 3043
rect 35483 3009 35492 3043
rect 35440 3000 35492 3009
rect 36176 3000 36228 3052
rect 37280 3000 37332 3052
rect 38660 3043 38712 3052
rect 38660 3009 38669 3043
rect 38669 3009 38703 3043
rect 38703 3009 38712 3043
rect 38660 3000 38712 3009
rect 31576 2932 31628 2984
rect 33600 2975 33652 2984
rect 33600 2941 33609 2975
rect 33609 2941 33643 2975
rect 33643 2941 33652 2975
rect 33600 2932 33652 2941
rect 35624 2975 35676 2984
rect 35624 2941 35633 2975
rect 35633 2941 35667 2975
rect 35667 2941 35676 2975
rect 35624 2932 35676 2941
rect 36544 2975 36596 2984
rect 36544 2941 36553 2975
rect 36553 2941 36587 2975
rect 36587 2941 36596 2975
rect 36544 2932 36596 2941
rect 36912 2932 36964 2984
rect 38936 2975 38988 2984
rect 38936 2941 38945 2975
rect 38945 2941 38979 2975
rect 38979 2941 38988 2975
rect 38936 2932 38988 2941
rect 38660 2864 38712 2916
rect 38844 2864 38896 2916
rect 39304 3000 39356 3052
rect 40132 3000 40184 3052
rect 41512 3000 41564 3052
rect 42984 3000 43036 3052
rect 43260 3043 43312 3052
rect 43260 3009 43269 3043
rect 43269 3009 43303 3043
rect 43303 3009 43312 3043
rect 43260 3000 43312 3009
rect 43628 3043 43680 3052
rect 43628 3009 43637 3043
rect 43637 3009 43671 3043
rect 43671 3009 43680 3043
rect 43628 3000 43680 3009
rect 43812 3000 43864 3052
rect 45008 3043 45060 3052
rect 45008 3009 45017 3043
rect 45017 3009 45051 3043
rect 45051 3009 45060 3043
rect 45008 3000 45060 3009
rect 46204 3000 46256 3052
rect 47032 3000 47084 3052
rect 48412 3000 48464 3052
rect 48964 3000 49016 3052
rect 40776 2932 40828 2984
rect 41236 2864 41288 2916
rect 43444 2932 43496 2984
rect 43904 2932 43956 2984
rect 45284 2932 45336 2984
rect 50988 3000 51040 3052
rect 51448 3000 51500 3052
rect 53932 3000 53984 3052
rect 54208 3000 54260 3052
rect 55312 3000 55364 3052
rect 58256 3000 58308 3052
rect 52092 2932 52144 2984
rect 26608 2796 26660 2848
rect 27528 2796 27580 2848
rect 29092 2796 29144 2848
rect 37464 2796 37516 2848
rect 40040 2796 40092 2848
rect 43076 2796 43128 2848
rect 49700 2796 49752 2848
rect 50160 2796 50212 2848
rect 50988 2796 51040 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 7196 2592 7248 2644
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 7840 2524 7892 2576
rect 8392 2524 8444 2576
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 7840 2388 7892 2440
rect 10140 2388 10192 2440
rect 13636 2592 13688 2644
rect 17408 2592 17460 2644
rect 17960 2592 18012 2644
rect 19064 2592 19116 2644
rect 19984 2635 20036 2644
rect 19984 2601 19993 2635
rect 19993 2601 20027 2635
rect 20027 2601 20036 2635
rect 19984 2592 20036 2601
rect 25780 2592 25832 2644
rect 25964 2592 26016 2644
rect 11060 2524 11112 2576
rect 14648 2524 14700 2576
rect 15016 2456 15068 2508
rect 17776 2456 17828 2508
rect 940 2320 992 2372
rect 3240 2363 3292 2372
rect 3240 2329 3249 2363
rect 3249 2329 3283 2363
rect 3283 2329 3292 2363
rect 3240 2320 3292 2329
rect 5356 2252 5408 2304
rect 5816 2363 5868 2372
rect 5816 2329 5825 2363
rect 5825 2329 5859 2363
rect 5859 2329 5868 2363
rect 5816 2320 5868 2329
rect 6920 2363 6972 2372
rect 6920 2329 6929 2363
rect 6929 2329 6963 2363
rect 6963 2329 6972 2363
rect 6920 2320 6972 2329
rect 7104 2363 7156 2372
rect 7104 2329 7113 2363
rect 7113 2329 7147 2363
rect 7147 2329 7156 2363
rect 7104 2320 7156 2329
rect 7656 2363 7708 2372
rect 7656 2329 7665 2363
rect 7665 2329 7699 2363
rect 7699 2329 7708 2363
rect 7656 2320 7708 2329
rect 11244 2388 11296 2440
rect 12348 2431 12400 2440
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 12992 2388 13044 2440
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 15476 2388 15528 2440
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 21364 2524 21416 2576
rect 20444 2499 20496 2508
rect 20444 2465 20453 2499
rect 20453 2465 20487 2499
rect 20487 2465 20496 2499
rect 20444 2456 20496 2465
rect 21180 2456 21232 2508
rect 6828 2252 6880 2304
rect 7748 2295 7800 2304
rect 7748 2261 7757 2295
rect 7757 2261 7791 2295
rect 7791 2261 7800 2295
rect 7748 2252 7800 2261
rect 13452 2320 13504 2372
rect 11060 2252 11112 2304
rect 15844 2252 15896 2304
rect 18236 2320 18288 2372
rect 20260 2388 20312 2440
rect 20536 2388 20588 2440
rect 22100 2388 22152 2440
rect 27436 2456 27488 2508
rect 23480 2388 23532 2440
rect 23664 2388 23716 2440
rect 28172 2456 28224 2508
rect 28908 2524 28960 2576
rect 30288 2524 30340 2576
rect 30472 2592 30524 2644
rect 32128 2524 32180 2576
rect 20720 2320 20772 2372
rect 23204 2320 23256 2372
rect 24768 2320 24820 2372
rect 25504 2363 25556 2372
rect 25504 2329 25513 2363
rect 25513 2329 25547 2363
rect 25547 2329 25556 2363
rect 25504 2320 25556 2329
rect 26424 2363 26476 2372
rect 26424 2329 26433 2363
rect 26433 2329 26467 2363
rect 26467 2329 26476 2363
rect 26424 2320 26476 2329
rect 27620 2320 27672 2372
rect 28356 2388 28408 2440
rect 30012 2388 30064 2440
rect 18880 2252 18932 2304
rect 19064 2252 19116 2304
rect 27528 2252 27580 2304
rect 28908 2320 28960 2372
rect 29920 2320 29972 2372
rect 29828 2252 29880 2304
rect 31116 2431 31168 2440
rect 31116 2397 31125 2431
rect 31125 2397 31159 2431
rect 31159 2397 31168 2431
rect 31116 2388 31168 2397
rect 32496 2388 32548 2440
rect 34888 2431 34940 2440
rect 34888 2397 34897 2431
rect 34897 2397 34931 2431
rect 34931 2397 34940 2431
rect 34888 2388 34940 2397
rect 39488 2524 39540 2576
rect 38660 2456 38712 2508
rect 30472 2363 30524 2372
rect 30472 2329 30481 2363
rect 30481 2329 30515 2363
rect 30515 2329 30524 2363
rect 30472 2320 30524 2329
rect 31024 2320 31076 2372
rect 32588 2363 32640 2372
rect 32588 2329 32597 2363
rect 32597 2329 32631 2363
rect 32631 2329 32640 2363
rect 32588 2320 32640 2329
rect 33508 2363 33560 2372
rect 33508 2329 33517 2363
rect 33517 2329 33551 2363
rect 33551 2329 33560 2363
rect 33508 2320 33560 2329
rect 35164 2363 35216 2372
rect 35164 2329 35173 2363
rect 35173 2329 35207 2363
rect 35207 2329 35216 2363
rect 35164 2320 35216 2329
rect 36084 2363 36136 2372
rect 36084 2329 36093 2363
rect 36093 2329 36127 2363
rect 36127 2329 36136 2363
rect 36084 2320 36136 2329
rect 37740 2363 37792 2372
rect 37740 2329 37749 2363
rect 37749 2329 37783 2363
rect 37783 2329 37792 2363
rect 37740 2320 37792 2329
rect 32220 2252 32272 2304
rect 35440 2252 35492 2304
rect 39120 2388 39172 2440
rect 38660 2363 38712 2372
rect 38660 2329 38669 2363
rect 38669 2329 38703 2363
rect 38703 2329 38712 2363
rect 38660 2320 38712 2329
rect 38844 2320 38896 2372
rect 41052 2363 41104 2372
rect 41052 2329 41061 2363
rect 41061 2329 41095 2363
rect 41095 2329 41104 2363
rect 41052 2320 41104 2329
rect 44088 2592 44140 2644
rect 44180 2592 44232 2644
rect 45836 2592 45888 2644
rect 47400 2592 47452 2644
rect 48872 2635 48924 2644
rect 48872 2601 48881 2635
rect 48881 2601 48915 2635
rect 48915 2601 48924 2635
rect 48872 2592 48924 2601
rect 49700 2592 49752 2644
rect 58256 2635 58308 2644
rect 58256 2601 58265 2635
rect 58265 2601 58299 2635
rect 58299 2601 58308 2635
rect 58256 2592 58308 2601
rect 51080 2524 51132 2576
rect 53472 2524 53524 2576
rect 43352 2388 43404 2440
rect 51816 2456 51868 2508
rect 55680 2499 55732 2508
rect 55680 2465 55689 2499
rect 55689 2465 55723 2499
rect 55723 2465 55732 2499
rect 55680 2456 55732 2465
rect 43904 2431 43956 2440
rect 43904 2397 43913 2431
rect 43913 2397 43947 2431
rect 43947 2397 43956 2431
rect 43904 2388 43956 2397
rect 44088 2388 44140 2440
rect 53840 2431 53892 2440
rect 53840 2397 53849 2431
rect 53849 2397 53883 2431
rect 53883 2397 53892 2431
rect 53840 2388 53892 2397
rect 55220 2388 55272 2440
rect 57244 2388 57296 2440
rect 58992 2388 59044 2440
rect 45192 2320 45244 2372
rect 45284 2363 45336 2372
rect 45284 2329 45293 2363
rect 45293 2329 45327 2363
rect 45327 2329 45336 2363
rect 45284 2320 45336 2329
rect 45928 2320 45980 2372
rect 46296 2320 46348 2372
rect 47400 2320 47452 2372
rect 48780 2363 48832 2372
rect 48780 2329 48789 2363
rect 48789 2329 48823 2363
rect 48823 2329 48832 2363
rect 48780 2320 48832 2329
rect 49700 2320 49752 2372
rect 51080 2320 51132 2372
rect 51908 2363 51960 2372
rect 51908 2329 51917 2363
rect 51917 2329 51951 2363
rect 51951 2329 51960 2363
rect 51908 2320 51960 2329
rect 52552 2320 52604 2372
rect 58900 2320 58952 2372
rect 43536 2252 43588 2304
rect 47216 2252 47268 2304
rect 52460 2252 52512 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 7656 2048 7708 2100
rect 11152 2048 11204 2100
rect 12348 2048 12400 2100
rect 15660 2048 15712 2100
rect 18236 2048 18288 2100
rect 21640 2048 21692 2100
rect 23480 2048 23532 2100
rect 40960 2048 41012 2100
rect 42432 2048 42484 2100
rect 44088 2048 44140 2100
rect 7748 1980 7800 2032
rect 12716 1980 12768 2032
rect 14372 1980 14424 2032
rect 23664 1980 23716 2032
rect 26976 1980 27028 2032
rect 34888 1980 34940 2032
rect 42708 1980 42760 2032
rect 47216 1980 47268 2032
rect 6920 1912 6972 1964
rect 10600 1912 10652 1964
rect 17500 1912 17552 1964
rect 23020 1912 23072 1964
rect 9128 1844 9180 1896
rect 27620 1844 27672 1896
rect 1584 1776 1636 1828
rect 26792 1776 26844 1828
rect 7104 1708 7156 1760
rect 12808 1708 12860 1760
rect 5356 1640 5408 1692
rect 9404 1640 9456 1692
rect 10140 1640 10192 1692
rect 11428 1640 11480 1692
rect 5816 1572 5868 1624
rect 10048 1572 10100 1624
rect 14924 1300 14976 1352
rect 37556 1300 37608 1352
rect 38752 1300 38804 1352
rect 56508 1300 56560 1352
rect 39856 1232 39908 1284
rect 43812 1232 43864 1284
rect 18144 1164 18196 1216
rect 21364 1164 21416 1216
rect 32404 1164 32456 1216
rect 36084 1164 36136 1216
rect 38752 1164 38804 1216
rect 39212 1164 39264 1216
rect 40960 1164 41012 1216
rect 45008 1164 45060 1216
rect 13452 1096 13504 1148
rect 14464 1096 14516 1148
rect 17592 1096 17644 1148
rect 20536 1096 20588 1148
rect 27804 1096 27856 1148
rect 29092 1096 29144 1148
rect 33784 1096 33836 1148
rect 36544 1096 36596 1148
rect 43444 1096 43496 1148
rect 46112 1096 46164 1148
rect 12624 1028 12676 1080
rect 14188 1028 14240 1080
rect 18972 1028 19024 1080
rect 21916 1028 21968 1080
rect 27344 1028 27396 1080
rect 28540 1028 28592 1080
rect 32128 1028 32180 1080
rect 35164 1028 35216 1080
rect 42616 1028 42668 1080
rect 44732 1028 44784 1080
rect 5080 960 5132 1012
rect 6736 960 6788 1012
rect 11060 960 11112 1012
rect 12808 960 12860 1012
rect 14280 960 14332 1012
rect 15568 960 15620 1012
rect 16304 960 16356 1012
rect 3240 892 3292 944
rect 4528 892 4580 944
rect 5172 892 5224 944
rect 6184 892 6236 944
rect 6920 892 6972 944
rect 9496 892 9548 944
rect 13728 892 13780 944
rect 14740 892 14792 944
rect 17316 892 17368 944
rect 18328 892 18380 944
rect 19248 960 19300 1012
rect 20812 960 20864 1012
rect 22008 960 22060 1012
rect 23020 960 23072 1012
rect 23204 960 23256 1012
rect 24400 960 24452 1012
rect 26424 960 26476 1012
rect 28816 960 28868 1012
rect 31852 960 31904 1012
rect 33508 960 33560 1012
rect 19432 892 19484 944
rect 20720 892 20772 944
rect 22192 892 22244 944
rect 23388 892 23440 944
rect 24124 892 24176 944
rect 27528 892 27580 944
rect 28264 892 28316 944
rect 28908 892 28960 944
rect 29368 892 29420 944
rect 31300 892 31352 944
rect 32588 892 32640 944
rect 32956 892 33008 944
rect 35624 960 35676 1012
rect 40684 960 40736 1012
rect 45284 960 45336 1012
rect 47308 960 47360 1012
rect 48780 960 48832 1012
rect 50068 960 50120 1012
rect 51908 960 51960 1012
rect 34060 892 34112 944
rect 37740 892 37792 944
rect 39580 892 39632 944
rect 41052 892 41104 944
rect 42340 892 42392 944
rect 46296 892 46348 944
rect 46480 892 46532 944
rect 47400 892 47452 944
rect 49240 892 49292 944
rect 51080 892 51132 944
rect 47952 824 48004 876
rect 49700 824 49752 876
rect 35256 348 35308 400
rect 38936 348 38988 400
rect 34980 144 35032 196
rect 38660 144 38712 196
rect 35532 76 35584 128
rect 38844 76 38896 128
<< metal2 >>
rect 846 63200 902 64000
rect 1582 63200 1638 64000
rect 2318 63322 2374 64000
rect 3054 63322 3110 64000
rect 3790 63322 3846 64000
rect 4526 63322 4582 64000
rect 5262 63322 5318 64000
rect 5998 63322 6054 64000
rect 6734 63322 6790 64000
rect 2318 63294 2636 63322
rect 2318 63200 2374 63294
rect 860 59022 888 63200
rect 938 61840 994 61849
rect 938 61775 994 61784
rect 952 61198 980 61775
rect 940 61192 992 61198
rect 940 61134 992 61140
rect 1030 61160 1086 61169
rect 1030 61095 1032 61104
rect 1084 61095 1086 61104
rect 1032 61066 1084 61072
rect 940 60716 992 60722
rect 940 60658 992 60664
rect 952 60489 980 60658
rect 938 60480 994 60489
rect 938 60415 994 60424
rect 940 60036 992 60042
rect 940 59978 992 59984
rect 952 59809 980 59978
rect 938 59800 994 59809
rect 938 59735 994 59744
rect 1596 59702 1624 63200
rect 2608 60110 2636 63294
rect 3054 63294 3280 63322
rect 3054 63200 3110 63294
rect 3252 60790 3280 63294
rect 3790 63294 4016 63322
rect 3790 63200 3846 63294
rect 3988 60790 4016 63294
rect 4526 63294 4660 63322
rect 4526 63200 4582 63294
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 4632 61198 4660 63294
rect 5092 63294 5318 63322
rect 5092 61198 5120 63294
rect 5262 63200 5318 63294
rect 5736 63294 6054 63322
rect 5172 61600 5224 61606
rect 5172 61542 5224 61548
rect 5184 61402 5212 61542
rect 5172 61396 5224 61402
rect 5172 61338 5224 61344
rect 5736 61198 5764 63294
rect 5998 63200 6054 63294
rect 6656 63294 6790 63322
rect 6656 61198 6684 63294
rect 6734 63200 6790 63294
rect 7470 63322 7526 64000
rect 8206 63322 8262 64000
rect 8942 63322 8998 64000
rect 7470 63294 7604 63322
rect 7470 63200 7526 63294
rect 7576 61198 7604 63294
rect 8206 63294 8432 63322
rect 8206 63200 8262 63294
rect 8208 61396 8260 61402
rect 8208 61338 8260 61344
rect 7656 61260 7708 61266
rect 7656 61202 7708 61208
rect 4620 61192 4672 61198
rect 4620 61134 4672 61140
rect 5080 61192 5132 61198
rect 5080 61134 5132 61140
rect 5724 61192 5776 61198
rect 5724 61134 5776 61140
rect 6644 61192 6696 61198
rect 6644 61134 6696 61140
rect 7564 61192 7616 61198
rect 7564 61134 7616 61140
rect 5632 61124 5684 61130
rect 5632 61066 5684 61072
rect 6184 61124 6236 61130
rect 6184 61066 6236 61072
rect 6920 61124 6972 61130
rect 6920 61066 6972 61072
rect 3240 60784 3292 60790
rect 3240 60726 3292 60732
rect 3976 60784 4028 60790
rect 3976 60726 4028 60732
rect 4620 60580 4672 60586
rect 4620 60522 4672 60528
rect 3332 60512 3384 60518
rect 3332 60454 3384 60460
rect 3344 60314 3372 60454
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 3332 60308 3384 60314
rect 3332 60250 3384 60256
rect 2596 60104 2648 60110
rect 2596 60046 2648 60052
rect 2044 60036 2096 60042
rect 2044 59978 2096 59984
rect 1584 59696 1636 59702
rect 1584 59638 1636 59644
rect 940 59628 992 59634
rect 940 59570 992 59576
rect 952 59129 980 59570
rect 1952 59424 2004 59430
rect 1952 59366 2004 59372
rect 938 59120 994 59129
rect 1964 59090 1992 59366
rect 938 59055 994 59064
rect 1952 59084 2004 59090
rect 1952 59026 2004 59032
rect 848 59016 900 59022
rect 848 58958 900 58964
rect 2056 58682 2084 59978
rect 2504 59968 2556 59974
rect 2504 59910 2556 59916
rect 2320 59424 2372 59430
rect 2320 59366 2372 59372
rect 2044 58676 2096 58682
rect 2044 58618 2096 58624
rect 940 58540 992 58546
rect 940 58482 992 58488
rect 952 58449 980 58482
rect 938 58440 994 58449
rect 938 58375 994 58384
rect 940 57928 992 57934
rect 940 57870 992 57876
rect 952 57769 980 57870
rect 938 57760 994 57769
rect 938 57695 994 57704
rect 940 57452 992 57458
rect 940 57394 992 57400
rect 952 57089 980 57394
rect 1768 57248 1820 57254
rect 1768 57190 1820 57196
rect 938 57080 994 57089
rect 938 57015 994 57024
rect 940 56772 992 56778
rect 940 56714 992 56720
rect 952 56409 980 56714
rect 938 56400 994 56409
rect 938 56335 994 56344
rect 1780 55894 1808 57190
rect 1768 55888 1820 55894
rect 1768 55830 1820 55836
rect 938 55720 994 55729
rect 938 55655 940 55664
rect 992 55655 994 55664
rect 940 55626 992 55632
rect 940 55276 992 55282
rect 940 55218 992 55224
rect 952 55049 980 55218
rect 938 55040 994 55049
rect 938 54975 994 54984
rect 940 54596 992 54602
rect 940 54538 992 54544
rect 952 54369 980 54538
rect 938 54360 994 54369
rect 938 54295 994 54304
rect 940 54188 992 54194
rect 940 54130 992 54136
rect 952 53689 980 54130
rect 1768 53984 1820 53990
rect 1768 53926 1820 53932
rect 938 53680 994 53689
rect 938 53615 994 53624
rect 1780 53446 1808 53926
rect 1768 53440 1820 53446
rect 1768 53382 1820 53388
rect 940 53100 992 53106
rect 940 53042 992 53048
rect 952 53009 980 53042
rect 938 53000 994 53009
rect 938 52935 994 52944
rect 2042 52592 2098 52601
rect 2042 52527 2098 52536
rect 2056 52494 2084 52527
rect 2044 52488 2096 52494
rect 2044 52430 2096 52436
rect 940 52420 992 52426
rect 940 52362 992 52368
rect 952 52329 980 52362
rect 938 52320 994 52329
rect 938 52255 994 52264
rect 940 52012 992 52018
rect 940 51954 992 51960
rect 952 51649 980 51954
rect 938 51640 994 51649
rect 938 51575 994 51584
rect 940 51332 992 51338
rect 940 51274 992 51280
rect 952 50969 980 51274
rect 938 50960 994 50969
rect 938 50895 994 50904
rect 938 50280 994 50289
rect 938 50215 940 50224
rect 992 50215 994 50224
rect 2044 50244 2096 50250
rect 940 50186 992 50192
rect 2044 50186 2096 50192
rect 940 49836 992 49842
rect 940 49778 992 49784
rect 952 49609 980 49778
rect 938 49600 994 49609
rect 938 49535 994 49544
rect 940 49224 992 49230
rect 940 49166 992 49172
rect 952 48929 980 49166
rect 938 48920 994 48929
rect 938 48855 994 48864
rect 940 48748 992 48754
rect 940 48690 992 48696
rect 952 48249 980 48690
rect 1952 48612 2004 48618
rect 1952 48554 2004 48560
rect 938 48240 994 48249
rect 938 48175 994 48184
rect 1584 48000 1636 48006
rect 1584 47942 1636 47948
rect 940 47660 992 47666
rect 940 47602 992 47608
rect 952 47569 980 47602
rect 938 47560 994 47569
rect 938 47495 994 47504
rect 940 47048 992 47054
rect 940 46990 992 46996
rect 952 46889 980 46990
rect 938 46880 994 46889
rect 938 46815 994 46824
rect 940 46572 992 46578
rect 940 46514 992 46520
rect 952 46209 980 46514
rect 938 46200 994 46209
rect 938 46135 994 46144
rect 940 45892 992 45898
rect 940 45834 992 45840
rect 952 45529 980 45834
rect 938 45520 994 45529
rect 938 45455 994 45464
rect 940 44872 992 44878
rect 938 44840 940 44849
rect 992 44840 994 44849
rect 938 44775 994 44784
rect 940 44396 992 44402
rect 940 44338 992 44344
rect 952 44169 980 44338
rect 938 44160 994 44169
rect 938 44095 994 44104
rect 940 43716 992 43722
rect 940 43658 992 43664
rect 952 43489 980 43658
rect 938 43480 994 43489
rect 938 43415 994 43424
rect 940 43308 992 43314
rect 940 43250 992 43256
rect 952 42809 980 43250
rect 938 42800 994 42809
rect 938 42735 994 42744
rect 940 42220 992 42226
rect 940 42162 992 42168
rect 952 42129 980 42162
rect 938 42120 994 42129
rect 938 42055 994 42064
rect 940 41540 992 41546
rect 940 41482 992 41488
rect 952 41449 980 41482
rect 938 41440 994 41449
rect 938 41375 994 41384
rect 940 41132 992 41138
rect 940 41074 992 41080
rect 952 40769 980 41074
rect 938 40760 994 40769
rect 938 40695 994 40704
rect 940 40452 992 40458
rect 940 40394 992 40400
rect 952 40089 980 40394
rect 1032 40112 1084 40118
rect 938 40080 994 40089
rect 1032 40054 1084 40060
rect 938 40015 994 40024
rect 1044 39409 1072 40054
rect 1030 39400 1086 39409
rect 940 39364 992 39370
rect 1030 39335 1086 39344
rect 940 39306 992 39312
rect 952 38729 980 39306
rect 1032 38956 1084 38962
rect 1032 38898 1084 38904
rect 938 38720 994 38729
rect 938 38655 994 38664
rect 1044 38049 1072 38898
rect 1030 38040 1086 38049
rect 1030 37975 1086 37984
rect 940 37868 992 37874
rect 940 37810 992 37816
rect 952 37369 980 37810
rect 938 37360 994 37369
rect 938 37295 994 37304
rect 940 36780 992 36786
rect 940 36722 992 36728
rect 952 36689 980 36722
rect 938 36680 994 36689
rect 938 36615 994 36624
rect 940 36100 992 36106
rect 940 36042 992 36048
rect 952 36009 980 36042
rect 938 36000 994 36009
rect 938 35935 994 35944
rect 1596 35834 1624 47942
rect 1768 47456 1820 47462
rect 1768 47398 1820 47404
rect 1780 43194 1808 47398
rect 1860 44872 1912 44878
rect 1858 44840 1860 44849
rect 1912 44840 1914 44849
rect 1858 44775 1914 44784
rect 1780 43166 1900 43194
rect 1768 43104 1820 43110
rect 1768 43046 1820 43052
rect 1780 42226 1808 43046
rect 1768 42220 1820 42226
rect 1768 42162 1820 42168
rect 1872 38486 1900 43166
rect 1860 38480 1912 38486
rect 1860 38422 1912 38428
rect 1676 38412 1728 38418
rect 1676 38354 1728 38360
rect 1584 35828 1636 35834
rect 1584 35770 1636 35776
rect 940 35692 992 35698
rect 940 35634 992 35640
rect 952 35329 980 35634
rect 938 35320 994 35329
rect 938 35255 994 35264
rect 940 35012 992 35018
rect 940 34954 992 34960
rect 952 34649 980 34954
rect 938 34640 994 34649
rect 938 34575 994 34584
rect 940 33992 992 33998
rect 938 33960 940 33969
rect 992 33960 994 33969
rect 938 33895 994 33904
rect 940 33516 992 33522
rect 940 33458 992 33464
rect 952 33289 980 33458
rect 938 33280 994 33289
rect 938 33215 994 33224
rect 940 32836 992 32842
rect 940 32778 992 32784
rect 952 32609 980 32778
rect 938 32600 994 32609
rect 938 32535 994 32544
rect 940 32428 992 32434
rect 940 32370 992 32376
rect 952 31929 980 32370
rect 938 31920 994 31929
rect 938 31855 994 31864
rect 940 31340 992 31346
rect 940 31282 992 31288
rect 952 31249 980 31282
rect 938 31240 994 31249
rect 938 31175 994 31184
rect 940 30660 992 30666
rect 940 30602 992 30608
rect 952 30569 980 30602
rect 938 30560 994 30569
rect 938 30495 994 30504
rect 940 30184 992 30190
rect 940 30126 992 30132
rect 952 29889 980 30126
rect 938 29880 994 29889
rect 938 29815 994 29824
rect 940 29572 992 29578
rect 940 29514 992 29520
rect 952 29209 980 29514
rect 938 29200 994 29209
rect 938 29135 994 29144
rect 1688 28694 1716 38354
rect 1964 38350 1992 48554
rect 2056 48142 2084 50186
rect 2044 48136 2096 48142
rect 2044 48078 2096 48084
rect 2136 42016 2188 42022
rect 2136 41958 2188 41964
rect 1952 38344 2004 38350
rect 1952 38286 2004 38292
rect 1860 37732 1912 37738
rect 1860 37674 1912 37680
rect 1872 32434 1900 37674
rect 1860 32428 1912 32434
rect 1860 32370 1912 32376
rect 1952 29640 2004 29646
rect 1952 29582 2004 29588
rect 1676 28688 1728 28694
rect 1676 28630 1728 28636
rect 940 28620 992 28626
rect 940 28562 992 28568
rect 952 28529 980 28562
rect 938 28520 994 28529
rect 938 28455 994 28464
rect 940 28008 992 28014
rect 940 27950 992 27956
rect 952 27849 980 27950
rect 938 27840 994 27849
rect 938 27775 994 27784
rect 1584 27464 1636 27470
rect 1584 27406 1636 27412
rect 940 27396 992 27402
rect 940 27338 992 27344
rect 952 27169 980 27338
rect 938 27160 994 27169
rect 1596 27130 1624 27406
rect 938 27095 994 27104
rect 1584 27124 1636 27130
rect 1584 27066 1636 27072
rect 1676 26988 1728 26994
rect 1676 26930 1728 26936
rect 940 26920 992 26926
rect 940 26862 992 26868
rect 952 26489 980 26862
rect 938 26480 994 26489
rect 938 26415 994 26424
rect 940 25832 992 25838
rect 938 25800 940 25809
rect 992 25800 994 25809
rect 938 25735 994 25744
rect 940 25220 992 25226
rect 940 25162 992 25168
rect 952 25129 980 25162
rect 938 25120 994 25129
rect 938 25055 994 25064
rect 940 24744 992 24750
rect 940 24686 992 24692
rect 952 24449 980 24686
rect 938 24440 994 24449
rect 938 24375 994 24384
rect 940 24132 992 24138
rect 940 24074 992 24080
rect 952 23769 980 24074
rect 938 23760 994 23769
rect 938 23695 994 23704
rect 940 23180 992 23186
rect 940 23122 992 23128
rect 952 23089 980 23122
rect 938 23080 994 23089
rect 938 23015 994 23024
rect 940 22568 992 22574
rect 940 22510 992 22516
rect 952 22409 980 22510
rect 938 22400 994 22409
rect 938 22335 994 22344
rect 940 21956 992 21962
rect 940 21898 992 21904
rect 952 21729 980 21898
rect 938 21720 994 21729
rect 938 21655 994 21664
rect 940 21344 992 21350
rect 940 21286 992 21292
rect 952 21049 980 21286
rect 938 21040 994 21049
rect 938 20975 994 20984
rect 940 20392 992 20398
rect 938 20360 940 20369
rect 992 20360 994 20369
rect 938 20295 994 20304
rect 940 19780 992 19786
rect 940 19722 992 19728
rect 952 19689 980 19722
rect 938 19680 994 19689
rect 938 19615 994 19624
rect 940 19440 992 19446
rect 940 19382 992 19388
rect 952 19009 980 19382
rect 938 19000 994 19009
rect 938 18935 994 18944
rect 940 18692 992 18698
rect 940 18634 992 18640
rect 952 18329 980 18634
rect 938 18320 994 18329
rect 938 18255 994 18264
rect 940 17740 992 17746
rect 940 17682 992 17688
rect 952 17649 980 17682
rect 938 17640 994 17649
rect 938 17575 994 17584
rect 940 17128 992 17134
rect 940 17070 992 17076
rect 952 16969 980 17070
rect 938 16960 994 16969
rect 938 16895 994 16904
rect 940 16516 992 16522
rect 940 16458 992 16464
rect 952 16289 980 16458
rect 938 16280 994 16289
rect 938 16215 994 16224
rect 940 16040 992 16046
rect 940 15982 992 15988
rect 952 15609 980 15982
rect 938 15600 994 15609
rect 938 15535 994 15544
rect 940 14952 992 14958
rect 938 14920 940 14929
rect 992 14920 994 14929
rect 938 14855 994 14864
rect 1582 14512 1638 14521
rect 1582 14447 1638 14456
rect 1596 14414 1624 14447
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 940 14340 992 14346
rect 940 14282 992 14288
rect 952 14249 980 14282
rect 938 14240 994 14249
rect 938 14175 994 14184
rect 940 13864 992 13870
rect 940 13806 992 13812
rect 952 13569 980 13806
rect 938 13560 994 13569
rect 938 13495 994 13504
rect 1582 13424 1638 13433
rect 1582 13359 1638 13368
rect 1596 13326 1624 13359
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 940 13252 992 13258
rect 940 13194 992 13200
rect 952 12889 980 13194
rect 938 12880 994 12889
rect 938 12815 994 12824
rect 938 12200 994 12209
rect 938 12135 994 12144
rect 952 11830 980 12135
rect 940 11824 992 11830
rect 940 11766 992 11772
rect 938 11520 994 11529
rect 938 11455 994 11464
rect 952 11218 980 11455
rect 940 11212 992 11218
rect 940 11154 992 11160
rect 938 10840 994 10849
rect 938 10775 994 10784
rect 952 10742 980 10775
rect 940 10736 992 10742
rect 940 10678 992 10684
rect 1688 10606 1716 26930
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 938 10160 994 10169
rect 938 10095 940 10104
rect 992 10095 994 10104
rect 940 10066 992 10072
rect 940 9512 992 9518
rect 938 9480 940 9489
rect 992 9480 994 9489
rect 938 9415 994 9424
rect 940 8900 992 8906
rect 940 8842 992 8848
rect 952 8809 980 8842
rect 938 8800 994 8809
rect 938 8735 994 8744
rect 940 8424 992 8430
rect 940 8366 992 8372
rect 952 8129 980 8366
rect 938 8120 994 8129
rect 938 8055 994 8064
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 940 7812 992 7818
rect 940 7754 992 7760
rect 952 7449 980 7754
rect 938 7440 994 7449
rect 1596 7410 1624 7822
rect 938 7375 994 7384
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 940 6860 992 6866
rect 940 6802 992 6808
rect 952 6769 980 6802
rect 1872 6769 1900 16050
rect 1964 9926 1992 29582
rect 2148 26926 2176 41958
rect 2228 39500 2280 39506
rect 2228 39442 2280 39448
rect 2240 36106 2268 39442
rect 2332 39438 2360 59366
rect 2412 48136 2464 48142
rect 2412 48078 2464 48084
rect 2320 39432 2372 39438
rect 2320 39374 2372 39380
rect 2424 38350 2452 48078
rect 2412 38344 2464 38350
rect 2412 38286 2464 38292
rect 2320 38276 2372 38282
rect 2320 38218 2372 38224
rect 2228 36100 2280 36106
rect 2228 36042 2280 36048
rect 2332 33590 2360 38218
rect 2424 37194 2452 38286
rect 2412 37188 2464 37194
rect 2412 37130 2464 37136
rect 2424 36242 2452 37130
rect 2412 36236 2464 36242
rect 2412 36178 2464 36184
rect 2320 33584 2372 33590
rect 2320 33526 2372 33532
rect 2320 28076 2372 28082
rect 2320 28018 2372 28024
rect 2136 26920 2188 26926
rect 2136 26862 2188 26868
rect 2332 12374 2360 28018
rect 2424 27062 2452 36178
rect 2516 36174 2544 59910
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 3424 58472 3476 58478
rect 3424 58414 3476 58420
rect 2688 50992 2740 50998
rect 2688 50934 2740 50940
rect 2596 39840 2648 39846
rect 2596 39782 2648 39788
rect 2608 39438 2636 39782
rect 2700 39574 2728 50934
rect 3436 47598 3464 58414
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 3976 51332 4028 51338
rect 3976 51274 4028 51280
rect 3988 50998 4016 51274
rect 3976 50992 4028 50998
rect 3976 50934 4028 50940
rect 4068 50924 4120 50930
rect 4068 50866 4120 50872
rect 4080 49842 4108 50866
rect 4632 50862 4660 60522
rect 5644 60110 5672 61066
rect 5908 61056 5960 61062
rect 5908 60998 5960 61004
rect 5632 60104 5684 60110
rect 5632 60046 5684 60052
rect 4620 50856 4672 50862
rect 4620 50798 4672 50804
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4068 49836 4120 49842
rect 4068 49778 4120 49784
rect 4080 48210 4108 49778
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4068 48204 4120 48210
rect 4068 48146 4120 48152
rect 3424 47592 3476 47598
rect 3424 47534 3476 47540
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 2688 39568 2740 39574
rect 2688 39510 2740 39516
rect 2596 39432 2648 39438
rect 2596 39374 2648 39380
rect 2688 39432 2740 39438
rect 2688 39374 2740 39380
rect 2700 38350 2728 39374
rect 3056 39296 3108 39302
rect 3056 39238 3108 39244
rect 3068 38418 3096 39238
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 3056 38412 3108 38418
rect 3056 38354 3108 38360
rect 2688 38344 2740 38350
rect 2688 38286 2740 38292
rect 2596 38208 2648 38214
rect 2596 38150 2648 38156
rect 2608 38010 2636 38150
rect 2596 38004 2648 38010
rect 2596 37946 2648 37952
rect 5920 37942 5948 60998
rect 6000 57860 6052 57866
rect 6000 57802 6052 57808
rect 6012 50386 6040 57802
rect 6000 50380 6052 50386
rect 6000 50322 6052 50328
rect 5908 37936 5960 37942
rect 5908 37878 5960 37884
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 6000 37256 6052 37262
rect 6000 37198 6052 37204
rect 5540 37120 5592 37126
rect 5540 37062 5592 37068
rect 3424 36576 3476 36582
rect 3424 36518 3476 36524
rect 2504 36168 2556 36174
rect 2504 36110 2556 36116
rect 2780 36100 2832 36106
rect 2780 36042 2832 36048
rect 2792 35222 2820 36042
rect 2780 35216 2832 35222
rect 2780 35158 2832 35164
rect 2596 28688 2648 28694
rect 2596 28630 2648 28636
rect 2608 28558 2636 28630
rect 2596 28552 2648 28558
rect 2596 28494 2648 28500
rect 2412 27056 2464 27062
rect 2412 26998 2464 27004
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 2596 26988 2648 26994
rect 2596 26930 2648 26936
rect 2516 25294 2544 26930
rect 2504 25288 2556 25294
rect 2504 25230 2556 25236
rect 2516 24070 2544 25230
rect 2504 24064 2556 24070
rect 2504 24006 2556 24012
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 2424 16998 2452 17138
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2320 12368 2372 12374
rect 2320 12310 2372 12316
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 2424 9489 2452 16934
rect 2608 16574 2636 26930
rect 2688 25288 2740 25294
rect 2688 25230 2740 25236
rect 2700 24342 2728 25230
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 2884 24410 2912 24754
rect 2872 24404 2924 24410
rect 2872 24346 2924 24352
rect 2688 24336 2740 24342
rect 2688 24278 2740 24284
rect 2688 24200 2740 24206
rect 2688 24142 2740 24148
rect 2700 24070 2728 24142
rect 2688 24064 2740 24070
rect 2688 24006 2740 24012
rect 2608 16546 2728 16574
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 2410 9480 2466 9489
rect 2410 9415 2466 9424
rect 2516 8945 2544 13806
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2608 11898 2636 12174
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2502 8936 2558 8945
rect 2502 8871 2558 8880
rect 2700 7818 2728 16546
rect 3436 13802 3464 36518
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3528 10810 3556 20402
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 5276 17882 5304 18702
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5552 17785 5580 37062
rect 6012 36922 6040 37198
rect 6000 36916 6052 36922
rect 6000 36858 6052 36864
rect 6196 35193 6224 61066
rect 6276 50720 6328 50726
rect 6276 50662 6328 50668
rect 6288 37262 6316 50662
rect 6828 49836 6880 49842
rect 6828 49778 6880 49784
rect 6460 49088 6512 49094
rect 6460 49030 6512 49036
rect 6472 42090 6500 49030
rect 6840 48210 6868 49778
rect 6828 48204 6880 48210
rect 6828 48146 6880 48152
rect 6460 42084 6512 42090
rect 6460 42026 6512 42032
rect 6368 41540 6420 41546
rect 6368 41482 6420 41488
rect 6276 37256 6328 37262
rect 6276 37198 6328 37204
rect 6182 35184 6238 35193
rect 6182 35119 6238 35128
rect 6380 29782 6408 41482
rect 6736 37256 6788 37262
rect 6736 37198 6788 37204
rect 6748 36378 6776 37198
rect 6736 36372 6788 36378
rect 6736 36314 6788 36320
rect 6368 29776 6420 29782
rect 6368 29718 6420 29724
rect 6932 22094 6960 61066
rect 7564 60036 7616 60042
rect 7564 59978 7616 59984
rect 7576 59702 7604 59978
rect 7564 59696 7616 59702
rect 7564 59638 7616 59644
rect 7668 55214 7696 61202
rect 7932 60648 7984 60654
rect 7932 60590 7984 60596
rect 7748 60104 7800 60110
rect 7748 60046 7800 60052
rect 7760 59770 7788 60046
rect 7748 59764 7800 59770
rect 7748 59706 7800 59712
rect 7668 55186 7788 55214
rect 7760 44305 7788 55186
rect 7840 51808 7892 51814
rect 7840 51750 7892 51756
rect 7746 44296 7802 44305
rect 7746 44231 7802 44240
rect 7852 26994 7880 51750
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 7944 24274 7972 60590
rect 8220 60042 8248 61338
rect 8404 60790 8432 63294
rect 8942 63294 9076 63322
rect 8942 63200 8998 63294
rect 8392 60784 8444 60790
rect 8392 60726 8444 60732
rect 9048 60722 9076 63294
rect 9678 63200 9734 64000
rect 10414 63322 10470 64000
rect 10244 63294 10470 63322
rect 9692 61198 9720 63200
rect 9772 61668 9824 61674
rect 9772 61610 9824 61616
rect 9784 61334 9812 61610
rect 9772 61328 9824 61334
rect 9772 61270 9824 61276
rect 10244 61198 10272 63294
rect 10414 63200 10470 63294
rect 11150 63200 11206 64000
rect 11886 63322 11942 64000
rect 12622 63322 12678 64000
rect 13358 63322 13414 64000
rect 14094 63322 14150 64000
rect 14830 63322 14886 64000
rect 15566 63322 15622 64000
rect 16302 63322 16358 64000
rect 11886 63294 12020 63322
rect 11886 63200 11942 63294
rect 11164 61198 11192 63200
rect 11992 61198 12020 63294
rect 12622 63294 12756 63322
rect 12622 63200 12678 63294
rect 12728 61198 12756 63294
rect 13358 63294 13584 63322
rect 13358 63200 13414 63294
rect 9680 61192 9732 61198
rect 9680 61134 9732 61140
rect 10232 61192 10284 61198
rect 10232 61134 10284 61140
rect 11152 61192 11204 61198
rect 11152 61134 11204 61140
rect 11980 61192 12032 61198
rect 11980 61134 12032 61140
rect 12716 61192 12768 61198
rect 12716 61134 12768 61140
rect 9128 61124 9180 61130
rect 9128 61066 9180 61072
rect 9036 60716 9088 60722
rect 9036 60658 9088 60664
rect 8208 60036 8260 60042
rect 8208 59978 8260 59984
rect 8024 59968 8076 59974
rect 8024 59910 8076 59916
rect 8036 52018 8064 59910
rect 8024 52012 8076 52018
rect 8024 51954 8076 51960
rect 8300 52012 8352 52018
rect 8300 51954 8352 51960
rect 8312 49842 8340 51954
rect 8300 49836 8352 49842
rect 8300 49778 8352 49784
rect 9036 48204 9088 48210
rect 9036 48146 9088 48152
rect 8944 47184 8996 47190
rect 8944 47126 8996 47132
rect 8956 30054 8984 47126
rect 9048 45354 9076 48146
rect 9140 47666 9168 61066
rect 12164 61056 12216 61062
rect 12164 60998 12216 61004
rect 9220 60512 9272 60518
rect 9220 60454 9272 60460
rect 9128 47660 9180 47666
rect 9128 47602 9180 47608
rect 9036 45348 9088 45354
rect 9036 45290 9088 45296
rect 9232 44810 9260 60454
rect 9220 44804 9272 44810
rect 9220 44746 9272 44752
rect 9588 44260 9640 44266
rect 9588 44202 9640 44208
rect 9600 43790 9628 44202
rect 9588 43784 9640 43790
rect 9588 43726 9640 43732
rect 11704 40384 11756 40390
rect 11704 40326 11756 40332
rect 11716 38418 11744 40326
rect 11704 38412 11756 38418
rect 11704 38354 11756 38360
rect 12176 33590 12204 60998
rect 13556 60790 13584 63294
rect 14094 63294 14320 63322
rect 14094 63200 14150 63294
rect 13636 61124 13688 61130
rect 13636 61066 13688 61072
rect 13544 60784 13596 60790
rect 13544 60726 13596 60732
rect 13084 49768 13136 49774
rect 13084 49710 13136 49716
rect 13096 42158 13124 49710
rect 13084 42152 13136 42158
rect 13084 42094 13136 42100
rect 12164 33584 12216 33590
rect 12164 33526 12216 33532
rect 9772 30252 9824 30258
rect 9772 30194 9824 30200
rect 8944 30048 8996 30054
rect 8944 29990 8996 29996
rect 9784 29306 9812 30194
rect 9772 29300 9824 29306
rect 9772 29242 9824 29248
rect 9404 29164 9456 29170
rect 9404 29106 9456 29112
rect 9416 28626 9444 29106
rect 9404 28620 9456 28626
rect 9404 28562 9456 28568
rect 9416 25906 9444 28562
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 10692 25900 10744 25906
rect 10692 25842 10744 25848
rect 7932 24268 7984 24274
rect 7932 24210 7984 24216
rect 8944 24064 8996 24070
rect 8944 24006 8996 24012
rect 6932 22066 7052 22094
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6840 21690 6868 21966
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 6104 19310 6132 21490
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 6092 19304 6144 19310
rect 6092 19246 6144 19252
rect 6104 18834 6132 19246
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5736 18290 5764 18566
rect 6104 18358 6132 18770
rect 6932 18698 6960 19722
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6092 18352 6144 18358
rect 6092 18294 6144 18300
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 5538 17776 5594 17785
rect 5538 17711 5594 17720
rect 6564 17678 6592 18022
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6472 17270 6500 17614
rect 6748 17542 6776 18634
rect 6932 18222 6960 18634
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6460 17264 6512 17270
rect 6460 17206 6512 17212
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 7024 13297 7052 22066
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 8128 19990 8156 20198
rect 8116 19984 8168 19990
rect 8116 19926 8168 19932
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7116 19378 7144 19654
rect 7576 19514 7604 19790
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 8404 18970 8432 19790
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 7116 18222 7144 18702
rect 8220 18578 8248 18702
rect 8404 18630 8432 18702
rect 8128 18550 8248 18578
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8128 18426 8156 18550
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 8128 17746 8156 18362
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8496 17338 8524 18158
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8588 17202 8616 17478
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8864 14074 8892 14350
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 7010 13288 7066 13297
rect 7010 13223 7066 13232
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 6184 12368 6236 12374
rect 6184 12310 6236 12316
rect 4066 12200 4122 12209
rect 4066 12135 4122 12144
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 4080 9586 4108 12135
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 938 6760 994 6769
rect 938 6695 994 6704
rect 1858 6760 1914 6769
rect 1858 6695 1914 6704
rect 940 6248 992 6254
rect 940 6190 992 6196
rect 952 6089 980 6190
rect 938 6080 994 6089
rect 938 6015 994 6024
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 940 5636 992 5642
rect 940 5578 992 5584
rect 952 5409 980 5578
rect 938 5400 994 5409
rect 938 5335 994 5344
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 952 4729 980 5102
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 5262 4992 5318 5001
rect 4214 4924 4522 4933
rect 5262 4927 5318 4936
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 940 4072 992 4078
rect 938 4040 940 4049
rect 992 4040 994 4049
rect 938 3975 994 3984
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 5276 3670 5304 4927
rect 5908 4548 5960 4554
rect 5908 4490 5960 4496
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5736 4049 5764 4082
rect 5722 4040 5778 4049
rect 5722 3975 5778 3984
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 940 3460 992 3466
rect 940 3402 992 3408
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 952 3369 980 3402
rect 938 3360 994 3369
rect 938 3295 994 3304
rect 940 2984 992 2990
rect 940 2926 992 2932
rect 952 2689 980 2926
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 938 2680 994 2689
rect 4214 2683 4522 2692
rect 938 2615 994 2624
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 940 2372 992 2378
rect 940 2314 992 2320
rect 952 2009 980 2314
rect 938 2000 994 2009
rect 938 1935 994 1944
rect 1596 1834 1624 2382
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 1584 1828 1636 1834
rect 1584 1770 1636 1776
rect 3252 950 3280 2314
rect 5092 1018 5120 3402
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5172 3120 5224 3126
rect 5828 3097 5856 3130
rect 5172 3062 5224 3068
rect 5814 3088 5870 3097
rect 5080 1012 5132 1018
rect 5080 954 5132 960
rect 5184 950 5212 3062
rect 5814 3023 5870 3032
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 5368 1698 5396 2246
rect 5356 1692 5408 1698
rect 5356 1634 5408 1640
rect 5828 1630 5856 2314
rect 5816 1624 5868 1630
rect 5816 1566 5868 1572
rect 3240 944 3292 950
rect 3240 886 3292 892
rect 4528 944 4580 950
rect 4528 886 4580 892
rect 5172 944 5224 950
rect 5172 886 5224 892
rect 4540 800 4568 886
rect 5920 800 5948 4490
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 6012 2961 6040 3946
rect 6104 3194 6132 5034
rect 6196 3670 6224 12310
rect 8956 11082 8984 24006
rect 10704 23118 10732 25842
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 12176 23322 12204 24074
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 12164 23316 12216 23322
rect 12164 23258 12216 23264
rect 12820 23118 12848 23598
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9784 22098 9812 22578
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 10152 21962 10180 23054
rect 10140 21956 10192 21962
rect 10140 21898 10192 21904
rect 10152 21554 10180 21898
rect 10140 21548 10192 21554
rect 10140 21490 10192 21496
rect 9678 20496 9734 20505
rect 9312 20460 9364 20466
rect 9678 20431 9734 20440
rect 9312 20402 9364 20408
rect 9324 20058 9352 20402
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 9692 19514 9720 20431
rect 10152 20210 10180 21490
rect 13268 21344 13320 21350
rect 13268 21286 13320 21292
rect 13176 21140 13228 21146
rect 13176 21082 13228 21088
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 9784 20182 10180 20210
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9048 18958 9352 18986
rect 9048 18902 9076 18958
rect 9324 18902 9352 18958
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9036 18896 9088 18902
rect 9036 18838 9088 18844
rect 9312 18896 9364 18902
rect 9312 18838 9364 18844
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9324 18222 9352 18566
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9600 18086 9628 18906
rect 9692 18290 9720 19110
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9784 17490 9812 20182
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9876 18426 9904 19790
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10060 19378 10088 19654
rect 10152 19514 10180 19994
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 10244 18970 10272 20402
rect 10324 20256 10376 20262
rect 10324 20198 10376 20204
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9968 18358 9996 18566
rect 9956 18352 10008 18358
rect 9956 18294 10008 18300
rect 9968 17746 9996 18294
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 10060 17678 10088 18634
rect 10152 18358 10180 18702
rect 10140 18352 10192 18358
rect 10140 18294 10192 18300
rect 10244 17882 10272 18770
rect 10336 18290 10364 20198
rect 10692 19440 10744 19446
rect 10692 19382 10744 19388
rect 10704 18630 10732 19382
rect 10980 19242 11008 20198
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 11164 19514 11192 19790
rect 11152 19508 11204 19514
rect 11152 19450 11204 19456
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10336 17746 10364 17818
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 9784 17462 9996 17490
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9324 14482 9352 14962
rect 9692 14958 9720 15846
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 13326 9720 14214
rect 9784 13870 9812 15438
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9784 12986 9812 13806
rect 9876 13530 9904 14350
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9968 12306 9996 17462
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10336 15706 10364 16050
rect 10428 15706 10456 16526
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 11072 15570 11100 19382
rect 11152 17264 11204 17270
rect 11256 17241 11284 19858
rect 11532 19854 11560 20470
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 11612 19916 11664 19922
rect 11612 19858 11664 19864
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11428 19236 11480 19242
rect 11428 19178 11480 19184
rect 11440 18766 11468 19178
rect 11624 18970 11652 19858
rect 11716 19378 11744 20266
rect 11900 19990 11928 20878
rect 11980 20800 12032 20806
rect 11980 20742 12032 20748
rect 11888 19984 11940 19990
rect 11888 19926 11940 19932
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11886 19000 11942 19009
rect 11612 18964 11664 18970
rect 11886 18935 11942 18944
rect 11612 18906 11664 18912
rect 11900 18902 11928 18935
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11992 18290 12020 20742
rect 13188 20482 13216 21082
rect 13004 20466 13216 20482
rect 13280 20466 13308 21286
rect 13004 20460 13228 20466
rect 13004 20454 13176 20460
rect 12900 20392 12952 20398
rect 12820 20340 12900 20346
rect 12820 20334 12952 20340
rect 12820 20318 12940 20334
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12360 19446 12388 19790
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12084 18834 12112 19382
rect 12820 19174 12848 20318
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12622 18864 12678 18873
rect 12072 18828 12124 18834
rect 12622 18799 12678 18808
rect 12072 18770 12124 18776
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 12176 18426 12204 18634
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 12636 18154 12664 18799
rect 12900 18284 12952 18290
rect 13004 18272 13032 20454
rect 13176 20402 13228 20408
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 13096 19334 13124 20334
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13096 19306 13216 19334
rect 13188 18766 13216 19306
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13188 18630 13216 18702
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13188 18290 13216 18566
rect 13372 18358 13400 19110
rect 13360 18352 13412 18358
rect 13360 18294 13412 18300
rect 12952 18244 13032 18272
rect 13176 18284 13228 18290
rect 12900 18226 12952 18232
rect 13176 18226 13228 18232
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 13280 17882 13308 18226
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 11152 17206 11204 17212
rect 11242 17232 11298 17241
rect 11164 16522 11192 17206
rect 11242 17167 11298 17176
rect 12808 16720 12860 16726
rect 12808 16662 12860 16668
rect 13450 16688 13506 16697
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11716 16114 11744 16390
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7116 4758 7144 7822
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 5998 2952 6054 2961
rect 5998 2887 6054 2896
rect 6184 944 6236 950
rect 6184 886 6236 892
rect 6196 800 6224 886
rect 6472 800 6500 4150
rect 6918 3224 6974 3233
rect 6918 3159 6974 3168
rect 6932 2854 6960 3159
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6840 1850 6868 2246
rect 6932 1970 6960 2314
rect 6920 1964 6972 1970
rect 6920 1906 6972 1912
rect 6840 1822 6960 1850
rect 6736 1012 6788 1018
rect 6736 954 6788 960
rect 6748 800 6776 954
rect 6932 950 6960 1822
rect 6920 944 6972 950
rect 6920 886 6972 892
rect 7024 800 7052 4558
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7116 3194 7144 3402
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7208 2650 7236 9386
rect 7930 7984 7986 7993
rect 7930 7919 7986 7928
rect 7944 7886 7972 7919
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7116 1766 7144 2314
rect 7104 1760 7156 1766
rect 7104 1702 7156 1708
rect 7300 800 7328 3334
rect 7392 2854 7420 7142
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7484 3738 7512 3878
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7576 3670 7604 4422
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7576 800 7604 2926
rect 7668 2825 7696 2994
rect 7654 2816 7710 2825
rect 7654 2751 7710 2760
rect 7852 2582 7880 5782
rect 7944 2854 7972 6054
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8128 4826 8156 5170
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8036 2854 8064 2994
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 7668 2106 7696 2314
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7760 2038 7788 2246
rect 7748 2032 7800 2038
rect 7748 1974 7800 1980
rect 7852 800 7880 2382
rect 8128 800 8156 4014
rect 8220 3466 8248 4082
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8220 3126 8248 3402
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8312 1442 8340 4490
rect 8404 4146 8432 4966
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8404 2582 8432 3946
rect 8496 2650 8524 10134
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8772 7886 8800 9454
rect 8956 7954 8984 11018
rect 9680 10736 9732 10742
rect 9586 10704 9642 10713
rect 9496 10668 9548 10674
rect 9680 10678 9732 10684
rect 9586 10639 9588 10648
rect 9496 10610 9548 10616
rect 9640 10639 9642 10648
rect 9588 10610 9640 10616
rect 9508 10418 9536 10610
rect 9588 10464 9640 10470
rect 9508 10412 9588 10418
rect 9508 10406 9640 10412
rect 9508 10390 9628 10406
rect 9692 9518 9720 10678
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8772 7478 8800 7822
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8772 6866 8800 7414
rect 9876 7274 9904 7754
rect 10060 7750 10088 13738
rect 10152 13530 10180 15438
rect 11072 15026 11100 15506
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10244 12434 10272 14214
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10520 12442 10548 12786
rect 10508 12436 10560 12442
rect 10244 12406 10364 12434
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9140 6458 9168 6734
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 5914 9168 6258
rect 9508 6254 9536 6598
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9324 5710 9352 6190
rect 9508 5710 9536 6190
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9508 5166 9536 5646
rect 9600 5370 9628 5646
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9770 4720 9826 4729
rect 9876 4690 9904 7210
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 10060 5166 10088 5578
rect 10152 5234 10180 7822
rect 10336 5574 10364 12406
rect 10508 12378 10560 12384
rect 10612 12238 10640 13194
rect 10704 12238 10732 13194
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11830 10732 12174
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10888 10441 10916 14758
rect 11440 14482 11468 14826
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11164 12850 11192 13670
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11624 12442 11652 13738
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 10968 10464 11020 10470
rect 10874 10432 10930 10441
rect 10968 10406 11020 10412
rect 10874 10367 10930 10376
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10612 7546 10640 8434
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10796 7410 10824 9386
rect 10980 9382 11008 10406
rect 11072 9518 11100 11834
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11164 11218 11192 11562
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11348 11218 11376 11494
rect 11808 11286 11836 13942
rect 11900 12986 11928 14282
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11992 13190 12020 13942
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11992 12866 12020 13126
rect 11900 12838 12020 12866
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11900 11218 11928 12838
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11992 12238 12020 12582
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 12084 11694 12112 15506
rect 12268 14890 12296 16526
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12636 15434 12664 15846
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12256 13864 12308 13870
rect 12176 13824 12256 13852
rect 12176 13190 12204 13824
rect 12256 13806 12308 13812
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 12360 13258 12388 13738
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12176 12434 12204 13126
rect 12452 12850 12480 14010
rect 12636 13734 12664 14962
rect 12728 14074 12756 14962
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12636 13326 12664 13670
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12176 12406 12296 12434
rect 12268 11694 12296 12406
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12084 11558 12112 11630
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11348 10674 11376 11154
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10704 6866 10732 7346
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10796 6746 10824 7346
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10888 6934 10916 7278
rect 10980 7274 11008 7482
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10876 6792 10928 6798
rect 10796 6740 10876 6746
rect 10796 6734 10928 6740
rect 10796 6718 10916 6734
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10244 5370 10272 5510
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9770 4655 9772 4664
rect 9824 4655 9826 4664
rect 9864 4684 9916 4690
rect 9772 4626 9824 4632
rect 9864 4626 9916 4632
rect 10060 4622 10088 5102
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8588 3670 8616 4490
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8576 3664 8628 3670
rect 8576 3606 8628 3612
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8588 2774 8616 3130
rect 8680 2922 8708 3878
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8864 2774 8892 4218
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9324 4078 9352 4150
rect 8944 4072 8996 4078
rect 8942 4040 8944 4049
rect 9128 4072 9180 4078
rect 8996 4040 8998 4049
rect 9128 4014 9180 4020
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 8942 3975 8998 3984
rect 8588 2746 8708 2774
rect 8864 2746 8984 2774
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 8312 1414 8432 1442
rect 8404 800 8432 1414
rect 8680 800 8708 2746
rect 8956 800 8984 2746
rect 9140 1902 9168 4014
rect 9324 3398 9352 4014
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9310 3088 9366 3097
rect 9220 3052 9272 3058
rect 9310 3023 9366 3032
rect 9220 2994 9272 3000
rect 9128 1896 9180 1902
rect 9128 1838 9180 1844
rect 9232 800 9260 2994
rect 9324 2990 9352 3023
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9416 1698 9444 3878
rect 9508 3466 9536 4014
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9494 3088 9550 3097
rect 9600 3074 9628 3470
rect 9550 3046 9628 3074
rect 9494 3023 9496 3032
rect 9548 3023 9550 3032
rect 9496 2994 9548 3000
rect 9692 2774 9720 4558
rect 10428 4078 10456 6190
rect 11072 5914 11100 7278
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10612 5166 10640 5578
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 10612 4622 10640 5102
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9784 3058 9812 3946
rect 10888 3738 10916 5102
rect 11164 4282 11192 10406
rect 11348 10062 11376 10610
rect 11440 10266 11468 11086
rect 12176 10810 12204 11630
rect 12820 11014 12848 16662
rect 13450 16623 13452 16632
rect 13504 16623 13506 16632
rect 13452 16594 13504 16600
rect 13360 16584 13412 16590
rect 13358 16552 13360 16561
rect 13412 16552 13414 16561
rect 13358 16487 13414 16496
rect 13372 16114 13400 16487
rect 13556 16250 13584 19790
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13268 15496 13320 15502
rect 13372 15484 13400 16050
rect 13320 15456 13400 15484
rect 13268 15438 13320 15444
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 11428 10260 11480 10266
rect 11428 10202 11480 10208
rect 12820 10062 12848 10610
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11256 4826 11284 6734
rect 11348 6730 11376 7346
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11716 6662 11744 9998
rect 12820 9586 12848 9998
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12360 9042 12388 9454
rect 13004 9330 13032 14826
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13372 12170 13400 13874
rect 13464 13326 13492 14758
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 13360 12164 13412 12170
rect 13360 12106 13412 12112
rect 13188 11218 13216 12106
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 12728 9302 13032 9330
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12636 7954 12664 8842
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12532 7812 12584 7818
rect 12532 7754 12584 7760
rect 12544 7546 12572 7754
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12636 7410 12664 7890
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12636 7002 12664 7346
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 12636 6322 12664 6938
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12728 5642 12756 9302
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11992 5098 12020 5306
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 12072 5092 12124 5098
rect 12072 5034 12124 5040
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11704 4208 11756 4214
rect 11704 4150 11756 4156
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9876 3194 9904 3470
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 10876 2848 10928 2854
rect 10322 2816 10378 2825
rect 9692 2746 9812 2774
rect 10876 2790 10928 2796
rect 10322 2751 10378 2760
rect 9404 1692 9456 1698
rect 9404 1634 9456 1640
rect 9496 944 9548 950
rect 9496 886 9548 892
rect 9508 800 9536 886
rect 9784 800 9812 2746
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10152 1698 10180 2382
rect 10140 1692 10192 1698
rect 10140 1634 10192 1640
rect 10048 1624 10100 1630
rect 10048 1566 10100 1572
rect 10060 800 10088 1566
rect 10336 800 10364 2751
rect 10600 1964 10652 1970
rect 10600 1906 10652 1912
rect 10612 800 10640 1906
rect 10888 800 10916 2790
rect 11072 2582 11100 3674
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11256 2446 11284 4082
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11072 1018 11100 2246
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11060 1012 11112 1018
rect 11060 954 11112 960
rect 11164 800 11192 2042
rect 11428 1692 11480 1698
rect 11428 1634 11480 1640
rect 11440 800 11468 1634
rect 11716 800 11744 4150
rect 11992 800 12020 4422
rect 12084 3670 12112 5034
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 12268 800 12296 5170
rect 12728 4706 12756 5578
rect 12636 4678 12756 4706
rect 12348 4208 12400 4214
rect 12400 4168 12480 4196
rect 12348 4150 12400 4156
rect 12452 2774 12480 4168
rect 12532 3664 12584 3670
rect 12636 3641 12664 4678
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12728 4010 12756 4558
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12820 3890 12848 7958
rect 12912 7342 12940 8230
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12900 4072 12952 4078
rect 12898 4040 12900 4049
rect 12952 4040 12954 4049
rect 12898 3975 12954 3984
rect 12728 3862 12848 3890
rect 12532 3606 12584 3612
rect 12622 3632 12678 3641
rect 12544 3194 12572 3606
rect 12622 3567 12678 3576
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12452 2746 12572 2774
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12360 2106 12388 2382
rect 12348 2100 12400 2106
rect 12348 2042 12400 2048
rect 12544 800 12572 2746
rect 12636 1086 12664 3402
rect 12728 2038 12756 3862
rect 13004 3754 13032 9046
rect 13096 4706 13124 10950
rect 13188 10538 13216 11154
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13188 10198 13216 10474
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13452 10056 13504 10062
rect 13266 10024 13322 10033
rect 13452 9998 13504 10004
rect 13266 9959 13322 9968
rect 13280 9110 13308 9959
rect 13464 9586 13492 9998
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13464 8974 13492 9522
rect 13648 9217 13676 61066
rect 14292 60790 14320 63294
rect 14830 63294 14964 63322
rect 14830 63200 14886 63294
rect 14936 61198 14964 63294
rect 15566 63294 15792 63322
rect 15566 63200 15622 63294
rect 14924 61192 14976 61198
rect 14924 61134 14976 61140
rect 15200 61124 15252 61130
rect 15200 61066 15252 61072
rect 14280 60784 14332 60790
rect 14280 60726 14332 60732
rect 15108 60512 15160 60518
rect 15108 60454 15160 60460
rect 15120 60246 15148 60454
rect 15108 60240 15160 60246
rect 15108 60182 15160 60188
rect 15212 47569 15240 61066
rect 15764 60790 15792 63294
rect 16132 63294 16358 63322
rect 16132 61198 16160 63294
rect 16302 63200 16358 63294
rect 17038 63322 17094 64000
rect 17774 63322 17830 64000
rect 18510 63322 18566 64000
rect 19246 63322 19302 64000
rect 19982 63322 20038 64000
rect 17038 63294 17172 63322
rect 17038 63200 17094 63294
rect 17144 61198 17172 63294
rect 17774 63294 18000 63322
rect 17774 63200 17830 63294
rect 17868 61600 17920 61606
rect 17868 61542 17920 61548
rect 16120 61192 16172 61198
rect 16120 61134 16172 61140
rect 17132 61192 17184 61198
rect 17132 61134 17184 61140
rect 17500 61124 17552 61130
rect 17500 61066 17552 61072
rect 17316 61056 17368 61062
rect 17316 60998 17368 61004
rect 15752 60784 15804 60790
rect 15752 60726 15804 60732
rect 15198 47560 15254 47569
rect 15198 47495 15254 47504
rect 15200 45824 15252 45830
rect 15200 45766 15252 45772
rect 15212 45558 15240 45766
rect 15200 45552 15252 45558
rect 15200 45494 15252 45500
rect 16212 38548 16264 38554
rect 16212 38490 16264 38496
rect 16224 38010 16252 38490
rect 16212 38004 16264 38010
rect 16212 37946 16264 37952
rect 16672 37868 16724 37874
rect 16672 37810 16724 37816
rect 16580 36780 16632 36786
rect 16580 36722 16632 36728
rect 16592 32774 16620 36722
rect 16684 36106 16712 37810
rect 16672 36100 16724 36106
rect 16672 36042 16724 36048
rect 16580 32768 16632 32774
rect 16580 32710 16632 32716
rect 16684 31090 16712 36042
rect 17328 34134 17356 60998
rect 17512 45558 17540 61066
rect 17880 60722 17908 61542
rect 17972 61198 18000 63294
rect 18510 63294 18736 63322
rect 18510 63200 18566 63294
rect 18052 61260 18104 61266
rect 18052 61202 18104 61208
rect 17960 61192 18012 61198
rect 17960 61134 18012 61140
rect 17868 60716 17920 60722
rect 17868 60658 17920 60664
rect 17868 60512 17920 60518
rect 17868 60454 17920 60460
rect 17880 60178 17908 60454
rect 17868 60172 17920 60178
rect 17868 60114 17920 60120
rect 17592 59968 17644 59974
rect 17592 59910 17644 59916
rect 17604 50289 17632 59910
rect 18064 59634 18092 61202
rect 18708 61198 18736 63294
rect 19246 63294 19472 63322
rect 19246 63200 19302 63294
rect 19340 61328 19392 61334
rect 19340 61270 19392 61276
rect 18696 61192 18748 61198
rect 18696 61134 18748 61140
rect 18788 61056 18840 61062
rect 18788 60998 18840 61004
rect 18420 60648 18472 60654
rect 18420 60590 18472 60596
rect 18144 60172 18196 60178
rect 18144 60114 18196 60120
rect 18052 59628 18104 59634
rect 18052 59570 18104 59576
rect 17868 51944 17920 51950
rect 17868 51886 17920 51892
rect 17590 50280 17646 50289
rect 17590 50215 17646 50224
rect 17880 48278 17908 51886
rect 17868 48272 17920 48278
rect 17868 48214 17920 48220
rect 17500 45552 17552 45558
rect 17500 45494 17552 45500
rect 17776 45280 17828 45286
rect 17776 45222 17828 45228
rect 17316 34128 17368 34134
rect 17316 34070 17368 34076
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 16592 31062 16712 31090
rect 15660 21616 15712 21622
rect 15660 21558 15712 21564
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14004 20800 14056 20806
rect 14004 20742 14056 20748
rect 14016 20466 14044 20742
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13740 19990 13768 20334
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13924 18970 13952 19110
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 14108 18154 14136 21490
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 15200 21072 15252 21078
rect 15200 21014 15252 21020
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14200 19378 14228 20198
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14096 18148 14148 18154
rect 14096 18090 14148 18096
rect 14292 17882 14320 20878
rect 15212 20534 15240 21014
rect 15396 20942 15424 21422
rect 15384 20936 15436 20942
rect 15384 20878 15436 20884
rect 15292 20800 15344 20806
rect 15292 20742 15344 20748
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 15304 20466 15332 20742
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14384 19378 14412 19790
rect 15488 19786 15516 20198
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14832 18828 14884 18834
rect 14832 18770 14884 18776
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14476 18193 14504 18226
rect 14462 18184 14518 18193
rect 14462 18119 14518 18128
rect 14556 18148 14608 18154
rect 14476 18086 14504 18119
rect 14556 18090 14608 18096
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 13818 16144 13874 16153
rect 13924 16114 13952 16458
rect 13818 16079 13820 16088
rect 13872 16079 13874 16088
rect 13912 16108 13964 16114
rect 13820 16050 13872 16056
rect 13912 16050 13964 16056
rect 13924 15586 13952 16050
rect 14096 16040 14148 16046
rect 14096 15982 14148 15988
rect 13832 15570 13952 15586
rect 13820 15564 13952 15570
rect 13872 15558 13952 15564
rect 13820 15506 13872 15512
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13740 13394 13768 14758
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 11898 13860 12786
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13634 9208 13690 9217
rect 13634 9143 13690 9152
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13464 8634 13492 8910
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13832 8022 13860 11154
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13372 5234 13400 6394
rect 13924 5370 13952 15438
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 14016 12986 14044 14418
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10266 14044 10610
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14016 8498 14044 10202
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13096 4678 13216 4706
rect 13372 4690 13400 5170
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13464 4758 13492 4966
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 12820 3726 13032 3754
rect 12716 2032 12768 2038
rect 12716 1974 12768 1980
rect 12820 1766 12848 3726
rect 12990 3632 13046 3641
rect 12990 3567 13046 3576
rect 13004 2446 13032 3567
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 12808 1760 12860 1766
rect 12808 1702 12860 1708
rect 12624 1080 12676 1086
rect 12624 1022 12676 1028
rect 12808 1012 12860 1018
rect 12808 954 12860 960
rect 12820 800 12848 954
rect 13096 800 13124 4490
rect 13188 3194 13216 4678
rect 13360 4684 13412 4690
rect 13360 4626 13412 4632
rect 13372 4214 13400 4626
rect 13360 4208 13412 4214
rect 13280 4168 13360 4196
rect 13280 3466 13308 4168
rect 13360 4150 13412 4156
rect 13268 3460 13320 3466
rect 13268 3402 13320 3408
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13280 2990 13308 3402
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13372 800 13400 3334
rect 13556 2990 13584 4966
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13740 3738 13768 3946
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 13464 1154 13492 2314
rect 13452 1148 13504 1154
rect 13452 1090 13504 1096
rect 13648 800 13676 2586
rect 13740 950 13768 2994
rect 13728 944 13780 950
rect 13728 886 13780 892
rect 13924 800 13952 5170
rect 14108 3602 14136 15982
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14200 14482 14228 14962
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14200 13938 14228 14418
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14292 13530 14320 15438
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14384 13410 14412 14962
rect 14476 14958 14504 15302
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14568 14804 14596 18090
rect 14844 17678 14872 18770
rect 15120 17678 15148 19654
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 15212 17882 15240 19314
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15304 17202 15332 18022
rect 15396 17338 15424 19654
rect 15580 19446 15608 19722
rect 15568 19440 15620 19446
rect 15568 19382 15620 19388
rect 15580 18766 15608 19382
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15488 18426 15516 18634
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15580 17202 15608 18702
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 14200 13382 14412 13410
rect 14476 14776 14596 14804
rect 15016 14816 15068 14822
rect 14200 12442 14228 13382
rect 14476 13274 14504 14776
rect 15016 14758 15068 14764
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14384 13246 14504 13274
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14384 11762 14412 13246
rect 14568 12918 14596 13874
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14556 12912 14608 12918
rect 14556 12854 14608 12860
rect 14844 12442 14872 13806
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 15028 12306 15056 14758
rect 15108 13320 15160 13326
rect 15212 13274 15240 15846
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15488 15162 15516 15302
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15488 13734 15516 15098
rect 15568 14272 15620 14278
rect 15568 14214 15620 14220
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15160 13268 15240 13274
rect 15108 13262 15240 13268
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15120 13246 15240 13262
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15212 12986 15240 13126
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15108 12844 15160 12850
rect 15304 12832 15332 13262
rect 15396 12918 15424 13262
rect 15488 12986 15516 13262
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15160 12804 15332 12832
rect 15108 12786 15160 12792
rect 15120 12753 15148 12786
rect 15106 12744 15162 12753
rect 15396 12714 15424 12854
rect 15106 12679 15162 12688
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 15580 12434 15608 14214
rect 15304 12406 15608 12434
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11762 14504 12038
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14936 10674 14964 11834
rect 15212 11354 15240 12106
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14752 10198 14780 10610
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14740 10192 14792 10198
rect 14740 10134 14792 10140
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14476 9586 14504 9930
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 14200 3670 14228 4490
rect 14188 3664 14240 3670
rect 14188 3606 14240 3612
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14188 1080 14240 1086
rect 14188 1022 14240 1028
rect 14200 800 14228 1022
rect 14292 1018 14320 2926
rect 14384 2038 14412 9318
rect 14752 7954 14780 10134
rect 14844 10062 14872 10406
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14936 9874 14964 10610
rect 15200 9920 15252 9926
rect 15198 9888 15200 9897
rect 15252 9888 15254 9897
rect 14936 9846 15148 9874
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14936 8906 14964 9386
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 15120 8838 15148 9846
rect 15198 9823 15254 9832
rect 15304 9674 15332 12406
rect 15672 12322 15700 21558
rect 16396 21412 16448 21418
rect 16396 21354 16448 21360
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 16224 20602 16252 20810
rect 16212 20596 16264 20602
rect 16212 20538 16264 20544
rect 16408 19990 16436 21354
rect 16592 21350 16620 31062
rect 16776 26234 16804 31758
rect 17788 30666 17816 45222
rect 17776 30660 17828 30666
rect 17776 30602 17828 30608
rect 16684 26206 16804 26234
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16396 19984 16448 19990
rect 16396 19926 16448 19932
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 16592 18970 16620 19314
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16224 16794 16252 17614
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16408 16590 16436 18362
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15764 13530 15792 16050
rect 16486 16008 16542 16017
rect 16486 15943 16542 15952
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15488 12294 15700 12322
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15396 10266 15424 11494
rect 15488 10606 15516 12294
rect 15856 12238 15884 13126
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15304 9646 15424 9674
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 14844 8129 14872 8774
rect 15120 8634 15148 8774
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15304 8430 15332 8570
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 14830 8120 14886 8129
rect 14830 8055 14886 8064
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15120 7478 15148 7890
rect 15304 7886 15332 8366
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15108 7472 15160 7478
rect 15200 7472 15252 7478
rect 15108 7414 15160 7420
rect 15198 7440 15200 7449
rect 15252 7440 15254 7449
rect 15120 6934 15148 7414
rect 15198 7375 15254 7384
rect 15304 7342 15332 7822
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15108 6928 15160 6934
rect 15108 6870 15160 6876
rect 15120 6474 15148 6870
rect 15120 6446 15240 6474
rect 15212 6390 15240 6446
rect 15396 6440 15424 9646
rect 15488 9586 15516 9930
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15580 9450 15608 11766
rect 15764 11354 15792 12174
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15658 11248 15714 11257
rect 15658 11183 15714 11192
rect 15672 11082 15700 11183
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15304 6412 15424 6440
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15304 6202 15332 6412
rect 15382 6352 15438 6361
rect 15382 6287 15384 6296
rect 15436 6287 15438 6296
rect 15384 6258 15436 6264
rect 15304 6174 15424 6202
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14476 3058 14504 5510
rect 14922 5264 14978 5273
rect 14922 5199 14978 5208
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14830 4720 14886 4729
rect 14568 4282 14596 4694
rect 14830 4655 14886 4664
rect 14738 4584 14794 4593
rect 14738 4519 14794 4528
rect 14752 4486 14780 4519
rect 14844 4486 14872 4655
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14936 4078 14964 5199
rect 15290 4856 15346 4865
rect 15290 4791 15346 4800
rect 15304 4690 15332 4791
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15396 4622 15424 6174
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15212 4282 15240 4558
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15200 4276 15252 4282
rect 15200 4218 15252 4224
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 14648 3664 14700 3670
rect 14648 3606 14700 3612
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14660 2582 14688 3606
rect 14844 3534 14872 3946
rect 15198 3768 15254 3777
rect 15198 3703 15254 3712
rect 15212 3602 15240 3703
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14830 2952 14886 2961
rect 14830 2887 14886 2896
rect 14844 2854 14872 2887
rect 14832 2848 14884 2854
rect 14832 2790 14884 2796
rect 14648 2576 14700 2582
rect 14648 2518 14700 2524
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 14372 2032 14424 2038
rect 14372 1974 14424 1980
rect 14936 1358 14964 2382
rect 14924 1352 14976 1358
rect 14924 1294 14976 1300
rect 14464 1148 14516 1154
rect 14464 1090 14516 1096
rect 14280 1012 14332 1018
rect 14280 954 14332 960
rect 14476 800 14504 1090
rect 14740 944 14792 950
rect 14740 886 14792 892
rect 14752 800 14780 886
rect 15028 800 15056 2450
rect 15304 800 15332 4490
rect 15488 2446 15516 9046
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15580 7410 15608 7754
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15580 3194 15608 5306
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15672 2106 15700 11018
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15948 9654 15976 10542
rect 15936 9648 15988 9654
rect 15842 9616 15898 9625
rect 15936 9590 15988 9596
rect 15842 9551 15844 9560
rect 15896 9551 15898 9560
rect 15844 9522 15896 9528
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15856 7478 15884 7822
rect 15844 7472 15896 7478
rect 15896 7420 15976 7426
rect 15844 7414 15976 7420
rect 15856 7398 15976 7414
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15750 6896 15806 6905
rect 15750 6831 15752 6840
rect 15804 6831 15806 6840
rect 15752 6802 15804 6808
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 6322 15792 6598
rect 15856 6322 15884 7278
rect 15948 6866 15976 7398
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15948 6322 15976 6802
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 15934 6216 15990 6225
rect 15934 6151 15990 6160
rect 15844 4072 15896 4078
rect 15844 4014 15896 4020
rect 15856 3602 15884 4014
rect 15948 3942 15976 6151
rect 16040 5370 16068 13806
rect 16132 12442 16160 15438
rect 16500 15434 16528 15943
rect 16488 15428 16540 15434
rect 16488 15370 16540 15376
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14074 16252 14758
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16120 12436 16172 12442
rect 16500 12434 16528 15098
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16592 13462 16620 13738
rect 16580 13456 16632 13462
rect 16580 13398 16632 13404
rect 16684 12434 16712 26206
rect 17684 24336 17736 24342
rect 17684 24278 17736 24284
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16776 19802 16804 21286
rect 16960 20534 16988 22374
rect 17316 22092 17368 22098
rect 17696 22094 17724 24278
rect 18052 22636 18104 22642
rect 18052 22578 18104 22584
rect 17960 22160 18012 22166
rect 17960 22102 18012 22108
rect 17316 22034 17368 22040
rect 17604 22066 17724 22094
rect 17328 21146 17356 22034
rect 17408 21956 17460 21962
rect 17408 21898 17460 21904
rect 17420 21486 17448 21898
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 17316 21140 17368 21146
rect 17316 21082 17368 21088
rect 17328 21026 17356 21082
rect 17236 20998 17356 21026
rect 17236 20942 17264 20998
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 17144 20466 17172 20742
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 16868 19922 16896 20402
rect 17314 19952 17370 19961
rect 16856 19916 16908 19922
rect 17314 19887 17370 19896
rect 16856 19858 16908 19864
rect 16776 19774 16896 19802
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16776 17882 16804 18158
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16868 16402 16896 19774
rect 17222 19408 17278 19417
rect 17222 19343 17278 19352
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16960 17882 16988 18702
rect 17052 18290 17080 19246
rect 17236 19009 17264 19343
rect 17328 19174 17356 19887
rect 17512 19854 17540 20742
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17222 19000 17278 19009
rect 17222 18935 17278 18944
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16948 16584 17000 16590
rect 17052 16572 17080 18226
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17144 16590 17172 16934
rect 17000 16544 17080 16572
rect 16948 16526 17000 16532
rect 16868 16374 16988 16402
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16776 15178 16804 15302
rect 16776 15150 16896 15178
rect 16868 15026 16896 15150
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16776 14278 16804 14418
rect 16868 14414 16896 14758
rect 16960 14498 16988 16374
rect 17052 16114 17080 16544
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 17236 16522 17264 16934
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17040 16108 17092 16114
rect 17040 16050 17092 16056
rect 17052 14958 17080 16050
rect 17132 15632 17184 15638
rect 17132 15574 17184 15580
rect 17144 15434 17172 15574
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 17052 14618 17080 14894
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 16960 14470 17080 14498
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 13938 16804 14214
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16762 13832 16818 13841
rect 16762 13767 16818 13776
rect 16120 12378 16172 12384
rect 16408 12406 16528 12434
rect 16592 12406 16712 12434
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16316 11150 16344 11494
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16120 10532 16172 10538
rect 16120 10474 16172 10480
rect 16132 10062 16160 10474
rect 16408 10418 16436 12406
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16500 11286 16528 11494
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16316 10390 16436 10418
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16132 7886 16160 9998
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16224 8430 16252 9522
rect 16316 9110 16344 10390
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16408 10062 16436 10202
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16500 9926 16528 10202
rect 16592 9926 16620 12406
rect 16670 12336 16726 12345
rect 16670 12271 16726 12280
rect 16684 11150 16712 12271
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 16684 10062 16712 10134
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16488 9920 16540 9926
rect 16394 9888 16450 9897
rect 16488 9862 16540 9868
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16394 9823 16450 9832
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16316 8566 16344 8910
rect 16304 8560 16356 8566
rect 16304 8502 16356 8508
rect 16316 8430 16344 8502
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16408 6866 16436 9823
rect 16684 8974 16712 9998
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16684 8838 16712 8910
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16488 7744 16540 7750
rect 16540 7704 16712 7732
rect 16488 7686 16540 7692
rect 16684 7478 16712 7704
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 16132 4826 16160 6666
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16592 5778 16620 6598
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16132 4078 16160 4762
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15842 3496 15898 3505
rect 15842 3431 15898 3440
rect 15856 3058 15884 3431
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16040 2774 16068 2926
rect 16040 2746 16160 2774
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15660 2100 15712 2106
rect 15660 2042 15712 2048
rect 15568 1012 15620 1018
rect 15568 954 15620 960
rect 15580 800 15608 954
rect 15856 800 15884 2246
rect 16132 800 16160 2746
rect 16316 1018 16344 2926
rect 16592 2774 16620 5034
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16408 2746 16620 2774
rect 16304 1012 16356 1018
rect 16304 954 16356 960
rect 16408 800 16436 2746
rect 16684 800 16712 4966
rect 16776 3534 16804 13767
rect 16868 11150 16896 14010
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16960 12238 16988 13126
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16868 10470 16896 11086
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16868 8022 16896 9862
rect 16960 8906 16988 10542
rect 17052 10198 17080 14470
rect 17604 14074 17632 22066
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17880 21622 17908 21966
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 17972 20874 18000 22102
rect 18064 21298 18092 22578
rect 18156 22094 18184 60114
rect 18432 60110 18460 60590
rect 18420 60104 18472 60110
rect 18420 60046 18472 60052
rect 18512 60104 18564 60110
rect 18512 60046 18564 60052
rect 18524 58886 18552 60046
rect 18512 58880 18564 58886
rect 18512 58822 18564 58828
rect 18800 35766 18828 60998
rect 19248 60240 19300 60246
rect 19248 60182 19300 60188
rect 19156 60036 19208 60042
rect 19156 59978 19208 59984
rect 19168 59702 19196 59978
rect 19156 59696 19208 59702
rect 19156 59638 19208 59644
rect 19260 59430 19288 60182
rect 19352 59650 19380 61270
rect 19444 60790 19472 63294
rect 19812 63294 20038 63322
rect 19812 61198 19840 63294
rect 19982 63200 20038 63294
rect 20718 63200 20774 64000
rect 21454 63322 21510 64000
rect 21284 63294 21510 63322
rect 20732 61198 20760 63200
rect 21284 61198 21312 63294
rect 21454 63200 21510 63294
rect 22190 63200 22246 64000
rect 22926 63322 22982 64000
rect 22926 63294 23244 63322
rect 22926 63200 22982 63294
rect 22100 61328 22152 61334
rect 22100 61270 22152 61276
rect 19800 61192 19852 61198
rect 19800 61134 19852 61140
rect 20720 61192 20772 61198
rect 20720 61134 20772 61140
rect 21272 61192 21324 61198
rect 21272 61134 21324 61140
rect 19984 61124 20036 61130
rect 19984 61066 20036 61072
rect 21180 61124 21232 61130
rect 21180 61066 21232 61072
rect 19574 60956 19882 60965
rect 19574 60954 19580 60956
rect 19636 60954 19660 60956
rect 19716 60954 19740 60956
rect 19796 60954 19820 60956
rect 19876 60954 19882 60956
rect 19636 60902 19638 60954
rect 19818 60902 19820 60954
rect 19574 60900 19580 60902
rect 19636 60900 19660 60902
rect 19716 60900 19740 60902
rect 19796 60900 19820 60902
rect 19876 60900 19882 60902
rect 19574 60891 19882 60900
rect 19432 60784 19484 60790
rect 19432 60726 19484 60732
rect 19616 60648 19668 60654
rect 19616 60590 19668 60596
rect 19628 60110 19656 60590
rect 19996 60110 20024 61066
rect 20996 61056 21048 61062
rect 20996 60998 21048 61004
rect 20076 60512 20128 60518
rect 20076 60454 20128 60460
rect 19616 60104 19668 60110
rect 19616 60046 19668 60052
rect 19892 60104 19944 60110
rect 19892 60046 19944 60052
rect 19984 60104 20036 60110
rect 19984 60046 20036 60052
rect 19904 59974 19932 60046
rect 19892 59968 19944 59974
rect 19892 59910 19944 59916
rect 19984 59968 20036 59974
rect 19984 59910 20036 59916
rect 19574 59868 19882 59877
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59803 19882 59812
rect 19996 59770 20024 59910
rect 19984 59764 20036 59770
rect 19984 59706 20036 59712
rect 19352 59622 19748 59650
rect 19248 59424 19300 59430
rect 19248 59366 19300 59372
rect 19524 59152 19576 59158
rect 19524 59094 19576 59100
rect 19536 58970 19564 59094
rect 19720 59022 19748 59622
rect 19352 58942 19564 58970
rect 19708 59016 19760 59022
rect 20088 58970 20116 60454
rect 20260 60308 20312 60314
rect 20260 60250 20312 60256
rect 20168 60240 20220 60246
rect 20168 60182 20220 60188
rect 19708 58958 19760 58964
rect 19996 58942 20116 58970
rect 19248 38276 19300 38282
rect 19248 38218 19300 38224
rect 19260 37466 19288 38218
rect 19352 37874 19380 58942
rect 19574 58780 19882 58789
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58715 19882 58724
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19996 38826 20024 58942
rect 20076 58880 20128 58886
rect 20076 58822 20128 58828
rect 19984 38820 20036 38826
rect 19984 38762 20036 38768
rect 19432 38752 19484 38758
rect 20088 38706 20116 58822
rect 19432 38694 19484 38700
rect 19444 37890 19472 38694
rect 19996 38678 20116 38706
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19708 37936 19760 37942
rect 19444 37884 19708 37890
rect 19444 37878 19760 37884
rect 19996 37890 20024 38678
rect 20180 38282 20208 60182
rect 20272 52154 20300 60250
rect 20812 60036 20864 60042
rect 20812 59978 20864 59984
rect 20904 60036 20956 60042
rect 20904 59978 20956 59984
rect 20824 59566 20852 59978
rect 20916 59770 20944 59978
rect 20904 59764 20956 59770
rect 20904 59706 20956 59712
rect 20812 59560 20864 59566
rect 20812 59502 20864 59508
rect 20260 52148 20312 52154
rect 20260 52090 20312 52096
rect 20536 51808 20588 51814
rect 20536 51750 20588 51756
rect 20548 38962 20576 51750
rect 21008 45554 21036 60998
rect 21192 59634 21220 61066
rect 22008 61056 22060 61062
rect 22008 60998 22060 61004
rect 21916 60240 21968 60246
rect 21916 60182 21968 60188
rect 21272 59968 21324 59974
rect 21272 59910 21324 59916
rect 21824 59968 21876 59974
rect 21824 59910 21876 59916
rect 21284 59634 21312 59910
rect 21364 59696 21416 59702
rect 21364 59638 21416 59644
rect 21180 59628 21232 59634
rect 21180 59570 21232 59576
rect 21272 59628 21324 59634
rect 21272 59570 21324 59576
rect 21284 53514 21312 59570
rect 21376 59022 21404 59638
rect 21836 59401 21864 59910
rect 21822 59392 21878 59401
rect 21822 59327 21878 59336
rect 21364 59016 21416 59022
rect 21364 58958 21416 58964
rect 21272 53508 21324 53514
rect 21272 53450 21324 53456
rect 21376 45554 21404 58958
rect 21456 52420 21508 52426
rect 21456 52362 21508 52368
rect 20916 45526 21036 45554
rect 21284 45526 21404 45554
rect 20916 40186 20944 45526
rect 21088 45484 21140 45490
rect 21088 45426 21140 45432
rect 20904 40180 20956 40186
rect 20904 40122 20956 40128
rect 21100 40118 21128 45426
rect 21284 44946 21312 45526
rect 21468 45422 21496 52362
rect 21456 45416 21508 45422
rect 21456 45358 21508 45364
rect 21272 44940 21324 44946
rect 21272 44882 21324 44888
rect 21180 40928 21232 40934
rect 21180 40870 21232 40876
rect 21192 40118 21220 40870
rect 21088 40112 21140 40118
rect 21088 40054 21140 40060
rect 21180 40112 21232 40118
rect 21180 40054 21232 40060
rect 20536 38956 20588 38962
rect 20536 38898 20588 38904
rect 20260 38820 20312 38826
rect 20260 38762 20312 38768
rect 20168 38276 20220 38282
rect 20168 38218 20220 38224
rect 19340 37868 19392 37874
rect 19444 37862 19748 37878
rect 19996 37862 20116 37890
rect 19340 37810 19392 37816
rect 19800 37732 19852 37738
rect 19800 37674 19852 37680
rect 19248 37460 19300 37466
rect 19248 37402 19300 37408
rect 19812 37398 19840 37674
rect 19984 37664 20036 37670
rect 19984 37606 20036 37612
rect 19800 37392 19852 37398
rect 19800 37334 19852 37340
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 18880 37188 18932 37194
rect 18880 37130 18932 37136
rect 18892 36786 18920 37130
rect 18880 36780 18932 36786
rect 18880 36722 18932 36728
rect 19248 36712 19300 36718
rect 19248 36654 19300 36660
rect 18788 35760 18840 35766
rect 18788 35702 18840 35708
rect 18880 35692 18932 35698
rect 18880 35634 18932 35640
rect 18892 35494 18920 35634
rect 18880 35488 18932 35494
rect 18880 35430 18932 35436
rect 18788 30252 18840 30258
rect 18788 30194 18840 30200
rect 18800 29782 18828 30194
rect 18788 29776 18840 29782
rect 18788 29718 18840 29724
rect 18512 26308 18564 26314
rect 18512 26250 18564 26256
rect 18524 22094 18552 26250
rect 18892 24342 18920 35430
rect 19156 30592 19208 30598
rect 19156 30534 19208 30540
rect 19168 30326 19196 30534
rect 19156 30320 19208 30326
rect 19156 30262 19208 30268
rect 19260 30258 19288 36654
rect 18972 30252 19024 30258
rect 18972 30194 19024 30200
rect 19064 30252 19116 30258
rect 19064 30194 19116 30200
rect 19248 30252 19300 30258
rect 19248 30194 19300 30200
rect 18880 24336 18932 24342
rect 18880 24278 18932 24284
rect 18984 24138 19012 30194
rect 19076 29714 19104 30194
rect 19064 29708 19116 29714
rect 19064 29650 19116 29656
rect 19076 29170 19104 29650
rect 19260 29306 19288 30194
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 19064 29164 19116 29170
rect 19064 29106 19116 29112
rect 19076 26234 19104 29106
rect 19352 26234 19380 37198
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36780 19484 36786
rect 19432 36722 19484 36728
rect 19444 34678 19472 36722
rect 19996 36106 20024 37606
rect 19984 36100 20036 36106
rect 19984 36042 20036 36048
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19432 34672 19484 34678
rect 19432 34614 19484 34620
rect 20088 34542 20116 37862
rect 20168 37188 20220 37194
rect 20168 37130 20220 37136
rect 20180 35698 20208 37130
rect 20168 35692 20220 35698
rect 20168 35634 20220 35640
rect 20272 34746 20300 38762
rect 21100 38554 21128 40054
rect 20904 38548 20956 38554
rect 20904 38490 20956 38496
rect 21088 38548 21140 38554
rect 21088 38490 21140 38496
rect 20720 38412 20772 38418
rect 20720 38354 20772 38360
rect 20352 38344 20404 38350
rect 20352 38286 20404 38292
rect 20364 38214 20392 38286
rect 20352 38208 20404 38214
rect 20352 38150 20404 38156
rect 20364 37890 20392 38150
rect 20626 37904 20682 37913
rect 20364 37862 20484 37890
rect 20352 37392 20404 37398
rect 20352 37334 20404 37340
rect 20260 34740 20312 34746
rect 20260 34682 20312 34688
rect 20076 34536 20128 34542
rect 20076 34478 20128 34484
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 20364 33454 20392 37334
rect 20456 37126 20484 37862
rect 20732 37874 20760 38354
rect 20812 38004 20864 38010
rect 20812 37946 20864 37952
rect 20824 37874 20852 37946
rect 20626 37839 20682 37848
rect 20720 37868 20772 37874
rect 20640 37806 20668 37839
rect 20720 37810 20772 37816
rect 20812 37868 20864 37874
rect 20812 37810 20864 37816
rect 20628 37800 20680 37806
rect 20628 37742 20680 37748
rect 20812 37732 20864 37738
rect 20812 37674 20864 37680
rect 20628 37664 20680 37670
rect 20628 37606 20680 37612
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 20444 37120 20496 37126
rect 20444 37062 20496 37068
rect 20352 33448 20404 33454
rect 20352 33390 20404 33396
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 30864 19484 30870
rect 19432 30806 19484 30812
rect 19444 30394 19472 30806
rect 19984 30592 20036 30598
rect 19984 30534 20036 30540
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19076 26206 19196 26234
rect 19352 26206 19472 26234
rect 18972 24132 19024 24138
rect 18972 24074 19024 24080
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 18156 22066 18460 22094
rect 18524 22066 18644 22094
rect 18236 21616 18288 21622
rect 18236 21558 18288 21564
rect 18248 21418 18276 21558
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 18236 21412 18288 21418
rect 18236 21354 18288 21360
rect 18064 21270 18184 21298
rect 18156 21078 18184 21270
rect 18248 21146 18276 21354
rect 18236 21140 18288 21146
rect 18236 21082 18288 21088
rect 18144 21072 18196 21078
rect 18144 21014 18196 21020
rect 18156 20942 18184 21014
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 17960 20868 18012 20874
rect 17960 20810 18012 20816
rect 18248 20602 18276 21082
rect 18340 20806 18368 21490
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 18142 20360 18198 20369
rect 18142 20295 18198 20304
rect 17958 20088 18014 20097
rect 17958 20023 17960 20032
rect 18012 20023 18014 20032
rect 17960 19994 18012 20000
rect 18156 19514 18184 20295
rect 18144 19508 18196 19514
rect 18144 19450 18196 19456
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 18408 18000 18566
rect 18340 18426 18368 19178
rect 18328 18420 18380 18426
rect 17972 18380 18092 18408
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17788 17202 17816 17478
rect 17972 17338 18000 18226
rect 18064 17678 18092 18380
rect 18328 18362 18380 18368
rect 18142 18184 18198 18193
rect 18142 18119 18198 18128
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 18156 17610 18184 18119
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 18326 16960 18382 16969
rect 18326 16895 18382 16904
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17788 15706 17816 16050
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17972 14550 18000 15302
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 17960 14544 18012 14550
rect 17960 14486 18012 14492
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17328 12850 17356 13330
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 11762 17264 12582
rect 17420 11898 17448 13874
rect 17788 13394 17816 14418
rect 18156 14074 18184 15030
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18156 12850 18184 13126
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 17682 12744 17738 12753
rect 17682 12679 17738 12688
rect 17696 12238 17724 12679
rect 18064 12442 18092 12786
rect 18340 12753 18368 16895
rect 18432 16454 18460 22066
rect 18512 20868 18564 20874
rect 18512 20810 18564 20816
rect 18524 20534 18552 20810
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18524 18154 18552 18702
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18432 13326 18460 13670
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18524 13326 18552 13398
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18142 12744 18198 12753
rect 18326 12744 18382 12753
rect 18142 12679 18198 12688
rect 18236 12708 18288 12714
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17972 12102 18000 12242
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17866 11384 17922 11393
rect 17866 11319 17922 11328
rect 17500 11280 17552 11286
rect 17500 11222 17552 11228
rect 17512 11082 17540 11222
rect 17590 11112 17646 11121
rect 17500 11076 17552 11082
rect 17590 11047 17646 11056
rect 17500 11018 17552 11024
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17420 10674 17448 10950
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17130 10568 17186 10577
rect 17236 10538 17264 10610
rect 17130 10503 17186 10512
rect 17224 10532 17276 10538
rect 17040 10192 17092 10198
rect 17040 10134 17092 10140
rect 17144 9110 17172 10503
rect 17224 10474 17276 10480
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17222 10296 17278 10305
rect 17222 10231 17278 10240
rect 17236 10130 17264 10231
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17328 9518 17356 10406
rect 17420 9994 17448 10610
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 17132 9104 17184 9110
rect 17132 9046 17184 9052
rect 17420 8974 17448 9930
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 17316 8900 17368 8906
rect 17316 8842 17368 8848
rect 17328 8616 17356 8842
rect 17512 8634 17540 10610
rect 17408 8628 17460 8634
rect 17328 8588 17408 8616
rect 17408 8570 17460 8576
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 17130 8528 17186 8537
rect 16856 8016 16908 8022
rect 16856 7958 16908 7964
rect 16868 7478 16896 7958
rect 16960 7886 16988 8502
rect 17420 8514 17448 8570
rect 17420 8486 17540 8514
rect 17130 8463 17186 8472
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 17052 7546 17080 7686
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 16960 6798 16988 7414
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16960 800 16988 4966
rect 17144 4146 17172 8463
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17328 6866 17356 7346
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17328 5710 17356 6802
rect 17420 6798 17448 8298
rect 17512 7886 17540 8486
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17512 7546 17540 7822
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17512 6934 17540 7346
rect 17604 7342 17632 11047
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17696 10810 17724 10950
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17682 10160 17738 10169
rect 17682 10095 17738 10104
rect 17696 10062 17724 10095
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 17590 6896 17646 6905
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17512 6322 17540 6870
rect 17590 6831 17646 6840
rect 17604 6798 17632 6831
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17696 5846 17724 9998
rect 17880 9704 17908 11319
rect 17880 9676 18000 9704
rect 17972 9602 18000 9676
rect 17972 9574 18092 9602
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17788 9081 17816 9454
rect 17774 9072 17830 9081
rect 17774 9007 17830 9016
rect 18064 8786 18092 9574
rect 17788 8758 18092 8786
rect 17684 5840 17736 5846
rect 17684 5782 17736 5788
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17132 4140 17184 4146
rect 17132 4082 17184 4088
rect 17236 800 17264 4558
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17328 950 17356 4014
rect 17500 3460 17552 3466
rect 17500 3402 17552 3408
rect 17512 2922 17540 3402
rect 17788 3040 17816 8758
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17880 7818 17908 8434
rect 17958 8120 18014 8129
rect 17958 8055 18014 8064
rect 17972 8022 18000 8055
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 18064 7886 18092 8570
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17880 7342 17908 7754
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17880 6730 17908 7278
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17880 5642 17908 6666
rect 17972 6186 18000 6666
rect 18064 6390 18092 7822
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 18064 5710 18092 6326
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 17958 4720 18014 4729
rect 17958 4655 18014 4664
rect 17972 4010 18000 4655
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17868 3052 17920 3058
rect 17788 3012 17868 3040
rect 17868 2994 17920 3000
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17420 1306 17448 2586
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17512 1970 17540 2382
rect 17500 1964 17552 1970
rect 17500 1906 17552 1912
rect 17420 1278 17540 1306
rect 17316 944 17368 950
rect 17316 886 17368 892
rect 17512 800 17540 1278
rect 17604 1154 17632 2926
rect 17972 2650 18000 2926
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 17592 1148 17644 1154
rect 17592 1090 17644 1096
rect 17788 800 17816 2450
rect 18064 800 18092 4490
rect 18156 4146 18184 12679
rect 18326 12679 18382 12688
rect 18236 12650 18288 12656
rect 18248 11812 18276 12650
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18432 12238 18460 12582
rect 18524 12306 18552 12582
rect 18512 12300 18564 12306
rect 18512 12242 18564 12248
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18616 11914 18644 22066
rect 18800 20942 18828 22510
rect 18880 22228 18932 22234
rect 18880 22170 18932 22176
rect 18892 21962 18920 22170
rect 19168 22094 19196 26206
rect 19444 23730 19472 26206
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19444 23526 19472 23666
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19076 22066 19196 22094
rect 18880 21956 18932 21962
rect 18880 21898 18932 21904
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18800 20346 18828 20878
rect 18972 20800 19024 20806
rect 18972 20742 19024 20748
rect 18984 20534 19012 20742
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 18800 20330 18920 20346
rect 18800 20324 18932 20330
rect 18800 20318 18880 20324
rect 18880 20266 18932 20272
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18800 18970 18828 20198
rect 18892 19718 18920 20266
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18788 18964 18840 18970
rect 18788 18906 18840 18912
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18708 17746 18736 17818
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18708 16726 18736 17478
rect 18800 17202 18828 17682
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18788 17196 18840 17202
rect 18788 17138 18840 17144
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18696 16720 18748 16726
rect 18800 16697 18828 16730
rect 18696 16662 18748 16668
rect 18786 16688 18842 16697
rect 18786 16623 18842 16632
rect 18892 16590 18920 17274
rect 18880 16584 18932 16590
rect 18880 16526 18932 16532
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18708 15094 18736 16050
rect 18696 15088 18748 15094
rect 18696 15030 18748 15036
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18708 14414 18736 14554
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18694 13832 18750 13841
rect 18694 13767 18750 13776
rect 18524 11886 18644 11914
rect 18328 11824 18380 11830
rect 18248 11784 18328 11812
rect 18248 11150 18276 11784
rect 18328 11766 18380 11772
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18234 9344 18290 9353
rect 18234 9279 18290 9288
rect 18248 6730 18276 9279
rect 18340 8838 18368 9522
rect 18432 8974 18460 10542
rect 18524 10538 18552 11886
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18524 10130 18552 10474
rect 18512 10124 18564 10130
rect 18512 10066 18564 10072
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18524 9042 18552 9318
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18420 8968 18472 8974
rect 18420 8910 18472 8916
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18432 8566 18460 8774
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 18432 7818 18460 8502
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18236 6724 18288 6730
rect 18236 6666 18288 6672
rect 18432 5710 18460 7754
rect 18524 7478 18552 7822
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 18616 6338 18644 10542
rect 18524 6310 18644 6338
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18524 5137 18552 6310
rect 18604 5160 18656 5166
rect 18510 5128 18566 5137
rect 18604 5102 18656 5108
rect 18510 5063 18566 5072
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18524 3534 18552 5063
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 18156 1222 18184 2926
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 18248 2106 18276 2314
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 18144 1216 18196 1222
rect 18144 1158 18196 1164
rect 18328 944 18380 950
rect 18328 886 18380 892
rect 18340 800 18368 886
rect 18616 800 18644 5102
rect 18708 3058 18736 13767
rect 18800 10266 18828 16390
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18892 15094 18920 15438
rect 18984 15162 19012 16118
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18880 15088 18932 15094
rect 18880 15030 18932 15036
rect 18892 14414 18920 15030
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18892 13462 18920 14350
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 19076 10198 19104 22066
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19616 21548 19668 21554
rect 19616 21490 19668 21496
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19168 19514 19196 20402
rect 19260 20262 19288 21422
rect 19628 21146 19656 21490
rect 19708 21344 19760 21350
rect 19706 21312 19708 21321
rect 19760 21312 19762 21321
rect 19706 21247 19762 21256
rect 19616 21140 19668 21146
rect 19616 21082 19668 21088
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19444 20602 19472 20878
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19248 20256 19300 20262
rect 19248 20198 19300 20204
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19156 19372 19208 19378
rect 19260 19360 19288 19654
rect 19208 19332 19288 19360
rect 19156 19314 19208 19320
rect 19352 19310 19380 19722
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19260 18086 19288 18566
rect 19352 18086 19380 18634
rect 19444 18272 19472 20538
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19890 19272 19946 19281
rect 19890 19207 19946 19216
rect 19904 19174 19932 19207
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19524 18284 19576 18290
rect 19444 18244 19524 18272
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19168 16266 19196 17274
rect 19352 17202 19380 18022
rect 19444 17678 19472 18244
rect 19524 18226 19576 18232
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19628 17678 19656 18158
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19260 16658 19288 17002
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19536 16726 19564 16934
rect 19524 16720 19576 16726
rect 19524 16662 19576 16668
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19524 16584 19576 16590
rect 19352 16544 19524 16572
rect 19168 16238 19288 16266
rect 19260 16182 19288 16238
rect 19248 16176 19300 16182
rect 19248 16118 19300 16124
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 19168 15570 19196 16050
rect 19352 15586 19380 16544
rect 19524 16526 19576 16532
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19260 15558 19380 15586
rect 19904 15570 19932 15846
rect 19892 15564 19944 15570
rect 19168 14822 19196 15506
rect 19260 15434 19288 15558
rect 19892 15506 19944 15512
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19260 15162 19288 15370
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19444 15026 19472 15302
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19996 15042 20024 30534
rect 20444 23520 20496 23526
rect 20444 23462 20496 23468
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 20074 21040 20130 21049
rect 20074 20975 20130 20984
rect 20088 20058 20116 20975
rect 20180 20942 20208 21286
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20168 20528 20220 20534
rect 20168 20470 20220 20476
rect 20180 20058 20208 20470
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 20088 19378 20116 19858
rect 20180 19378 20208 19994
rect 20272 19990 20300 21490
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 20168 18692 20220 18698
rect 20168 18634 20220 18640
rect 20180 18222 20208 18634
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 20272 18086 20300 19926
rect 20364 18834 20392 20198
rect 20352 18828 20404 18834
rect 20352 18770 20404 18776
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20364 17134 20392 18770
rect 20456 17610 20484 23462
rect 20548 22094 20576 37198
rect 20640 36242 20668 37606
rect 20720 37392 20772 37398
rect 20720 37334 20772 37340
rect 20732 36786 20760 37334
rect 20720 36780 20772 36786
rect 20720 36722 20772 36728
rect 20628 36236 20680 36242
rect 20628 36178 20680 36184
rect 20720 36236 20772 36242
rect 20720 36178 20772 36184
rect 20628 33448 20680 33454
rect 20628 33390 20680 33396
rect 20640 25702 20668 33390
rect 20628 25696 20680 25702
rect 20628 25638 20680 25644
rect 20732 22094 20760 36178
rect 20824 34649 20852 37674
rect 20916 37330 20944 38490
rect 20996 38480 21048 38486
rect 20996 38422 21048 38428
rect 21008 38010 21036 38422
rect 20996 38004 21048 38010
rect 20996 37946 21048 37952
rect 21088 37868 21140 37874
rect 21088 37810 21140 37816
rect 21100 37466 21128 37810
rect 21088 37460 21140 37466
rect 21088 37402 21140 37408
rect 21100 37330 21128 37402
rect 20904 37324 20956 37330
rect 20904 37266 20956 37272
rect 21088 37324 21140 37330
rect 21088 37266 21140 37272
rect 20996 36576 21048 36582
rect 20996 36518 21048 36524
rect 21008 35834 21036 36518
rect 20996 35828 21048 35834
rect 20996 35770 21048 35776
rect 21100 35766 21128 37266
rect 21180 36712 21232 36718
rect 21180 36654 21232 36660
rect 21088 35760 21140 35766
rect 21088 35702 21140 35708
rect 21088 35624 21140 35630
rect 21088 35566 21140 35572
rect 20810 34640 20866 34649
rect 20810 34575 20866 34584
rect 21100 34202 21128 35566
rect 21192 35086 21220 36654
rect 21180 35080 21232 35086
rect 21180 35022 21232 35028
rect 21088 34196 21140 34202
rect 21088 34138 21140 34144
rect 21100 33522 21128 34138
rect 21284 33522 21312 44882
rect 21468 41414 21496 45358
rect 21376 41386 21496 41414
rect 21376 37874 21404 41386
rect 21640 40044 21692 40050
rect 21640 39986 21692 39992
rect 21546 37904 21602 37913
rect 21364 37868 21416 37874
rect 21546 37839 21602 37848
rect 21364 37810 21416 37816
rect 21456 37800 21508 37806
rect 21456 37742 21508 37748
rect 21364 36576 21416 36582
rect 21364 36518 21416 36524
rect 21376 36310 21404 36518
rect 21468 36310 21496 37742
rect 21364 36304 21416 36310
rect 21364 36246 21416 36252
rect 21456 36304 21508 36310
rect 21456 36246 21508 36252
rect 21560 33998 21588 37839
rect 21456 33992 21508 33998
rect 21456 33934 21508 33940
rect 21548 33992 21600 33998
rect 21548 33934 21600 33940
rect 20904 33516 20956 33522
rect 20904 33458 20956 33464
rect 21088 33516 21140 33522
rect 21088 33458 21140 33464
rect 21272 33516 21324 33522
rect 21272 33458 21324 33464
rect 20916 22982 20944 33458
rect 21284 31754 21312 33458
rect 21192 31726 21312 31754
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 21192 22094 21220 31726
rect 21468 29578 21496 33934
rect 21560 31278 21588 33934
rect 21548 31272 21600 31278
rect 21548 31214 21600 31220
rect 21456 29572 21508 29578
rect 21456 29514 21508 29520
rect 21652 28626 21680 39986
rect 21732 38208 21784 38214
rect 21732 38150 21784 38156
rect 21744 32910 21772 38150
rect 21824 36848 21876 36854
rect 21824 36790 21876 36796
rect 21836 36650 21864 36790
rect 21824 36644 21876 36650
rect 21824 36586 21876 36592
rect 21928 34066 21956 60182
rect 22020 60178 22048 60998
rect 22008 60172 22060 60178
rect 22008 60114 22060 60120
rect 22112 59634 22140 61270
rect 22204 61198 22232 63200
rect 23020 61260 23072 61266
rect 23020 61202 23072 61208
rect 22192 61192 22244 61198
rect 22192 61134 22244 61140
rect 22192 60784 22244 60790
rect 22190 60752 22192 60761
rect 22244 60752 22246 60761
rect 22190 60687 22246 60696
rect 22192 60648 22244 60654
rect 22192 60590 22244 60596
rect 22100 59628 22152 59634
rect 22100 59570 22152 59576
rect 22100 54596 22152 54602
rect 22100 54538 22152 54544
rect 21916 34060 21968 34066
rect 21916 34002 21968 34008
rect 21824 33992 21876 33998
rect 21824 33934 21876 33940
rect 21732 32904 21784 32910
rect 21732 32846 21784 32852
rect 21836 31822 21864 33934
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 21824 31816 21876 31822
rect 21824 31758 21876 31764
rect 22020 30666 22048 32370
rect 22008 30660 22060 30666
rect 22008 30602 22060 30608
rect 21916 30592 21968 30598
rect 21916 30534 21968 30540
rect 21640 28620 21692 28626
rect 21640 28562 21692 28568
rect 21652 27062 21680 28562
rect 21640 27056 21692 27062
rect 21640 26998 21692 27004
rect 20548 22066 20668 22094
rect 20732 22066 20944 22094
rect 21192 22066 21312 22094
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20444 17604 20496 17610
rect 20444 17546 20496 17552
rect 20548 17202 20576 20266
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20364 16590 20392 16934
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20364 16250 20392 16526
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20548 16182 20576 17138
rect 20536 16176 20588 16182
rect 20536 16118 20588 16124
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 19432 15020 19484 15026
rect 19996 15014 20116 15042
rect 20272 15026 20300 15438
rect 20456 15162 20484 15438
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 19432 14962 19484 14968
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19168 14618 19196 14758
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19352 13394 19380 14350
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19352 12986 19380 13330
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19156 12708 19208 12714
rect 19156 12650 19208 12656
rect 19168 11354 19196 12650
rect 19248 12436 19300 12442
rect 19444 12434 19472 13806
rect 19524 13796 19576 13802
rect 19524 13738 19576 13744
rect 19708 13796 19760 13802
rect 19708 13738 19760 13744
rect 19536 13705 19564 13738
rect 19616 13728 19668 13734
rect 19522 13696 19578 13705
rect 19616 13670 19668 13676
rect 19522 13631 19578 13640
rect 19628 13326 19656 13670
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 19720 13258 19748 13738
rect 19708 13252 19760 13258
rect 19708 13194 19760 13200
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19248 12378 19300 12384
rect 19352 12406 19472 12434
rect 19156 11348 19208 11354
rect 19156 11290 19208 11296
rect 19260 11218 19288 12378
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19352 10810 19380 12406
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19616 11688 19668 11694
rect 19522 11656 19578 11665
rect 19616 11630 19668 11636
rect 19522 11591 19578 11600
rect 19536 11558 19564 11591
rect 19524 11552 19576 11558
rect 19430 11520 19486 11529
rect 19524 11494 19576 11500
rect 19430 11455 19486 11464
rect 19444 11286 19472 11455
rect 19432 11280 19484 11286
rect 19432 11222 19484 11228
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19444 10674 19472 11086
rect 19628 11014 19656 11630
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19904 11082 19932 11494
rect 19996 11370 20024 14894
rect 20088 12306 20116 15014
rect 20260 15020 20312 15026
rect 20260 14962 20312 14968
rect 20272 14414 20300 14962
rect 20640 14793 20668 22066
rect 20916 21622 20944 22066
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 20904 21616 20956 21622
rect 20904 21558 20956 21564
rect 20812 21548 20864 21554
rect 20812 21490 20864 21496
rect 20720 21344 20772 21350
rect 20720 21286 20772 21292
rect 20732 18766 20760 21286
rect 20824 19854 20852 21490
rect 21100 21146 21128 21966
rect 21088 21140 21140 21146
rect 21088 21082 21140 21088
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20916 20398 20944 20878
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20916 18970 20944 19314
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20732 18086 20760 18226
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 21008 17762 21036 20334
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21192 19281 21220 19314
rect 21178 19272 21234 19281
rect 21178 19207 21234 19216
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21100 18970 21128 19110
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 21192 18630 21220 19110
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 20916 17734 21036 17762
rect 20916 17678 20944 17734
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 20812 16652 20864 16658
rect 20812 16594 20864 16600
rect 20626 14784 20682 14793
rect 20626 14719 20682 14728
rect 20640 14498 20668 14719
rect 20456 14470 20668 14498
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20180 14113 20208 14214
rect 20166 14104 20222 14113
rect 20166 14039 20222 14048
rect 20180 13938 20208 14039
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20272 13462 20300 14350
rect 20352 14000 20404 14006
rect 20352 13942 20404 13948
rect 20260 13456 20312 13462
rect 20260 13398 20312 13404
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20272 12374 20300 13262
rect 20260 12368 20312 12374
rect 20260 12310 20312 12316
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20272 11694 20300 12174
rect 20364 11762 20392 13942
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20088 11558 20116 11630
rect 20076 11552 20128 11558
rect 20364 11529 20392 11698
rect 20076 11494 20128 11500
rect 20350 11520 20406 11529
rect 20350 11455 20406 11464
rect 20456 11370 20484 14470
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20640 13802 20668 14214
rect 20824 14074 20852 16594
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20628 13796 20680 13802
rect 20628 13738 20680 13744
rect 20824 13394 20852 14010
rect 20916 13852 20944 17614
rect 21008 17338 21036 17614
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 21100 16590 21128 17478
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 20996 13864 21048 13870
rect 20916 13824 20996 13852
rect 20916 13462 20944 13824
rect 20996 13806 21048 13812
rect 21284 13818 21312 22066
rect 21364 22092 21416 22098
rect 21928 22094 21956 30534
rect 22112 22094 22140 54538
rect 22204 52018 22232 60590
rect 22284 60512 22336 60518
rect 22284 60454 22336 60460
rect 22296 60110 22324 60454
rect 23032 60110 23060 61202
rect 23216 60110 23244 63294
rect 23662 63200 23718 64000
rect 24398 63200 24454 64000
rect 25134 63200 25190 64000
rect 25870 63322 25926 64000
rect 25870 63294 26280 63322
rect 25870 63200 25926 63294
rect 23480 61668 23532 61674
rect 23480 61610 23532 61616
rect 23296 60240 23348 60246
rect 23296 60182 23348 60188
rect 22284 60104 22336 60110
rect 22284 60046 22336 60052
rect 22560 60104 22612 60110
rect 22560 60046 22612 60052
rect 22836 60104 22888 60110
rect 22836 60046 22888 60052
rect 23020 60104 23072 60110
rect 23020 60046 23072 60052
rect 23204 60104 23256 60110
rect 23204 60046 23256 60052
rect 22296 59974 22324 60046
rect 22284 59968 22336 59974
rect 22284 59910 22336 59916
rect 22572 59498 22600 60046
rect 22848 59702 22876 60046
rect 22836 59696 22888 59702
rect 22836 59638 22888 59644
rect 23308 59634 23336 60182
rect 23388 59968 23440 59974
rect 23388 59910 23440 59916
rect 23400 59634 23428 59910
rect 23492 59634 23520 61610
rect 23676 61198 23704 63200
rect 23664 61192 23716 61198
rect 23664 61134 23716 61140
rect 24412 60790 24440 63200
rect 25148 61198 25176 63200
rect 26252 61198 26280 63294
rect 26606 63200 26662 64000
rect 27342 63322 27398 64000
rect 27342 63294 27568 63322
rect 27342 63200 27398 63294
rect 26620 61198 26648 63200
rect 26884 61328 26936 61334
rect 26884 61270 26936 61276
rect 25136 61192 25188 61198
rect 25136 61134 25188 61140
rect 26240 61192 26292 61198
rect 26240 61134 26292 61140
rect 26608 61192 26660 61198
rect 26608 61134 26660 61140
rect 24768 61124 24820 61130
rect 24768 61066 24820 61072
rect 24676 61056 24728 61062
rect 24676 60998 24728 61004
rect 24688 60790 24716 60998
rect 24400 60784 24452 60790
rect 24400 60726 24452 60732
rect 24676 60784 24728 60790
rect 24676 60726 24728 60732
rect 23664 60716 23716 60722
rect 23664 60658 23716 60664
rect 23676 59974 23704 60658
rect 24400 60512 24452 60518
rect 24400 60454 24452 60460
rect 24676 60512 24728 60518
rect 24676 60454 24728 60460
rect 23664 59968 23716 59974
rect 23664 59910 23716 59916
rect 23756 59968 23808 59974
rect 23756 59910 23808 59916
rect 23296 59628 23348 59634
rect 23296 59570 23348 59576
rect 23388 59628 23440 59634
rect 23388 59570 23440 59576
rect 23480 59628 23532 59634
rect 23480 59570 23532 59576
rect 23572 59628 23624 59634
rect 23572 59570 23624 59576
rect 23400 59498 23428 59570
rect 22560 59492 22612 59498
rect 22560 59434 22612 59440
rect 23388 59492 23440 59498
rect 23388 59434 23440 59440
rect 22468 59424 22520 59430
rect 22468 59366 22520 59372
rect 22928 59424 22980 59430
rect 22928 59366 22980 59372
rect 22480 56846 22508 59366
rect 22468 56840 22520 56846
rect 22468 56782 22520 56788
rect 22192 52012 22244 52018
rect 22192 51954 22244 51960
rect 22836 52012 22888 52018
rect 22836 51954 22888 51960
rect 22192 42628 22244 42634
rect 22192 42570 22244 42576
rect 22204 37398 22232 42570
rect 22560 42084 22612 42090
rect 22560 42026 22612 42032
rect 22284 39840 22336 39846
rect 22284 39782 22336 39788
rect 22296 38962 22324 39782
rect 22284 38956 22336 38962
rect 22284 38898 22336 38904
rect 22468 38888 22520 38894
rect 22468 38830 22520 38836
rect 22480 38729 22508 38830
rect 22466 38720 22522 38729
rect 22466 38655 22522 38664
rect 22192 37392 22244 37398
rect 22192 37334 22244 37340
rect 22572 36174 22600 42026
rect 22652 39568 22704 39574
rect 22652 39510 22704 39516
rect 22284 36168 22336 36174
rect 22284 36110 22336 36116
rect 22560 36168 22612 36174
rect 22560 36110 22612 36116
rect 22192 36032 22244 36038
rect 22192 35974 22244 35980
rect 22204 30258 22232 35974
rect 22296 35222 22324 36110
rect 22284 35216 22336 35222
rect 22284 35158 22336 35164
rect 22664 35018 22692 39510
rect 22848 37942 22876 51954
rect 22940 38350 22968 59366
rect 23584 59022 23612 59570
rect 23572 59016 23624 59022
rect 23572 58958 23624 58964
rect 23572 55956 23624 55962
rect 23572 55898 23624 55904
rect 23584 54670 23612 55898
rect 23572 54664 23624 54670
rect 23572 54606 23624 54612
rect 23584 53990 23612 54606
rect 23572 53984 23624 53990
rect 23572 53926 23624 53932
rect 23676 53106 23704 59910
rect 23664 53100 23716 53106
rect 23664 53042 23716 53048
rect 23664 42152 23716 42158
rect 23664 42094 23716 42100
rect 23110 38856 23166 38865
rect 23110 38791 23112 38800
rect 23164 38791 23166 38800
rect 23112 38762 23164 38768
rect 23112 38480 23164 38486
rect 23112 38422 23164 38428
rect 23388 38480 23440 38486
rect 23388 38422 23440 38428
rect 22928 38344 22980 38350
rect 22928 38286 22980 38292
rect 22836 37936 22888 37942
rect 22836 37878 22888 37884
rect 22848 37670 22876 37878
rect 23020 37868 23072 37874
rect 23020 37810 23072 37816
rect 23032 37777 23060 37810
rect 23018 37768 23074 37777
rect 23018 37703 23074 37712
rect 22836 37664 22888 37670
rect 22836 37606 22888 37612
rect 23124 36122 23152 38422
rect 23400 38350 23428 38422
rect 23388 38344 23440 38350
rect 23388 38286 23440 38292
rect 23204 38276 23256 38282
rect 23204 38218 23256 38224
rect 23216 36258 23244 38218
rect 23572 38208 23624 38214
rect 23572 38150 23624 38156
rect 23480 36576 23532 36582
rect 23480 36518 23532 36524
rect 23492 36378 23520 36518
rect 23480 36372 23532 36378
rect 23480 36314 23532 36320
rect 23216 36230 23520 36258
rect 23584 36242 23612 38150
rect 23296 36168 23348 36174
rect 23124 36094 23244 36122
rect 23296 36110 23348 36116
rect 23388 36168 23440 36174
rect 23388 36110 23440 36116
rect 22744 36032 22796 36038
rect 22744 35974 22796 35980
rect 22756 35290 22784 35974
rect 22744 35284 22796 35290
rect 22744 35226 22796 35232
rect 22652 35012 22704 35018
rect 22652 34954 22704 34960
rect 22928 34944 22980 34950
rect 22928 34886 22980 34892
rect 22376 34740 22428 34746
rect 22376 34682 22428 34688
rect 22388 33590 22416 34682
rect 22940 33998 22968 34886
rect 22928 33992 22980 33998
rect 22928 33934 22980 33940
rect 23112 33924 23164 33930
rect 23112 33866 23164 33872
rect 22376 33584 22428 33590
rect 22376 33526 22428 33532
rect 22284 33516 22336 33522
rect 22284 33458 22336 33464
rect 22296 33425 22324 33458
rect 22282 33416 22338 33425
rect 22282 33351 22338 33360
rect 22652 33312 22704 33318
rect 22652 33254 22704 33260
rect 22664 33046 22692 33254
rect 22652 33040 22704 33046
rect 22652 32982 22704 32988
rect 22560 32836 22612 32842
rect 22560 32778 22612 32784
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22204 29714 22232 30194
rect 22192 29708 22244 29714
rect 22192 29650 22244 29656
rect 22468 23044 22520 23050
rect 22468 22986 22520 22992
rect 21928 22066 22048 22094
rect 22112 22066 22232 22094
rect 21364 22034 21416 22040
rect 21376 21418 21404 22034
rect 21640 21684 21692 21690
rect 21640 21626 21692 21632
rect 21364 21412 21416 21418
rect 21364 21354 21416 21360
rect 21652 20942 21680 21626
rect 21824 21616 21876 21622
rect 21824 21558 21876 21564
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21376 19854 21404 20198
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21456 19780 21508 19786
rect 21456 19722 21508 19728
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 21376 18766 21404 19246
rect 21468 19009 21496 19722
rect 21652 19718 21680 20878
rect 21732 20324 21784 20330
rect 21732 20266 21784 20272
rect 21744 19990 21772 20266
rect 21732 19984 21784 19990
rect 21732 19926 21784 19932
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21640 19508 21692 19514
rect 21744 19496 21772 19790
rect 21692 19468 21772 19496
rect 21640 19450 21692 19456
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21454 19000 21510 19009
rect 21454 18935 21510 18944
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21560 18358 21588 19110
rect 21548 18352 21600 18358
rect 21548 18294 21600 18300
rect 21652 18290 21680 19450
rect 21836 19334 21864 21558
rect 21744 19306 21864 19334
rect 21640 18284 21692 18290
rect 21640 18226 21692 18232
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21284 13790 21404 13818
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 20812 13388 20864 13394
rect 20812 13330 20864 13336
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20732 12986 20760 13262
rect 20916 13258 20944 13398
rect 20996 13388 21048 13394
rect 20996 13330 21048 13336
rect 20904 13252 20956 13258
rect 20904 13194 20956 13200
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 21008 12918 21036 13330
rect 21284 13326 21312 13670
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 19996 11342 20300 11370
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19982 10976 20038 10985
rect 19574 10908 19882 10917
rect 19982 10911 20038 10920
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10792 20024 10911
rect 19720 10764 20024 10792
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 18972 9988 19024 9994
rect 18972 9930 19024 9936
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18892 9110 18920 9318
rect 18880 9104 18932 9110
rect 18880 9046 18932 9052
rect 18984 7002 19012 9930
rect 19076 9926 19104 10134
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 19168 8634 19196 10202
rect 19444 10130 19472 10610
rect 19720 10538 19748 10764
rect 19708 10532 19760 10538
rect 19708 10474 19760 10480
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 20166 9888 20222 9897
rect 19574 9820 19882 9829
rect 20166 9823 20222 9832
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19982 9752 20038 9761
rect 19982 9687 20038 9696
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19444 9042 19472 9454
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 19076 4622 19104 7890
rect 19260 6458 19288 8502
rect 19338 8256 19394 8265
rect 19338 8191 19394 8200
rect 19352 8090 19380 8191
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19444 7342 19472 8978
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19996 6866 20024 9687
rect 20074 9072 20130 9081
rect 20074 9007 20130 9016
rect 20088 8809 20116 9007
rect 20074 8800 20130 8809
rect 20074 8735 20130 8744
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 20088 7002 20116 7278
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 19432 6724 19484 6730
rect 19432 6666 19484 6672
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19338 6080 19394 6089
rect 19338 6015 19394 6024
rect 19352 5352 19380 6015
rect 19444 5642 19472 6666
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6458 20024 6802
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19892 5364 19944 5370
rect 19352 5324 19656 5352
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 19260 4554 19288 5170
rect 19536 4826 19564 5170
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19352 4622 19380 4762
rect 19628 4758 19656 5324
rect 19996 5352 20024 6258
rect 19944 5324 20024 5352
rect 19892 5306 19944 5312
rect 20076 5160 20128 5166
rect 20076 5102 20128 5108
rect 20088 4758 20116 5102
rect 19616 4752 19668 4758
rect 19616 4694 19668 4700
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19156 4548 19208 4554
rect 19156 4490 19208 4496
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18984 3942 19012 4082
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 19076 3194 19104 3538
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18880 2304 18932 2310
rect 18880 2246 18932 2252
rect 18892 800 18920 2246
rect 18984 1086 19012 2926
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 19076 2310 19104 2586
rect 19064 2304 19116 2310
rect 19064 2246 19116 2252
rect 18972 1080 19024 1086
rect 18972 1022 19024 1028
rect 19168 800 19196 4490
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19892 4208 19944 4214
rect 20180 4196 20208 9823
rect 20272 9024 20300 11342
rect 20364 11342 20484 11370
rect 20364 11200 20392 11342
rect 20364 11172 20484 11200
rect 20350 10840 20406 10849
rect 20350 10775 20406 10784
rect 20364 9466 20392 10775
rect 20456 9586 20484 11172
rect 20548 10849 20576 12242
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20534 10840 20590 10849
rect 20534 10775 20590 10784
rect 20536 10736 20588 10742
rect 20536 10678 20588 10684
rect 20548 10062 20576 10678
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20364 9438 20484 9466
rect 20272 8996 20392 9024
rect 20260 8900 20312 8906
rect 20260 8842 20312 8848
rect 20272 8634 20300 8842
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20364 7546 20392 8996
rect 20456 7954 20484 9438
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20640 7562 20668 12174
rect 20824 11286 20852 12650
rect 21008 12434 21036 12854
rect 20916 12406 21036 12434
rect 20916 12238 20944 12406
rect 21100 12238 21128 13126
rect 21180 12776 21232 12782
rect 21178 12744 21180 12753
rect 21232 12744 21234 12753
rect 21178 12679 21234 12688
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21088 11824 21140 11830
rect 21088 11766 21140 11772
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 9110 20760 10950
rect 20916 10674 20944 11630
rect 20994 11520 21050 11529
rect 20994 11455 21050 11464
rect 21008 11354 21036 11455
rect 21100 11354 21128 11766
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 20916 9994 20944 10610
rect 21088 10600 21140 10606
rect 21088 10542 21140 10548
rect 21100 10198 21128 10542
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 21100 9382 21128 9998
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20916 8566 20944 8774
rect 20904 8560 20956 8566
rect 20904 8502 20956 8508
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20548 7534 20668 7562
rect 20260 6928 20312 6934
rect 20260 6870 20312 6876
rect 20272 6390 20300 6870
rect 20260 6384 20312 6390
rect 20260 6326 20312 6332
rect 20272 5642 20300 6326
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 20364 5386 20392 7482
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 20272 5358 20392 5386
rect 20456 5370 20484 6666
rect 20444 5364 20496 5370
rect 20272 4622 20300 5358
rect 20444 5306 20496 5312
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20364 4554 20392 5238
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 20444 4480 20496 4486
rect 20442 4448 20444 4457
rect 20496 4448 20498 4457
rect 20442 4383 20498 4392
rect 19944 4168 20208 4196
rect 19892 4150 19944 4156
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19260 1018 19288 4014
rect 19720 3641 19748 4082
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 19706 3632 19762 3641
rect 19432 3596 19484 3602
rect 19706 3567 19708 3576
rect 19432 3538 19484 3544
rect 19760 3567 19762 3576
rect 19708 3538 19760 3544
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19352 3233 19380 3334
rect 19338 3224 19394 3233
rect 19338 3159 19394 3168
rect 19444 3058 19472 3538
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19444 1442 19472 2858
rect 19996 2650 20024 2994
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19444 1414 19748 1442
rect 19248 1012 19300 1018
rect 19248 954 19300 960
rect 19432 944 19484 950
rect 19432 886 19484 892
rect 19444 800 19472 886
rect 19720 800 19748 1414
rect 20088 1034 20116 3878
rect 20456 3194 20484 4082
rect 20548 3369 20576 7534
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20640 7002 20668 7346
rect 20628 6996 20680 7002
rect 20628 6938 20680 6944
rect 21100 6866 21128 9318
rect 21192 8634 21220 12679
rect 21376 11914 21404 13790
rect 21468 13734 21496 17070
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 21468 12782 21496 13670
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21376 11886 21496 11914
rect 21364 11824 21416 11830
rect 21364 11766 21416 11772
rect 21376 11665 21404 11766
rect 21362 11656 21418 11665
rect 21362 11591 21418 11600
rect 21468 10742 21496 11886
rect 21456 10736 21508 10742
rect 21456 10678 21508 10684
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21284 8430 21312 10134
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21468 9761 21496 9862
rect 21454 9752 21510 9761
rect 21454 9687 21510 9696
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21284 6866 21312 8366
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 21008 6118 21036 6394
rect 21088 6180 21140 6186
rect 21088 6122 21140 6128
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 21100 5642 21128 6122
rect 21088 5636 21140 5642
rect 21088 5578 21140 5584
rect 21284 5574 21312 6802
rect 21468 6662 21496 7142
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 20916 5030 20944 5102
rect 21008 5098 21036 5510
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 20996 5092 21048 5098
rect 20996 5034 21048 5040
rect 21088 5092 21140 5098
rect 21088 5034 21140 5040
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20640 4214 20668 4422
rect 20732 4214 20760 4966
rect 21100 4758 21128 5034
rect 21088 4752 21140 4758
rect 21088 4694 21140 4700
rect 21192 4570 21220 5102
rect 21284 4690 21312 5510
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21100 4542 21220 4570
rect 20628 4208 20680 4214
rect 20628 4150 20680 4156
rect 20720 4208 20772 4214
rect 20720 4150 20772 4156
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20534 3360 20590 3369
rect 20534 3295 20590 3304
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20364 3058 20392 3130
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20456 2514 20484 3130
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 20548 2446 20576 3295
rect 20732 2961 20760 3878
rect 20718 2952 20774 2961
rect 20718 2887 20774 2896
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 19996 1006 20116 1034
rect 19996 800 20024 1006
rect 20272 800 20300 2382
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 20536 1148 20588 1154
rect 20536 1090 20588 1096
rect 20548 800 20576 1090
rect 20732 950 20760 2314
rect 20812 1012 20864 1018
rect 20812 954 20864 960
rect 20720 944 20772 950
rect 20720 886 20772 892
rect 20824 800 20852 954
rect 21100 800 21128 4542
rect 21180 4480 21232 4486
rect 21180 4422 21232 4428
rect 21192 4282 21220 4422
rect 21180 4276 21232 4282
rect 21180 4218 21232 4224
rect 21284 3058 21312 4626
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 21180 2508 21232 2514
rect 21284 2496 21312 2994
rect 21560 2774 21588 17546
rect 21744 15434 21772 19306
rect 21916 19236 21968 19242
rect 21916 19178 21968 19184
rect 21928 18222 21956 19178
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 21916 17196 21968 17202
rect 21916 17138 21968 17144
rect 21928 16454 21956 17138
rect 21916 16448 21968 16454
rect 21916 16390 21968 16396
rect 21928 16114 21956 16390
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 21928 15910 21956 16050
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 21732 15428 21784 15434
rect 21732 15370 21784 15376
rect 21638 13696 21694 13705
rect 21638 13631 21694 13640
rect 21652 12889 21680 13631
rect 21638 12880 21694 12889
rect 21638 12815 21640 12824
rect 21692 12815 21694 12824
rect 21640 12786 21692 12792
rect 21640 11144 21692 11150
rect 21638 11112 21640 11121
rect 21692 11112 21694 11121
rect 21638 11047 21694 11056
rect 21640 9920 21692 9926
rect 21744 9897 21772 15370
rect 21824 14884 21876 14890
rect 21824 14826 21876 14832
rect 21836 14618 21864 14826
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21822 12472 21878 12481
rect 21822 12407 21824 12416
rect 21876 12407 21878 12416
rect 21824 12378 21876 12384
rect 21824 10532 21876 10538
rect 21824 10474 21876 10480
rect 21836 10198 21864 10474
rect 21824 10192 21876 10198
rect 21824 10134 21876 10140
rect 21640 9862 21692 9868
rect 21730 9888 21786 9897
rect 21652 9654 21680 9862
rect 21730 9823 21786 9832
rect 21640 9648 21692 9654
rect 21640 9590 21692 9596
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21640 9104 21692 9110
rect 21640 9046 21692 9052
rect 21652 4865 21680 9046
rect 21836 5234 21864 9522
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21638 4856 21694 4865
rect 21638 4791 21694 4800
rect 21928 3534 21956 13126
rect 22020 11150 22048 22066
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 22112 19718 22140 20402
rect 22204 19825 22232 22066
rect 22480 20602 22508 22986
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22190 19816 22246 19825
rect 22190 19751 22246 19760
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22112 19378 22140 19654
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22112 18290 22140 19314
rect 22480 19310 22508 20538
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22284 17060 22336 17066
rect 22284 17002 22336 17008
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22008 9716 22060 9722
rect 22008 9658 22060 9664
rect 22020 9217 22048 9658
rect 22006 9208 22062 9217
rect 22006 9143 22062 9152
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22020 7313 22048 7346
rect 22006 7304 22062 7313
rect 22006 7239 22062 7248
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 21376 2746 21588 2774
rect 21376 2582 21404 2746
rect 21364 2576 21416 2582
rect 21364 2518 21416 2524
rect 21232 2468 21312 2496
rect 21180 2450 21232 2456
rect 21640 2100 21692 2106
rect 21640 2042 21692 2048
rect 21364 1216 21416 1222
rect 21364 1158 21416 1164
rect 21376 800 21404 1158
rect 21652 800 21680 2042
rect 21916 1080 21968 1086
rect 21916 1022 21968 1028
rect 21928 800 21956 1022
rect 22020 1018 22048 3402
rect 22112 2446 22140 14350
rect 22190 12880 22246 12889
rect 22190 12815 22192 12824
rect 22244 12815 22246 12824
rect 22192 12786 22244 12792
rect 22204 12442 22232 12786
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 22296 10810 22324 17002
rect 22572 15162 22600 32778
rect 23020 32224 23072 32230
rect 23020 32166 23072 32172
rect 23032 31822 23060 32166
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 23020 31272 23072 31278
rect 23020 31214 23072 31220
rect 22836 30728 22888 30734
rect 22836 30670 22888 30676
rect 22848 30394 22876 30670
rect 23032 30666 23060 31214
rect 23020 30660 23072 30666
rect 23020 30602 23072 30608
rect 22836 30388 22888 30394
rect 22836 30330 22888 30336
rect 23124 30138 23152 33866
rect 23216 30734 23244 36094
rect 23308 32502 23336 36110
rect 23400 35630 23428 36110
rect 23492 35894 23520 36230
rect 23572 36236 23624 36242
rect 23572 36178 23624 36184
rect 23676 36122 23704 42094
rect 23584 36106 23704 36122
rect 23572 36100 23704 36106
rect 23624 36094 23704 36100
rect 23572 36042 23624 36048
rect 23492 35866 23612 35894
rect 23388 35624 23440 35630
rect 23388 35566 23440 35572
rect 23584 35290 23612 35866
rect 23572 35284 23624 35290
rect 23572 35226 23624 35232
rect 23388 34536 23440 34542
rect 23388 34478 23440 34484
rect 23400 33318 23428 34478
rect 23584 34202 23612 35226
rect 23572 34196 23624 34202
rect 23572 34138 23624 34144
rect 23480 34128 23532 34134
rect 23480 34070 23532 34076
rect 23492 33522 23520 34070
rect 23480 33516 23532 33522
rect 23480 33458 23532 33464
rect 23388 33312 23440 33318
rect 23388 33254 23440 33260
rect 23296 32496 23348 32502
rect 23296 32438 23348 32444
rect 23400 31822 23428 33254
rect 23388 31816 23440 31822
rect 23308 31764 23388 31770
rect 23308 31758 23440 31764
rect 23308 31742 23428 31758
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23216 30598 23244 30670
rect 23204 30592 23256 30598
rect 23204 30534 23256 30540
rect 23204 30252 23256 30258
rect 23204 30194 23256 30200
rect 23032 30110 23152 30138
rect 22836 30048 22888 30054
rect 22836 29990 22888 29996
rect 22650 29880 22706 29889
rect 22650 29815 22706 29824
rect 22664 29646 22692 29815
rect 22848 29646 22876 29990
rect 22652 29640 22704 29646
rect 22652 29582 22704 29588
rect 22836 29640 22888 29646
rect 22836 29582 22888 29588
rect 22928 29504 22980 29510
rect 22928 29446 22980 29452
rect 22744 21956 22796 21962
rect 22744 21898 22796 21904
rect 22652 18828 22704 18834
rect 22652 18770 22704 18776
rect 22664 18086 22692 18770
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 22652 17264 22704 17270
rect 22652 17206 22704 17212
rect 22664 16794 22692 17206
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22664 15026 22692 16526
rect 22756 16425 22784 21898
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22848 18737 22876 20198
rect 22834 18728 22890 18737
rect 22834 18663 22890 18672
rect 22848 16697 22876 18663
rect 22834 16688 22890 16697
rect 22834 16623 22890 16632
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22742 16416 22798 16425
rect 22742 16351 22798 16360
rect 22848 15638 22876 16526
rect 22940 16250 22968 29446
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 23032 15892 23060 30110
rect 23112 30048 23164 30054
rect 23112 29990 23164 29996
rect 23124 29714 23152 29990
rect 23216 29714 23244 30194
rect 23112 29708 23164 29714
rect 23112 29650 23164 29656
rect 23204 29708 23256 29714
rect 23204 29650 23256 29656
rect 23204 26920 23256 26926
rect 23204 26862 23256 26868
rect 23216 20262 23244 26862
rect 23308 21962 23336 31742
rect 23492 31210 23520 33458
rect 23572 33380 23624 33386
rect 23572 33322 23624 33328
rect 23584 32910 23612 33322
rect 23572 32904 23624 32910
rect 23572 32846 23624 32852
rect 23584 31770 23612 32846
rect 23584 31742 23704 31770
rect 23572 31680 23624 31686
rect 23572 31622 23624 31628
rect 23480 31204 23532 31210
rect 23480 31146 23532 31152
rect 23388 30592 23440 30598
rect 23388 30534 23440 30540
rect 23400 30258 23428 30534
rect 23584 30258 23612 31622
rect 23388 30252 23440 30258
rect 23388 30194 23440 30200
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23676 30054 23704 31742
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23768 28914 23796 59910
rect 24124 55820 24176 55826
rect 24124 55762 24176 55768
rect 23938 55312 23994 55321
rect 23938 55247 23940 55256
rect 23992 55247 23994 55256
rect 24032 55276 24084 55282
rect 23940 55218 23992 55224
rect 24032 55218 24084 55224
rect 23848 52896 23900 52902
rect 23848 52838 23900 52844
rect 23860 37874 23888 52838
rect 24044 45554 24072 55218
rect 23952 45526 24072 45554
rect 23848 37868 23900 37874
rect 23848 37810 23900 37816
rect 23952 36786 23980 45526
rect 24136 37806 24164 55762
rect 24308 55412 24360 55418
rect 24308 55354 24360 55360
rect 24320 54670 24348 55354
rect 24412 55282 24440 60454
rect 24492 59424 24544 59430
rect 24492 59366 24544 59372
rect 24400 55276 24452 55282
rect 24400 55218 24452 55224
rect 24308 54664 24360 54670
rect 24308 54606 24360 54612
rect 24216 53984 24268 53990
rect 24216 53926 24268 53932
rect 24228 51814 24256 53926
rect 24216 51808 24268 51814
rect 24216 51750 24268 51756
rect 24124 37800 24176 37806
rect 24124 37742 24176 37748
rect 24032 37664 24084 37670
rect 24032 37606 24084 37612
rect 23940 36780 23992 36786
rect 23940 36722 23992 36728
rect 23848 36712 23900 36718
rect 23848 36654 23900 36660
rect 23860 36378 23888 36654
rect 23848 36372 23900 36378
rect 23848 36314 23900 36320
rect 23848 34196 23900 34202
rect 23848 34138 23900 34144
rect 23860 30258 23888 34138
rect 23848 30252 23900 30258
rect 23848 30194 23900 30200
rect 23860 30138 23888 30194
rect 23860 30110 23980 30138
rect 23848 30048 23900 30054
rect 23848 29990 23900 29996
rect 23400 28886 23796 28914
rect 23400 26382 23428 28886
rect 23754 27704 23810 27713
rect 23754 27639 23810 27648
rect 23480 26988 23532 26994
rect 23480 26930 23532 26936
rect 23664 26988 23716 26994
rect 23664 26930 23716 26936
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23296 21956 23348 21962
rect 23296 21898 23348 21904
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 23204 20256 23256 20262
rect 23204 20198 23256 20204
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23216 19825 23244 19858
rect 23202 19816 23258 19825
rect 23202 19751 23258 19760
rect 23202 19000 23258 19009
rect 23202 18935 23258 18944
rect 23216 18766 23244 18935
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 23308 17746 23336 21286
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23400 20058 23428 20334
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23400 19378 23428 19994
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23296 17740 23348 17746
rect 23296 17682 23348 17688
rect 23492 16266 23520 26930
rect 23676 26586 23704 26930
rect 23664 26580 23716 26586
rect 23664 26522 23716 26528
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23584 23662 23612 26318
rect 23572 23656 23624 23662
rect 23572 23598 23624 23604
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 23584 21146 23612 21490
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23664 17808 23716 17814
rect 23664 17750 23716 17756
rect 23676 16998 23704 17750
rect 23664 16992 23716 16998
rect 23664 16934 23716 16940
rect 23296 16244 23348 16250
rect 23492 16238 23704 16266
rect 23296 16186 23348 16192
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 22940 15864 23060 15892
rect 23112 15904 23164 15910
rect 22836 15632 22888 15638
rect 22836 15574 22888 15580
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22756 15026 22784 15098
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 22744 15020 22796 15026
rect 22744 14962 22796 14968
rect 22940 14414 22968 15864
rect 23112 15846 23164 15852
rect 23020 15428 23072 15434
rect 23020 15370 23072 15376
rect 22928 14408 22980 14414
rect 22466 14376 22522 14385
rect 22928 14350 22980 14356
rect 22466 14311 22522 14320
rect 22560 14340 22612 14346
rect 22374 14104 22430 14113
rect 22480 14074 22508 14311
rect 22560 14282 22612 14288
rect 22652 14340 22704 14346
rect 22652 14282 22704 14288
rect 22572 14074 22600 14282
rect 22374 14039 22376 14048
rect 22428 14039 22430 14048
rect 22468 14068 22520 14074
rect 22376 14010 22428 14016
rect 22468 14010 22520 14016
rect 22560 14068 22612 14074
rect 22560 14010 22612 14016
rect 22388 13530 22416 14010
rect 22376 13524 22428 13530
rect 22376 13466 22428 13472
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22480 9926 22508 14010
rect 22558 11520 22614 11529
rect 22558 11455 22614 11464
rect 22468 9920 22520 9926
rect 22468 9862 22520 9868
rect 22374 7032 22430 7041
rect 22374 6967 22430 6976
rect 22388 6730 22416 6967
rect 22376 6724 22428 6730
rect 22376 6666 22428 6672
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 22204 6361 22232 6598
rect 22190 6352 22246 6361
rect 22190 6287 22246 6296
rect 22374 5536 22430 5545
rect 22374 5471 22430 5480
rect 22388 4622 22416 5471
rect 22572 5234 22600 11455
rect 22664 8906 22692 14282
rect 23032 12850 23060 15370
rect 23124 14414 23152 15846
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23216 14346 23244 16050
rect 23308 14822 23336 16186
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 23388 15632 23440 15638
rect 23388 15574 23440 15580
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 23308 13977 23336 14758
rect 23400 14414 23428 15574
rect 23480 15020 23532 15026
rect 23480 14962 23532 14968
rect 23492 14482 23520 14962
rect 23480 14476 23532 14482
rect 23480 14418 23532 14424
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23294 13968 23350 13977
rect 23294 13903 23350 13912
rect 23386 13696 23442 13705
rect 23386 13631 23442 13640
rect 23400 12986 23428 13631
rect 23584 13258 23612 16118
rect 23676 15910 23704 16238
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23676 14482 23704 15098
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23572 13252 23624 13258
rect 23572 13194 23624 13200
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 23018 12744 23074 12753
rect 23018 12679 23074 12688
rect 22836 9716 22888 9722
rect 22836 9658 22888 9664
rect 22652 8900 22704 8906
rect 22652 8842 22704 8848
rect 22664 7834 22692 8842
rect 22664 7806 22784 7834
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22664 6730 22692 7686
rect 22652 6724 22704 6730
rect 22652 6666 22704 6672
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22468 5160 22520 5166
rect 22468 5102 22520 5108
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22008 1012 22060 1018
rect 22008 954 22060 960
rect 22192 944 22244 950
rect 22192 886 22244 892
rect 22204 800 22232 886
rect 22480 800 22508 5102
rect 22756 4865 22784 7806
rect 22742 4856 22798 4865
rect 22742 4791 22798 4800
rect 22560 4548 22612 4554
rect 22560 4490 22612 4496
rect 22744 4548 22796 4554
rect 22744 4490 22796 4496
rect 22572 4185 22600 4490
rect 22558 4176 22614 4185
rect 22558 4111 22614 4120
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 22664 4049 22692 4082
rect 22650 4040 22706 4049
rect 22650 3975 22706 3984
rect 22650 3632 22706 3641
rect 22650 3567 22706 3576
rect 22664 3534 22692 3567
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 22756 800 22784 4490
rect 22848 3058 22876 9658
rect 22926 8392 22982 8401
rect 22926 8327 22982 8336
rect 22940 8294 22968 8327
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 22940 7750 22968 7822
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22940 7478 22968 7686
rect 22928 7472 22980 7478
rect 22928 7414 22980 7420
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 23032 1970 23060 12679
rect 23202 11656 23258 11665
rect 23202 11591 23258 11600
rect 23112 7744 23164 7750
rect 23112 7686 23164 7692
rect 23124 6458 23152 7686
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23216 6390 23244 11591
rect 23294 10432 23350 10441
rect 23294 10367 23350 10376
rect 23308 8566 23336 10367
rect 23400 9586 23428 12922
rect 23584 10130 23612 13194
rect 23768 10674 23796 27639
rect 23860 27062 23888 29990
rect 23848 27056 23900 27062
rect 23848 26998 23900 27004
rect 23952 26314 23980 30110
rect 23940 26308 23992 26314
rect 23940 26250 23992 26256
rect 24044 22094 24072 37606
rect 24124 36780 24176 36786
rect 24124 36722 24176 36728
rect 24136 34649 24164 36722
rect 24122 34640 24178 34649
rect 24122 34575 24178 34584
rect 24228 31754 24256 51750
rect 24320 42770 24348 54606
rect 24400 53508 24452 53514
rect 24400 53450 24452 53456
rect 24412 53106 24440 53450
rect 24400 53100 24452 53106
rect 24400 53042 24452 53048
rect 24308 42764 24360 42770
rect 24308 42706 24360 42712
rect 24320 36174 24348 42706
rect 24412 42634 24440 53042
rect 24400 42628 24452 42634
rect 24400 42570 24452 42576
rect 24400 37800 24452 37806
rect 24400 37742 24452 37748
rect 24308 36168 24360 36174
rect 24308 36110 24360 36116
rect 24412 35086 24440 37742
rect 24400 35080 24452 35086
rect 24400 35022 24452 35028
rect 24504 33998 24532 59366
rect 24584 55684 24636 55690
rect 24584 55626 24636 55632
rect 24596 40746 24624 55626
rect 24688 45554 24716 60454
rect 24780 55282 24808 61066
rect 25412 61056 25464 61062
rect 25412 60998 25464 61004
rect 24860 60512 24912 60518
rect 24860 60454 24912 60460
rect 24872 60178 24900 60454
rect 24860 60172 24912 60178
rect 24912 60132 24992 60160
rect 24860 60114 24912 60120
rect 24860 59492 24912 59498
rect 24860 59434 24912 59440
rect 24872 56982 24900 59434
rect 24860 56976 24912 56982
rect 24860 56918 24912 56924
rect 24964 55282 24992 60132
rect 24768 55276 24820 55282
rect 24768 55218 24820 55224
rect 24952 55276 25004 55282
rect 24952 55218 25004 55224
rect 25320 55276 25372 55282
rect 25320 55218 25372 55224
rect 24952 53644 25004 53650
rect 24952 53586 25004 53592
rect 24964 53242 24992 53586
rect 24952 53236 25004 53242
rect 24952 53178 25004 53184
rect 24964 52698 24992 53178
rect 24952 52692 25004 52698
rect 24952 52634 25004 52640
rect 24688 45526 24808 45554
rect 24596 40718 24716 40746
rect 24584 36576 24636 36582
rect 24584 36518 24636 36524
rect 24596 36174 24624 36518
rect 24584 36168 24636 36174
rect 24584 36110 24636 36116
rect 24492 33992 24544 33998
rect 24492 33934 24544 33940
rect 24228 31726 24532 31754
rect 24228 31346 24256 31726
rect 24308 31476 24360 31482
rect 24308 31418 24360 31424
rect 24216 31340 24268 31346
rect 24216 31282 24268 31288
rect 24124 31204 24176 31210
rect 24124 31146 24176 31152
rect 24216 31204 24268 31210
rect 24216 31146 24268 31152
rect 24136 26382 24164 31146
rect 24228 26994 24256 31146
rect 24320 29306 24348 31418
rect 24400 31340 24452 31346
rect 24400 31282 24452 31288
rect 24412 30938 24440 31282
rect 24400 30932 24452 30938
rect 24400 30874 24452 30880
rect 24504 29782 24532 31726
rect 24492 29776 24544 29782
rect 24492 29718 24544 29724
rect 24308 29300 24360 29306
rect 24308 29242 24360 29248
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24124 26376 24176 26382
rect 24124 26318 24176 26324
rect 24228 23118 24256 26930
rect 24216 23112 24268 23118
rect 24216 23054 24268 23060
rect 23952 22066 24072 22094
rect 24320 22094 24348 29242
rect 24504 29034 24532 29718
rect 24492 29028 24544 29034
rect 24492 28970 24544 28976
rect 24400 26988 24452 26994
rect 24400 26930 24452 26936
rect 24412 26790 24440 26930
rect 24400 26784 24452 26790
rect 24400 26726 24452 26732
rect 24688 22094 24716 40718
rect 24780 37942 24808 45526
rect 25332 38554 25360 55218
rect 25424 49094 25452 60998
rect 25688 55752 25740 55758
rect 25688 55694 25740 55700
rect 25700 55418 25728 55694
rect 25688 55412 25740 55418
rect 25688 55354 25740 55360
rect 25412 49088 25464 49094
rect 25412 49030 25464 49036
rect 25320 38548 25372 38554
rect 25320 38490 25372 38496
rect 24768 37936 24820 37942
rect 24768 37878 24820 37884
rect 25134 37904 25190 37913
rect 25332 37874 25360 38490
rect 25134 37839 25136 37848
rect 25188 37839 25190 37848
rect 25320 37868 25372 37874
rect 25136 37810 25188 37816
rect 25320 37810 25372 37816
rect 24952 36032 25004 36038
rect 24952 35974 25004 35980
rect 24860 34672 24912 34678
rect 24860 34614 24912 34620
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 24780 32570 24808 33934
rect 24872 33658 24900 34614
rect 24964 34066 24992 35974
rect 25148 35834 25176 37810
rect 25228 36100 25280 36106
rect 25228 36042 25280 36048
rect 25240 35894 25268 36042
rect 25240 35866 25360 35894
rect 25136 35828 25188 35834
rect 25136 35770 25188 35776
rect 24952 34060 25004 34066
rect 24952 34002 25004 34008
rect 25044 33856 25096 33862
rect 25044 33798 25096 33804
rect 24860 33652 24912 33658
rect 24860 33594 24912 33600
rect 24952 33448 25004 33454
rect 24952 33390 25004 33396
rect 24768 32564 24820 32570
rect 24768 32506 24820 32512
rect 24860 32428 24912 32434
rect 24860 32370 24912 32376
rect 24872 31482 24900 32370
rect 24860 31476 24912 31482
rect 24860 31418 24912 31424
rect 24964 31210 24992 33390
rect 25056 32434 25084 33798
rect 25044 32428 25096 32434
rect 25044 32370 25096 32376
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 24952 31204 25004 31210
rect 24952 31146 25004 31152
rect 25240 27713 25268 32302
rect 25226 27704 25282 27713
rect 25226 27639 25282 27648
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 24780 23662 24808 24346
rect 24768 23656 24820 23662
rect 24768 23598 24820 23604
rect 24320 22066 24440 22094
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23860 20466 23888 20878
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23952 17678 23980 22066
rect 24030 20904 24086 20913
rect 24030 20839 24086 20848
rect 24044 19922 24072 20839
rect 24032 19916 24084 19922
rect 24032 19858 24084 19864
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 24228 17746 24256 18226
rect 24308 18148 24360 18154
rect 24308 18090 24360 18096
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24136 16250 24164 17138
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 23848 16108 23900 16114
rect 24228 16096 24256 17682
rect 24320 17610 24348 18090
rect 24308 17604 24360 17610
rect 24308 17546 24360 17552
rect 23900 16068 24256 16096
rect 23848 16050 23900 16056
rect 23848 15972 23900 15978
rect 23848 15914 23900 15920
rect 23860 15502 23888 15914
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23952 13938 23980 15846
rect 24032 15632 24084 15638
rect 24032 15574 24084 15580
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 24044 13462 24072 15574
rect 24124 15564 24176 15570
rect 24124 15506 24176 15512
rect 24136 15026 24164 15506
rect 24228 15434 24256 16068
rect 24308 16108 24360 16114
rect 24308 16050 24360 16056
rect 24320 15638 24348 16050
rect 24308 15632 24360 15638
rect 24308 15574 24360 15580
rect 24216 15428 24268 15434
rect 24216 15370 24268 15376
rect 24228 15026 24256 15370
rect 24308 15088 24360 15094
rect 24308 15030 24360 15036
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24032 13456 24084 13462
rect 24032 13398 24084 13404
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 23940 11280 23992 11286
rect 23940 11222 23992 11228
rect 23756 10668 23808 10674
rect 23756 10610 23808 10616
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23478 8936 23534 8945
rect 23478 8871 23480 8880
rect 23532 8871 23534 8880
rect 23480 8842 23532 8848
rect 23584 8786 23612 10066
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23676 8906 23704 9318
rect 23664 8900 23716 8906
rect 23664 8842 23716 8848
rect 23492 8758 23612 8786
rect 23386 8664 23442 8673
rect 23386 8599 23388 8608
rect 23440 8599 23442 8608
rect 23388 8570 23440 8576
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 23492 7954 23520 8758
rect 23676 8650 23704 8842
rect 23584 8622 23704 8650
rect 23584 8498 23612 8622
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23664 8492 23716 8498
rect 23664 8434 23716 8440
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23388 6996 23440 7002
rect 23308 6956 23388 6984
rect 23204 6384 23256 6390
rect 23204 6326 23256 6332
rect 23308 4146 23336 6956
rect 23388 6938 23440 6944
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23400 5001 23428 6258
rect 23492 5030 23520 7890
rect 23572 7472 23624 7478
rect 23572 7414 23624 7420
rect 23584 5914 23612 7414
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23572 5160 23624 5166
rect 23572 5102 23624 5108
rect 23480 5024 23532 5030
rect 23386 4992 23442 5001
rect 23480 4966 23532 4972
rect 23386 4927 23442 4936
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23492 4146 23520 4422
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23112 4072 23164 4078
rect 23112 4014 23164 4020
rect 23124 2774 23152 4014
rect 23308 3534 23336 4082
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23204 3460 23256 3466
rect 23204 3402 23256 3408
rect 23216 3194 23244 3402
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23124 2746 23336 2774
rect 23204 2372 23256 2378
rect 23204 2314 23256 2320
rect 23020 1964 23072 1970
rect 23020 1906 23072 1912
rect 23216 1018 23244 2314
rect 23020 1012 23072 1018
rect 23020 954 23072 960
rect 23204 1012 23256 1018
rect 23204 954 23256 960
rect 23032 800 23060 954
rect 23308 800 23336 2746
rect 23400 950 23428 2926
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23492 2106 23520 2382
rect 23480 2100 23532 2106
rect 23480 2042 23532 2048
rect 23388 944 23440 950
rect 23388 886 23440 892
rect 23584 800 23612 5102
rect 23676 4729 23704 8434
rect 23662 4720 23718 4729
rect 23662 4655 23718 4664
rect 23768 4570 23796 10610
rect 23848 10600 23900 10606
rect 23848 10542 23900 10548
rect 23860 8362 23888 10542
rect 23952 9058 23980 11222
rect 24044 9450 24072 11834
rect 24136 10606 24164 14962
rect 24228 14414 24256 14962
rect 24320 14822 24348 15030
rect 24308 14816 24360 14822
rect 24308 14758 24360 14764
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24124 10464 24176 10470
rect 24124 10406 24176 10412
rect 24032 9444 24084 9450
rect 24032 9386 24084 9392
rect 23952 9030 24072 9058
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 23848 8356 23900 8362
rect 23848 8298 23900 8304
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 23860 5710 23888 6598
rect 23952 5914 23980 8910
rect 24044 8838 24072 9030
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 24044 8566 24072 8774
rect 24032 8560 24084 8566
rect 24032 8502 24084 8508
rect 24044 6254 24072 8502
rect 24136 7818 24164 10406
rect 24228 9654 24256 13874
rect 24306 12336 24362 12345
rect 24306 12271 24362 12280
rect 24320 10538 24348 12271
rect 24412 11778 24440 22066
rect 24596 22066 24716 22094
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24504 19174 24532 19790
rect 24492 19168 24544 19174
rect 24492 19110 24544 19116
rect 24596 18578 24624 22066
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 24964 20534 24992 20742
rect 24952 20528 25004 20534
rect 24952 20470 25004 20476
rect 25136 20528 25188 20534
rect 25136 20470 25188 20476
rect 25148 20262 25176 20470
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 24872 19922 24900 20198
rect 25148 20058 25176 20198
rect 24952 20052 25004 20058
rect 24952 19994 25004 20000
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 24768 19780 24820 19786
rect 24768 19722 24820 19728
rect 24780 19514 24808 19722
rect 24768 19508 24820 19514
rect 24768 19450 24820 19456
rect 24674 19272 24730 19281
rect 24674 19207 24730 19216
rect 24688 18902 24716 19207
rect 24676 18896 24728 18902
rect 24676 18838 24728 18844
rect 24964 18698 24992 19994
rect 25136 19712 25188 19718
rect 25136 19654 25188 19660
rect 25148 19378 25176 19654
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 25228 19168 25280 19174
rect 25228 19110 25280 19116
rect 25240 18698 25268 19110
rect 24952 18692 25004 18698
rect 24952 18634 25004 18640
rect 25228 18692 25280 18698
rect 25228 18634 25280 18640
rect 24860 18624 24912 18630
rect 24596 18572 24860 18578
rect 24596 18566 24912 18572
rect 24596 18550 24900 18566
rect 24492 18148 24544 18154
rect 24492 18090 24544 18096
rect 24504 17882 24532 18090
rect 24780 17921 24808 18550
rect 25136 18148 25188 18154
rect 25136 18090 25188 18096
rect 24766 17912 24822 17921
rect 24492 17876 24544 17882
rect 24766 17847 24822 17856
rect 24952 17876 25004 17882
rect 24492 17818 24544 17824
rect 24952 17818 25004 17824
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24688 17270 24716 17478
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24872 17202 24900 17478
rect 24964 17338 24992 17818
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 24952 17332 25004 17338
rect 24952 17274 25004 17280
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24492 16448 24544 16454
rect 24492 16390 24544 16396
rect 24504 11898 24532 16390
rect 24596 15502 24624 16526
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24688 15910 24716 16186
rect 24676 15904 24728 15910
rect 24676 15846 24728 15852
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24596 13530 24624 15438
rect 24688 14890 24716 15438
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24676 14340 24728 14346
rect 24676 14282 24728 14288
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24596 12918 24624 13466
rect 24688 13394 24716 14282
rect 24780 13938 24808 17070
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 24780 13841 24808 13874
rect 24766 13832 24822 13841
rect 24766 13767 24822 13776
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24872 13326 24900 17138
rect 24952 15360 25004 15366
rect 24952 15302 25004 15308
rect 24964 15094 24992 15302
rect 24952 15088 25004 15094
rect 24952 15030 25004 15036
rect 24950 14512 25006 14521
rect 24950 14447 25006 14456
rect 24964 14414 24992 14447
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 25056 14056 25084 17546
rect 25148 16114 25176 18090
rect 25240 17542 25268 18634
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25240 17338 25268 17478
rect 25228 17332 25280 17338
rect 25228 17274 25280 17280
rect 25136 16108 25188 16114
rect 25136 16050 25188 16056
rect 25240 15314 25268 17274
rect 25332 16969 25360 35866
rect 25964 30388 26016 30394
rect 25964 30330 26016 30336
rect 25412 29708 25464 29714
rect 25412 29650 25464 29656
rect 25424 19310 25452 29650
rect 25976 28422 26004 30330
rect 25964 28416 26016 28422
rect 25964 28358 26016 28364
rect 26896 26994 26924 61270
rect 27344 61056 27396 61062
rect 27344 60998 27396 61004
rect 27356 50454 27384 60998
rect 27540 60722 27568 63294
rect 28078 63200 28134 64000
rect 28814 63322 28870 64000
rect 29550 63322 29606 64000
rect 30286 63322 30342 64000
rect 28814 63294 29040 63322
rect 28814 63200 28870 63294
rect 28092 61198 28120 63200
rect 28908 61600 28960 61606
rect 28908 61542 28960 61548
rect 28080 61192 28132 61198
rect 28080 61134 28132 61140
rect 28172 61124 28224 61130
rect 28172 61066 28224 61072
rect 27528 60716 27580 60722
rect 27528 60658 27580 60664
rect 28184 60110 28212 61066
rect 28448 61056 28500 61062
rect 28448 60998 28500 61004
rect 28172 60104 28224 60110
rect 28172 60046 28224 60052
rect 28356 59628 28408 59634
rect 28356 59570 28408 59576
rect 27344 50448 27396 50454
rect 27344 50390 27396 50396
rect 26976 38412 27028 38418
rect 26976 38354 27028 38360
rect 26988 35894 27016 38354
rect 28264 37800 28316 37806
rect 28264 37742 28316 37748
rect 26988 35866 27108 35894
rect 26976 35080 27028 35086
rect 26976 35022 27028 35028
rect 26884 26988 26936 26994
rect 26884 26930 26936 26936
rect 26884 25900 26936 25906
rect 26884 25842 26936 25848
rect 25596 24200 25648 24206
rect 25596 24142 25648 24148
rect 25608 23186 25636 24142
rect 25596 23180 25648 23186
rect 25596 23122 25648 23128
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25688 21072 25740 21078
rect 25688 21014 25740 21020
rect 25778 21040 25834 21049
rect 25596 20936 25648 20942
rect 25596 20878 25648 20884
rect 25608 20602 25636 20878
rect 25700 20754 25728 21014
rect 25778 20975 25834 20984
rect 25792 20942 25820 20975
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25700 20726 25820 20754
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25504 20392 25556 20398
rect 25504 20334 25556 20340
rect 25516 19922 25544 20334
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25412 17536 25464 17542
rect 25412 17478 25464 17484
rect 25424 17270 25452 17478
rect 25412 17264 25464 17270
rect 25412 17206 25464 17212
rect 25318 16960 25374 16969
rect 25318 16895 25374 16904
rect 25410 16416 25466 16425
rect 25410 16351 25466 16360
rect 25148 15286 25268 15314
rect 25148 15162 25176 15286
rect 25226 15192 25282 15201
rect 25136 15156 25188 15162
rect 25226 15127 25282 15136
rect 25136 15098 25188 15104
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 24964 14028 25084 14056
rect 24964 13938 24992 14028
rect 25042 13968 25098 13977
rect 24952 13932 25004 13938
rect 25042 13903 25044 13912
rect 24952 13874 25004 13880
rect 25096 13903 25098 13912
rect 25044 13874 25096 13880
rect 25148 13802 25176 14962
rect 25240 13938 25268 15127
rect 25320 14544 25372 14550
rect 25318 14512 25320 14521
rect 25372 14512 25374 14521
rect 25318 14447 25374 14456
rect 25320 14272 25372 14278
rect 25318 14240 25320 14249
rect 25372 14240 25374 14249
rect 25318 14175 25374 14184
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25136 13796 25188 13802
rect 25136 13738 25188 13744
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24584 12912 24636 12918
rect 24584 12854 24636 12860
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24412 11750 24624 11778
rect 24400 11620 24452 11626
rect 24400 11562 24452 11568
rect 24412 11082 24440 11562
rect 24400 11076 24452 11082
rect 24400 11018 24452 11024
rect 24308 10532 24360 10538
rect 24308 10474 24360 10480
rect 24216 9648 24268 9654
rect 24216 9590 24268 9596
rect 24308 8492 24360 8498
rect 24308 8434 24360 8440
rect 24214 8120 24270 8129
rect 24214 8055 24270 8064
rect 24124 7812 24176 7818
rect 24124 7754 24176 7760
rect 24032 6248 24084 6254
rect 24032 6190 24084 6196
rect 23940 5908 23992 5914
rect 23940 5850 23992 5856
rect 23940 5772 23992 5778
rect 23940 5714 23992 5720
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 23848 5024 23900 5030
rect 23848 4966 23900 4972
rect 23860 4690 23888 4966
rect 23848 4684 23900 4690
rect 23848 4626 23900 4632
rect 23676 4542 23796 4570
rect 23952 4554 23980 5714
rect 24124 5636 24176 5642
rect 24124 5578 24176 5584
rect 23940 4548 23992 4554
rect 23676 3505 23704 4542
rect 23940 4490 23992 4496
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23768 3738 23796 4422
rect 23756 3732 23808 3738
rect 23756 3674 23808 3680
rect 23848 3528 23900 3534
rect 23662 3496 23718 3505
rect 23848 3470 23900 3476
rect 23662 3431 23718 3440
rect 23662 3224 23718 3233
rect 23662 3159 23664 3168
rect 23716 3159 23718 3168
rect 23664 3130 23716 3136
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 23676 2038 23704 2382
rect 23664 2032 23716 2038
rect 23664 1974 23716 1980
rect 23860 800 23888 3470
rect 23952 2990 23980 4490
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 24044 3126 24072 3334
rect 24032 3120 24084 3126
rect 24032 3062 24084 3068
rect 23940 2984 23992 2990
rect 23940 2926 23992 2932
rect 24136 2825 24164 5578
rect 24228 5234 24256 8055
rect 24320 7954 24348 8434
rect 24308 7948 24360 7954
rect 24308 7890 24360 7896
rect 24412 7546 24440 11018
rect 24492 10532 24544 10538
rect 24492 10474 24544 10480
rect 24504 10266 24532 10474
rect 24596 10470 24624 11750
rect 24688 11082 24716 12174
rect 24780 12170 24808 12718
rect 24872 12374 24900 13262
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24860 12368 24912 12374
rect 24860 12310 24912 12316
rect 24768 12164 24820 12170
rect 24768 12106 24820 12112
rect 24858 12064 24914 12073
rect 24858 11999 24914 12008
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24780 11286 24808 11834
rect 24768 11280 24820 11286
rect 24768 11222 24820 11228
rect 24676 11076 24728 11082
rect 24676 11018 24728 11024
rect 24584 10464 24636 10470
rect 24584 10406 24636 10412
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 24688 10180 24716 11018
rect 24872 10198 24900 11999
rect 24964 11694 24992 13126
rect 25424 12434 25452 16351
rect 25516 15026 25544 19858
rect 25792 19854 25820 20726
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 25608 19417 25636 19450
rect 25594 19408 25650 19417
rect 25792 19378 25820 19790
rect 25594 19343 25596 19352
rect 25648 19343 25650 19352
rect 25780 19372 25832 19378
rect 25596 19314 25648 19320
rect 25780 19314 25832 19320
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25792 18970 25820 19110
rect 25780 18964 25832 18970
rect 25780 18906 25832 18912
rect 25688 18760 25740 18766
rect 25688 18702 25740 18708
rect 25700 18426 25728 18702
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25688 18420 25740 18426
rect 25688 18362 25740 18368
rect 25608 18290 25636 18362
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25608 17746 25636 18226
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 25596 16176 25648 16182
rect 25596 16118 25648 16124
rect 25504 15020 25556 15026
rect 25504 14962 25556 14968
rect 25504 14884 25556 14890
rect 25504 14826 25556 14832
rect 25516 14414 25544 14826
rect 25504 14408 25556 14414
rect 25504 14350 25556 14356
rect 25504 14272 25556 14278
rect 25504 14214 25556 14220
rect 25516 13938 25544 14214
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25056 12406 25452 12434
rect 24952 11688 25004 11694
rect 24952 11630 25004 11636
rect 24964 11286 24992 11630
rect 24952 11280 25004 11286
rect 24952 11222 25004 11228
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 24768 10192 24820 10198
rect 24688 10152 24768 10180
rect 24768 10134 24820 10140
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24492 8492 24544 8498
rect 24492 8434 24544 8440
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24412 7002 24440 7482
rect 24504 7002 24532 8434
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 24492 6996 24544 7002
rect 24492 6938 24544 6944
rect 24412 6322 24440 6938
rect 24400 6316 24452 6322
rect 24400 6258 24452 6264
rect 24308 6248 24360 6254
rect 24308 6190 24360 6196
rect 24320 5574 24348 6190
rect 24504 5846 24532 6938
rect 24596 6390 24624 9522
rect 24872 9382 24900 9998
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24964 9042 24992 10542
rect 25056 10441 25084 12406
rect 25320 12164 25372 12170
rect 25320 12106 25372 12112
rect 25136 12096 25188 12102
rect 25136 12038 25188 12044
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25148 11150 25176 12038
rect 25240 11762 25268 12038
rect 25332 11898 25360 12106
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25228 11756 25280 11762
rect 25228 11698 25280 11704
rect 25424 11642 25452 11834
rect 25240 11614 25452 11642
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 25136 10464 25188 10470
rect 25042 10432 25098 10441
rect 25136 10406 25188 10412
rect 25042 10367 25098 10376
rect 25056 10130 25084 10367
rect 25148 10130 25176 10406
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 25056 8974 25084 9318
rect 25136 9104 25188 9110
rect 25136 9046 25188 9052
rect 25148 8974 25176 9046
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24964 8430 24992 8774
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24766 7848 24822 7857
rect 24766 7783 24822 7792
rect 24780 7750 24808 7783
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24860 7540 24912 7546
rect 24860 7482 24912 7488
rect 24584 6384 24636 6390
rect 24584 6326 24636 6332
rect 24872 6202 24900 7482
rect 24688 6174 24900 6202
rect 24688 6118 24716 6174
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24492 5840 24544 5846
rect 24492 5782 24544 5788
rect 24308 5568 24360 5574
rect 24308 5510 24360 5516
rect 24216 5228 24268 5234
rect 24216 5170 24268 5176
rect 24964 4690 24992 8366
rect 25056 8242 25084 8910
rect 25056 8214 25176 8242
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 25056 7954 25084 8026
rect 25044 7948 25096 7954
rect 25044 7890 25096 7896
rect 25056 7274 25084 7890
rect 25148 7546 25176 8214
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25044 7268 25096 7274
rect 25044 7210 25096 7216
rect 25136 7268 25188 7274
rect 25136 7210 25188 7216
rect 25148 6662 25176 7210
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25056 6390 25084 6598
rect 25148 6458 25176 6598
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 25044 6384 25096 6390
rect 25044 6326 25096 6332
rect 25148 5370 25176 6394
rect 25240 6390 25268 11614
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 25332 8634 25360 11154
rect 25504 11008 25556 11014
rect 25504 10950 25556 10956
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25424 10062 25452 10406
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 25516 9926 25544 10950
rect 25504 9920 25556 9926
rect 25504 9862 25556 9868
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 25412 9512 25464 9518
rect 25412 9454 25464 9460
rect 25424 8906 25452 9454
rect 25516 9110 25544 9590
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 25412 8900 25464 8906
rect 25412 8842 25464 8848
rect 25320 8628 25372 8634
rect 25320 8570 25372 8576
rect 25424 7274 25452 8842
rect 25516 7478 25544 9046
rect 25608 8129 25636 16118
rect 25688 16040 25740 16046
rect 25688 15982 25740 15988
rect 25700 15502 25728 15982
rect 25688 15496 25740 15502
rect 25688 15438 25740 15444
rect 25778 15056 25834 15065
rect 25778 14991 25780 15000
rect 25832 14991 25834 15000
rect 25780 14962 25832 14968
rect 25780 14884 25832 14890
rect 25884 14872 25912 23054
rect 25964 21548 26016 21554
rect 25964 21490 26016 21496
rect 25976 20505 26004 21490
rect 26424 21412 26476 21418
rect 26424 21354 26476 21360
rect 26146 21312 26202 21321
rect 26146 21247 26202 21256
rect 26160 21146 26188 21247
rect 26148 21140 26200 21146
rect 26148 21082 26200 21088
rect 26436 21010 26464 21354
rect 26790 21040 26846 21049
rect 26424 21004 26476 21010
rect 26790 20975 26846 20984
rect 26424 20946 26476 20952
rect 26804 20942 26832 20975
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26792 20800 26844 20806
rect 26792 20742 26844 20748
rect 26804 20534 26832 20742
rect 26792 20528 26844 20534
rect 25962 20496 26018 20505
rect 26792 20470 26844 20476
rect 25962 20431 26018 20440
rect 26516 20392 26568 20398
rect 26516 20334 26568 20340
rect 26146 20088 26202 20097
rect 26146 20023 26148 20032
rect 26200 20023 26202 20032
rect 26148 19994 26200 20000
rect 26160 19378 26188 19994
rect 26528 19446 26556 20334
rect 26516 19440 26568 19446
rect 26516 19382 26568 19388
rect 25964 19372 26016 19378
rect 25964 19314 26016 19320
rect 26148 19372 26200 19378
rect 26148 19314 26200 19320
rect 25976 18154 26004 19314
rect 26528 18834 26556 19382
rect 26516 18828 26568 18834
rect 26516 18770 26568 18776
rect 26148 18216 26200 18222
rect 26148 18158 26200 18164
rect 25964 18148 26016 18154
rect 25964 18090 26016 18096
rect 26056 17264 26108 17270
rect 26056 17206 26108 17212
rect 26068 16969 26096 17206
rect 26054 16960 26110 16969
rect 26054 16895 26110 16904
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 26068 16114 26096 16458
rect 26160 16454 26188 18158
rect 26528 16590 26556 18770
rect 26896 17218 26924 25842
rect 26804 17190 26924 17218
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26608 16584 26660 16590
rect 26608 16526 26660 16532
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26620 16250 26648 16526
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 26608 15972 26660 15978
rect 26608 15914 26660 15920
rect 26332 15088 26384 15094
rect 26332 15030 26384 15036
rect 25832 14844 25912 14872
rect 25780 14826 25832 14832
rect 26056 14816 26108 14822
rect 26056 14758 26108 14764
rect 25964 14544 26016 14550
rect 25962 14512 25964 14521
rect 26016 14512 26018 14521
rect 25962 14447 26018 14456
rect 25688 14408 25740 14414
rect 25688 14350 25740 14356
rect 25964 14408 26016 14414
rect 25964 14350 26016 14356
rect 25700 11898 25728 14350
rect 25976 14074 26004 14350
rect 25964 14068 26016 14074
rect 25964 14010 26016 14016
rect 25976 13938 26004 14010
rect 25964 13932 26016 13938
rect 25964 13874 26016 13880
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25780 13728 25832 13734
rect 25780 13670 25832 13676
rect 25792 12918 25820 13670
rect 25780 12912 25832 12918
rect 25780 12854 25832 12860
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 25700 11665 25728 11698
rect 25686 11656 25742 11665
rect 25686 11591 25742 11600
rect 25700 11558 25728 11591
rect 25688 11552 25740 11558
rect 25688 11494 25740 11500
rect 25688 11348 25740 11354
rect 25688 11290 25740 11296
rect 25594 8120 25650 8129
rect 25700 8090 25728 11290
rect 25780 10600 25832 10606
rect 25780 10542 25832 10548
rect 25792 9518 25820 10542
rect 25780 9512 25832 9518
rect 25780 9454 25832 9460
rect 25792 8974 25820 9454
rect 25884 9217 25912 13806
rect 26068 13734 26096 14758
rect 26146 14104 26202 14113
rect 26146 14039 26148 14048
rect 26200 14039 26202 14048
rect 26148 14010 26200 14016
rect 26148 13864 26200 13870
rect 26148 13806 26200 13812
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 26160 12850 26188 13806
rect 26344 13394 26372 15030
rect 26332 13388 26384 13394
rect 26332 13330 26384 13336
rect 26238 12880 26294 12889
rect 26148 12844 26200 12850
rect 26238 12815 26294 12824
rect 26148 12786 26200 12792
rect 26252 12424 26280 12815
rect 26160 12396 26280 12424
rect 25964 12232 26016 12238
rect 25964 12174 26016 12180
rect 25976 9654 26004 12174
rect 26056 12096 26108 12102
rect 26056 12038 26108 12044
rect 26068 11830 26096 12038
rect 26160 11898 26188 12396
rect 26240 12300 26292 12306
rect 26240 12242 26292 12248
rect 26148 11892 26200 11898
rect 26148 11834 26200 11840
rect 26056 11824 26108 11830
rect 26056 11766 26108 11772
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 26068 11014 26096 11630
rect 26056 11008 26108 11014
rect 26056 10950 26108 10956
rect 26054 10432 26110 10441
rect 26054 10367 26110 10376
rect 26068 10062 26096 10367
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 26148 10056 26200 10062
rect 26148 9998 26200 10004
rect 26054 9752 26110 9761
rect 26054 9687 26110 9696
rect 26068 9654 26096 9687
rect 25964 9648 26016 9654
rect 25964 9590 26016 9596
rect 26056 9648 26108 9654
rect 26056 9590 26108 9596
rect 26056 9512 26108 9518
rect 26056 9454 26108 9460
rect 25870 9208 25926 9217
rect 25870 9143 25926 9152
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 25780 8968 25832 8974
rect 25778 8936 25780 8945
rect 25832 8936 25834 8945
rect 25778 8871 25834 8880
rect 25976 8634 26004 9114
rect 26068 9042 26096 9454
rect 26160 9353 26188 9998
rect 26252 9382 26280 12242
rect 26240 9376 26292 9382
rect 26146 9344 26202 9353
rect 26344 9353 26372 13330
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 26436 11354 26464 12582
rect 26514 12472 26570 12481
rect 26514 12407 26570 12416
rect 26528 12374 26556 12407
rect 26516 12368 26568 12374
rect 26516 12310 26568 12316
rect 26516 12096 26568 12102
rect 26514 12064 26516 12073
rect 26568 12064 26570 12073
rect 26514 11999 26570 12008
rect 26528 11898 26556 11999
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26424 11348 26476 11354
rect 26424 11290 26476 11296
rect 26516 10056 26568 10062
rect 26516 9998 26568 10004
rect 26528 9761 26556 9998
rect 26514 9752 26570 9761
rect 26514 9687 26570 9696
rect 26240 9318 26292 9324
rect 26330 9344 26386 9353
rect 26146 9279 26202 9288
rect 26330 9279 26386 9288
rect 26332 9104 26384 9110
rect 26332 9046 26384 9052
rect 26056 9036 26108 9042
rect 26056 8978 26108 8984
rect 26240 8900 26292 8906
rect 26240 8842 26292 8848
rect 26252 8786 26280 8842
rect 26068 8758 26280 8786
rect 25964 8628 26016 8634
rect 25964 8570 26016 8576
rect 26068 8498 26096 8758
rect 26344 8673 26372 9046
rect 26620 8974 26648 15914
rect 26700 15496 26752 15502
rect 26700 15438 26752 15444
rect 26712 15162 26740 15438
rect 26700 15156 26752 15162
rect 26700 15098 26752 15104
rect 26698 14784 26754 14793
rect 26698 14719 26754 14728
rect 26712 14618 26740 14719
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26700 12164 26752 12170
rect 26700 12106 26752 12112
rect 26712 9586 26740 12106
rect 26804 11762 26832 17190
rect 26884 12844 26936 12850
rect 26884 12786 26936 12792
rect 26896 12102 26924 12786
rect 26884 12096 26936 12102
rect 26884 12038 26936 12044
rect 26792 11756 26844 11762
rect 26792 11698 26844 11704
rect 26804 11218 26832 11698
rect 26792 11212 26844 11218
rect 26792 11154 26844 11160
rect 26700 9580 26752 9586
rect 26700 9522 26752 9528
rect 26608 8968 26660 8974
rect 26608 8910 26660 8916
rect 26712 8838 26740 9522
rect 26804 9518 26832 11154
rect 26896 9926 26924 12038
rect 26988 11286 27016 35022
rect 27080 29646 27108 35866
rect 27344 29844 27396 29850
rect 27344 29786 27396 29792
rect 27068 29640 27120 29646
rect 27068 29582 27120 29588
rect 27068 27056 27120 27062
rect 27068 26998 27120 27004
rect 27080 19334 27108 26998
rect 27080 19306 27200 19334
rect 27068 17672 27120 17678
rect 27066 17640 27068 17649
rect 27120 17640 27122 17649
rect 27066 17575 27122 17584
rect 27172 17542 27200 19306
rect 27252 18692 27304 18698
rect 27252 18634 27304 18640
rect 27264 18426 27292 18634
rect 27252 18420 27304 18426
rect 27252 18362 27304 18368
rect 27356 17678 27384 29786
rect 28276 28490 28304 37742
rect 28368 37262 28396 59570
rect 28460 40730 28488 60998
rect 28920 60042 28948 61542
rect 29012 60722 29040 63294
rect 29550 63294 29868 63322
rect 30208 63306 30342 63322
rect 31022 63322 31078 64000
rect 29550 63200 29606 63294
rect 29840 61198 29868 63294
rect 30196 63300 30342 63306
rect 30248 63294 30342 63300
rect 30196 63242 30248 63248
rect 30286 63200 30342 63294
rect 30472 63300 30524 63306
rect 30472 63242 30524 63248
rect 31022 63294 31248 63322
rect 30288 61736 30340 61742
rect 30288 61678 30340 61684
rect 29828 61192 29880 61198
rect 29828 61134 29880 61140
rect 29920 61056 29972 61062
rect 29920 60998 29972 61004
rect 29000 60716 29052 60722
rect 29000 60658 29052 60664
rect 29000 60512 29052 60518
rect 29828 60512 29880 60518
rect 29052 60460 29132 60466
rect 29000 60454 29132 60460
rect 29828 60454 29880 60460
rect 29012 60438 29132 60454
rect 29104 60330 29132 60438
rect 29104 60302 29224 60330
rect 29196 60178 29224 60302
rect 29092 60172 29144 60178
rect 29092 60114 29144 60120
rect 29184 60172 29236 60178
rect 29184 60114 29236 60120
rect 28908 60036 28960 60042
rect 28908 59978 28960 59984
rect 29104 59974 29132 60114
rect 28632 59968 28684 59974
rect 28632 59910 28684 59916
rect 28724 59968 28776 59974
rect 29092 59968 29144 59974
rect 28724 59910 28776 59916
rect 29090 59936 29092 59945
rect 29144 59936 29146 59945
rect 28644 59634 28672 59910
rect 28632 59628 28684 59634
rect 28632 59570 28684 59576
rect 28736 54738 28764 59910
rect 29090 59871 29146 59880
rect 29460 59696 29512 59702
rect 29512 59644 29684 59650
rect 29460 59638 29684 59644
rect 29472 59622 29684 59638
rect 29840 59634 29868 60454
rect 29656 59566 29684 59622
rect 29736 59628 29788 59634
rect 29736 59570 29788 59576
rect 29828 59628 29880 59634
rect 29828 59570 29880 59576
rect 29644 59560 29696 59566
rect 29748 59537 29776 59570
rect 29644 59502 29696 59508
rect 29734 59528 29790 59537
rect 29734 59463 29790 59472
rect 29748 59430 29776 59463
rect 29736 59424 29788 59430
rect 29736 59366 29788 59372
rect 29736 55684 29788 55690
rect 29736 55626 29788 55632
rect 28724 54732 28776 54738
rect 28724 54674 28776 54680
rect 29552 50380 29604 50386
rect 29552 50322 29604 50328
rect 28448 40724 28500 40730
rect 28448 40666 28500 40672
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 28264 28484 28316 28490
rect 28264 28426 28316 28432
rect 27896 26988 27948 26994
rect 27896 26930 27948 26936
rect 27804 20936 27856 20942
rect 27804 20878 27856 20884
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27526 19816 27582 19825
rect 27526 19751 27528 19760
rect 27580 19751 27582 19760
rect 27528 19722 27580 19728
rect 27436 19712 27488 19718
rect 27436 19654 27488 19660
rect 27448 19428 27476 19654
rect 27528 19440 27580 19446
rect 27448 19400 27528 19428
rect 27528 19382 27580 19388
rect 27436 19236 27488 19242
rect 27436 19178 27488 19184
rect 27448 18816 27476 19178
rect 27528 18828 27580 18834
rect 27448 18788 27528 18816
rect 27344 17672 27396 17678
rect 27344 17614 27396 17620
rect 27160 17536 27212 17542
rect 27160 17478 27212 17484
rect 27344 17536 27396 17542
rect 27344 17478 27396 17484
rect 27160 16516 27212 16522
rect 27160 16458 27212 16464
rect 27172 16250 27200 16458
rect 27252 16448 27304 16454
rect 27252 16390 27304 16396
rect 27160 16244 27212 16250
rect 27160 16186 27212 16192
rect 27264 16046 27292 16390
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 27068 12436 27120 12442
rect 27068 12378 27120 12384
rect 26976 11280 27028 11286
rect 26976 11222 27028 11228
rect 26884 9920 26936 9926
rect 26884 9862 26936 9868
rect 26792 9512 26844 9518
rect 26792 9454 26844 9460
rect 26790 9344 26846 9353
rect 26790 9279 26846 9288
rect 26700 8832 26752 8838
rect 26804 8809 26832 9279
rect 26988 9042 27016 11222
rect 27080 10674 27108 12378
rect 27160 11144 27212 11150
rect 27160 11086 27212 11092
rect 27068 10668 27120 10674
rect 27068 10610 27120 10616
rect 27172 10538 27200 11086
rect 27160 10532 27212 10538
rect 27160 10474 27212 10480
rect 27158 10432 27214 10441
rect 27158 10367 27214 10376
rect 27068 9920 27120 9926
rect 27068 9862 27120 9868
rect 26976 9036 27028 9042
rect 26976 8978 27028 8984
rect 26700 8774 26752 8780
rect 26790 8800 26846 8809
rect 26790 8735 26846 8744
rect 26330 8664 26386 8673
rect 26330 8599 26386 8608
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 25594 8055 25650 8064
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25504 7472 25556 7478
rect 25504 7414 25556 7420
rect 25412 7268 25464 7274
rect 25412 7210 25464 7216
rect 25516 7206 25544 7414
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25780 6656 25832 6662
rect 25780 6598 25832 6604
rect 25228 6384 25280 6390
rect 25228 6326 25280 6332
rect 25792 5914 25820 6598
rect 25780 5908 25832 5914
rect 25780 5850 25832 5856
rect 25320 5704 25372 5710
rect 25320 5646 25372 5652
rect 25136 5364 25188 5370
rect 25136 5306 25188 5312
rect 25226 5264 25282 5273
rect 25226 5199 25282 5208
rect 24952 4684 25004 4690
rect 24952 4626 25004 4632
rect 24676 4616 24728 4622
rect 24676 4558 24728 4564
rect 24688 4282 24716 4558
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 25240 4146 25268 5199
rect 25228 4140 25280 4146
rect 25228 4082 25280 4088
rect 24676 4072 24728 4078
rect 24676 4014 24728 4020
rect 24122 2816 24178 2825
rect 24122 2751 24178 2760
rect 24400 1012 24452 1018
rect 24400 954 24452 960
rect 24124 944 24176 950
rect 24124 886 24176 892
rect 24136 800 24164 886
rect 24412 800 24440 954
rect 24688 800 24716 4014
rect 25332 3738 25360 5646
rect 25884 5370 25912 8366
rect 26068 6798 26096 8434
rect 26528 8401 26556 8570
rect 26514 8392 26570 8401
rect 26514 8327 26570 8336
rect 26698 8120 26754 8129
rect 26698 8055 26754 8064
rect 26712 7886 26740 8055
rect 26424 7880 26476 7886
rect 26424 7822 26476 7828
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26056 6792 26108 6798
rect 25976 6740 26056 6746
rect 25976 6734 26108 6740
rect 25976 6718 26096 6734
rect 25872 5364 25924 5370
rect 25872 5306 25924 5312
rect 25778 4040 25834 4049
rect 25778 3975 25834 3984
rect 24952 3732 25004 3738
rect 24952 3674 25004 3680
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 24964 2922 24992 3674
rect 25136 3596 25188 3602
rect 25136 3538 25188 3544
rect 25148 3398 25176 3538
rect 25792 3534 25820 3975
rect 25780 3528 25832 3534
rect 25780 3470 25832 3476
rect 25044 3392 25096 3398
rect 25044 3334 25096 3340
rect 25136 3392 25188 3398
rect 25136 3334 25188 3340
rect 25056 3194 25084 3334
rect 25044 3188 25096 3194
rect 25044 3130 25096 3136
rect 24952 2916 25004 2922
rect 24952 2858 25004 2864
rect 25228 2916 25280 2922
rect 25228 2858 25280 2864
rect 24768 2372 24820 2378
rect 24768 2314 24820 2320
rect 24780 898 24808 2314
rect 24780 870 24992 898
rect 24964 800 24992 870
rect 25240 800 25268 2858
rect 25976 2650 26004 6718
rect 26056 6112 26108 6118
rect 26056 6054 26108 6060
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 26068 5914 26096 6054
rect 26056 5908 26108 5914
rect 26056 5850 26108 5856
rect 26056 5772 26108 5778
rect 26056 5714 26108 5720
rect 26068 5574 26096 5714
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 26068 3398 26096 5510
rect 26160 5234 26188 6054
rect 26436 5778 26464 7822
rect 26608 7812 26660 7818
rect 26608 7754 26660 7760
rect 26516 7200 26568 7206
rect 26516 7142 26568 7148
rect 26528 6866 26556 7142
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 26620 6254 26648 7754
rect 26712 7449 26740 7822
rect 26698 7440 26754 7449
rect 26698 7375 26754 7384
rect 26804 6730 26832 8735
rect 26882 8392 26938 8401
rect 26882 8327 26938 8336
rect 26792 6724 26844 6730
rect 26792 6666 26844 6672
rect 26608 6248 26660 6254
rect 26608 6190 26660 6196
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 26804 5642 26832 6666
rect 26792 5636 26844 5642
rect 26792 5578 26844 5584
rect 26896 5302 26924 8327
rect 26974 6896 27030 6905
rect 26974 6831 27030 6840
rect 26988 6798 27016 6831
rect 26976 6792 27028 6798
rect 26976 6734 27028 6740
rect 26988 5710 27016 6734
rect 26976 5704 27028 5710
rect 26976 5646 27028 5652
rect 26884 5296 26936 5302
rect 26884 5238 26936 5244
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 26240 5024 26292 5030
rect 26240 4966 26292 4972
rect 26056 3392 26108 3398
rect 26056 3334 26108 3340
rect 26252 2774 26280 4966
rect 26332 4616 26384 4622
rect 26332 4558 26384 4564
rect 26068 2746 26280 2774
rect 25780 2644 25832 2650
rect 25780 2586 25832 2592
rect 25964 2644 26016 2650
rect 25964 2586 26016 2592
rect 25504 2372 25556 2378
rect 25504 2314 25556 2320
rect 25516 800 25544 2314
rect 25792 800 25820 2586
rect 26068 800 26096 2746
rect 26344 800 26372 4558
rect 26884 4480 26936 4486
rect 26884 4422 26936 4428
rect 26792 3460 26844 3466
rect 26792 3402 26844 3408
rect 26608 2848 26660 2854
rect 26608 2790 26660 2796
rect 26424 2372 26476 2378
rect 26424 2314 26476 2320
rect 26436 1018 26464 2314
rect 26424 1012 26476 1018
rect 26424 954 26476 960
rect 26620 800 26648 2790
rect 26804 1834 26832 3402
rect 26792 1828 26844 1834
rect 26792 1770 26844 1776
rect 26896 800 26924 4422
rect 26976 3460 27028 3466
rect 26976 3402 27028 3408
rect 26988 3058 27016 3402
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 27080 2774 27108 9862
rect 27172 7750 27200 10367
rect 27264 8498 27292 15982
rect 27356 11812 27384 17478
rect 27448 15094 27476 18788
rect 27528 18770 27580 18776
rect 27632 18426 27660 20742
rect 27816 20602 27844 20878
rect 27804 20596 27856 20602
rect 27804 20538 27856 20544
rect 27804 18760 27856 18766
rect 27804 18702 27856 18708
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 27620 18420 27672 18426
rect 27620 18362 27672 18368
rect 27724 18222 27752 18566
rect 27712 18216 27764 18222
rect 27712 18158 27764 18164
rect 27712 18080 27764 18086
rect 27712 18022 27764 18028
rect 27620 17196 27672 17202
rect 27620 17138 27672 17144
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27540 16250 27568 16594
rect 27528 16244 27580 16250
rect 27528 16186 27580 16192
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27436 15088 27488 15094
rect 27436 15030 27488 15036
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27448 14278 27476 14894
rect 27436 14272 27488 14278
rect 27436 14214 27488 14220
rect 27540 13530 27568 15438
rect 27528 13524 27580 13530
rect 27528 13466 27580 13472
rect 27632 12442 27660 17138
rect 27724 17066 27752 18022
rect 27712 17060 27764 17066
rect 27712 17002 27764 17008
rect 27712 16448 27764 16454
rect 27712 16390 27764 16396
rect 27724 15026 27752 16390
rect 27712 15020 27764 15026
rect 27712 14962 27764 14968
rect 27710 14648 27766 14657
rect 27710 14583 27766 14592
rect 27724 13530 27752 14583
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27816 12986 27844 18702
rect 27908 17746 27936 26930
rect 29000 26444 29052 26450
rect 29000 26386 29052 26392
rect 29012 25770 29040 26386
rect 29000 25764 29052 25770
rect 29000 25706 29052 25712
rect 27988 23520 28040 23526
rect 27988 23462 28040 23468
rect 28000 19854 28028 23462
rect 29276 23180 29328 23186
rect 29276 23122 29328 23128
rect 28632 21548 28684 21554
rect 28632 21490 28684 21496
rect 28644 21146 28672 21490
rect 28908 21480 28960 21486
rect 28908 21422 28960 21428
rect 28632 21140 28684 21146
rect 28632 21082 28684 21088
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28448 20596 28500 20602
rect 28448 20538 28500 20544
rect 27988 19848 28040 19854
rect 27988 19790 28040 19796
rect 28000 17921 28028 19790
rect 28080 19712 28132 19718
rect 28080 19654 28132 19660
rect 28092 19174 28120 19654
rect 28080 19168 28132 19174
rect 28080 19110 28132 19116
rect 28092 18290 28120 19110
rect 28460 18766 28488 20538
rect 28644 19922 28672 20878
rect 28920 20602 28948 21422
rect 29184 21072 29236 21078
rect 29184 21014 29236 21020
rect 28998 20632 29054 20641
rect 28908 20596 28960 20602
rect 28998 20567 29054 20576
rect 28908 20538 28960 20544
rect 29012 20466 29040 20567
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29092 20392 29144 20398
rect 28920 20340 29092 20346
rect 28920 20334 29144 20340
rect 28920 20318 29132 20334
rect 28920 19961 28948 20318
rect 28906 19952 28962 19961
rect 28632 19916 28684 19922
rect 28906 19887 28962 19896
rect 28632 19858 28684 19864
rect 28448 18760 28500 18766
rect 28448 18702 28500 18708
rect 28538 18728 28594 18737
rect 28538 18663 28540 18672
rect 28592 18663 28594 18672
rect 28540 18634 28592 18640
rect 28080 18284 28132 18290
rect 28080 18226 28132 18232
rect 28080 18080 28132 18086
rect 28080 18022 28132 18028
rect 27986 17912 28042 17921
rect 27986 17847 28042 17856
rect 27896 17740 27948 17746
rect 27896 17682 27948 17688
rect 27988 17672 28040 17678
rect 27988 17614 28040 17620
rect 28000 17202 28028 17614
rect 27988 17196 28040 17202
rect 27988 17138 28040 17144
rect 27896 17060 27948 17066
rect 27896 17002 27948 17008
rect 27908 16046 27936 17002
rect 27896 16040 27948 16046
rect 27896 15982 27948 15988
rect 27986 15600 28042 15609
rect 27986 15535 28042 15544
rect 27896 15428 27948 15434
rect 27896 15370 27948 15376
rect 27908 15162 27936 15370
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 28000 14385 28028 15535
rect 27986 14376 28042 14385
rect 27986 14311 28042 14320
rect 27804 12980 27856 12986
rect 27804 12922 27856 12928
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 27620 12436 27672 12442
rect 27620 12378 27672 12384
rect 27816 12238 27844 12786
rect 27988 12708 28040 12714
rect 27988 12650 28040 12656
rect 27804 12232 27856 12238
rect 27804 12174 27856 12180
rect 27528 11824 27580 11830
rect 27356 11784 27528 11812
rect 27528 11766 27580 11772
rect 27344 11144 27396 11150
rect 27342 11112 27344 11121
rect 27436 11144 27488 11150
rect 27396 11112 27398 11121
rect 27436 11086 27488 11092
rect 27342 11047 27398 11056
rect 27448 10577 27476 11086
rect 27540 11082 27568 11766
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 27804 10736 27856 10742
rect 27804 10678 27856 10684
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27434 10568 27490 10577
rect 27434 10503 27490 10512
rect 27344 10056 27396 10062
rect 27344 9998 27396 10004
rect 27356 9353 27384 9998
rect 27528 9988 27580 9994
rect 27528 9930 27580 9936
rect 27540 9722 27568 9930
rect 27528 9716 27580 9722
rect 27528 9658 27580 9664
rect 27342 9344 27398 9353
rect 27342 9279 27398 9288
rect 27632 9194 27660 10610
rect 27816 10606 27844 10678
rect 27896 10668 27948 10674
rect 27896 10610 27948 10616
rect 27804 10600 27856 10606
rect 27804 10542 27856 10548
rect 27710 10296 27766 10305
rect 27710 10231 27766 10240
rect 27724 10198 27752 10231
rect 27712 10192 27764 10198
rect 27712 10134 27764 10140
rect 27712 9648 27764 9654
rect 27712 9590 27764 9596
rect 27540 9166 27660 9194
rect 27540 8922 27568 9166
rect 27618 9072 27674 9081
rect 27618 9007 27674 9016
rect 27448 8894 27568 8922
rect 27252 8492 27304 8498
rect 27252 8434 27304 8440
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 27160 7744 27212 7750
rect 27160 7686 27212 7692
rect 27172 6866 27200 7686
rect 27250 7168 27306 7177
rect 27250 7103 27306 7112
rect 27160 6860 27212 6866
rect 27160 6802 27212 6808
rect 27264 6304 27292 7103
rect 27356 6905 27384 8434
rect 27448 8294 27476 8894
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27436 8288 27488 8294
rect 27436 8230 27488 8236
rect 27436 7948 27488 7954
rect 27436 7890 27488 7896
rect 27342 6896 27398 6905
rect 27342 6831 27398 6840
rect 27344 6316 27396 6322
rect 27264 6276 27344 6304
rect 27344 6258 27396 6264
rect 27356 6089 27384 6258
rect 27342 6080 27398 6089
rect 27342 6015 27398 6024
rect 27448 4214 27476 7890
rect 27540 5234 27568 8774
rect 27632 8498 27660 9007
rect 27724 8906 27752 9590
rect 27712 8900 27764 8906
rect 27712 8842 27764 8848
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27724 8498 27752 8570
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27816 8378 27844 10542
rect 27908 9178 27936 10610
rect 28000 10470 28028 12650
rect 28092 12434 28120 18022
rect 28540 17808 28592 17814
rect 28540 17750 28592 17756
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 28172 17264 28224 17270
rect 28224 17212 28304 17218
rect 28172 17206 28304 17212
rect 28184 17190 28304 17206
rect 28276 16436 28304 17190
rect 28368 17105 28396 17614
rect 28448 17264 28500 17270
rect 28448 17206 28500 17212
rect 28354 17096 28410 17105
rect 28354 17031 28410 17040
rect 28460 16658 28488 17206
rect 28448 16652 28500 16658
rect 28448 16594 28500 16600
rect 28356 16448 28408 16454
rect 28276 16408 28356 16436
rect 28356 16390 28408 16396
rect 28368 16114 28396 16390
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28172 16040 28224 16046
rect 28172 15982 28224 15988
rect 28184 13870 28212 15982
rect 28368 15366 28396 16050
rect 28552 15722 28580 17750
rect 28644 16658 28672 19858
rect 29196 18970 29224 21014
rect 29288 19174 29316 23122
rect 29276 19168 29328 19174
rect 29276 19110 29328 19116
rect 29184 18964 29236 18970
rect 29184 18906 29236 18912
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 28724 17536 28776 17542
rect 28724 17478 28776 17484
rect 28632 16652 28684 16658
rect 28632 16594 28684 16600
rect 28736 15994 28764 17478
rect 28828 17202 28856 18702
rect 28908 17604 28960 17610
rect 28908 17546 28960 17552
rect 28816 17196 28868 17202
rect 28816 17138 28868 17144
rect 28920 16794 28948 17546
rect 29000 17128 29052 17134
rect 29000 17070 29052 17076
rect 29012 16794 29040 17070
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 28908 16788 28960 16794
rect 28908 16730 28960 16736
rect 29000 16788 29052 16794
rect 29000 16730 29052 16736
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 28736 15966 28948 15994
rect 28724 15904 28776 15910
rect 28724 15846 28776 15852
rect 28552 15694 28672 15722
rect 28540 15632 28592 15638
rect 28540 15574 28592 15580
rect 28356 15360 28408 15366
rect 28356 15302 28408 15308
rect 28172 13864 28224 13870
rect 28172 13806 28224 13812
rect 28552 13326 28580 15574
rect 28644 14940 28672 15694
rect 28736 15094 28764 15846
rect 28724 15088 28776 15094
rect 28724 15030 28776 15036
rect 28644 14912 28764 14940
rect 28540 13320 28592 13326
rect 28540 13262 28592 13268
rect 28632 13252 28684 13258
rect 28632 13194 28684 13200
rect 28644 12918 28672 13194
rect 28632 12912 28684 12918
rect 28632 12854 28684 12860
rect 28092 12406 28212 12434
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 27988 10464 28040 10470
rect 27988 10406 28040 10412
rect 27896 9172 27948 9178
rect 27896 9114 27948 9120
rect 27896 8968 27948 8974
rect 28000 8956 28028 10406
rect 27948 8928 28028 8956
rect 27896 8910 27948 8916
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 27724 8350 27844 8378
rect 27620 8288 27672 8294
rect 27620 8230 27672 8236
rect 27632 6866 27660 8230
rect 27724 7342 27752 8350
rect 27896 8288 27948 8294
rect 27896 8230 27948 8236
rect 27804 8016 27856 8022
rect 27804 7958 27856 7964
rect 27712 7336 27764 7342
rect 27712 7278 27764 7284
rect 27620 6860 27672 6866
rect 27620 6802 27672 6808
rect 27632 6322 27660 6802
rect 27816 6730 27844 7958
rect 27908 7818 27936 8230
rect 27896 7812 27948 7818
rect 27896 7754 27948 7760
rect 27908 7002 27936 7754
rect 28000 7342 28028 8434
rect 27988 7336 28040 7342
rect 27988 7278 28040 7284
rect 27988 7200 28040 7206
rect 27988 7142 28040 7148
rect 27896 6996 27948 7002
rect 27896 6938 27948 6944
rect 27804 6724 27856 6730
rect 27804 6666 27856 6672
rect 27802 6624 27858 6633
rect 27802 6559 27858 6568
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 27528 5228 27580 5234
rect 27528 5170 27580 5176
rect 27528 5024 27580 5030
rect 27528 4966 27580 4972
rect 27160 4208 27212 4214
rect 27160 4150 27212 4156
rect 27436 4208 27488 4214
rect 27436 4150 27488 4156
rect 26988 2746 27108 2774
rect 26988 2038 27016 2746
rect 26976 2032 27028 2038
rect 26976 1974 27028 1980
rect 27172 800 27200 4150
rect 27540 4146 27568 4966
rect 27632 4690 27660 6258
rect 27816 6254 27844 6559
rect 27804 6248 27856 6254
rect 27804 6190 27856 6196
rect 28000 6118 28028 7142
rect 28092 6866 28120 11018
rect 28184 9722 28212 12406
rect 28264 12232 28316 12238
rect 28264 12174 28316 12180
rect 28276 11082 28304 12174
rect 28448 12164 28500 12170
rect 28448 12106 28500 12112
rect 28264 11076 28316 11082
rect 28264 11018 28316 11024
rect 28264 10668 28316 10674
rect 28264 10610 28316 10616
rect 28276 10577 28304 10610
rect 28262 10568 28318 10577
rect 28262 10503 28318 10512
rect 28264 10124 28316 10130
rect 28264 10066 28316 10072
rect 28172 9716 28224 9722
rect 28172 9658 28224 9664
rect 28172 9580 28224 9586
rect 28172 9522 28224 9528
rect 28184 8498 28212 9522
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 28276 8430 28304 10066
rect 28356 9920 28408 9926
rect 28356 9862 28408 9868
rect 28264 8424 28316 8430
rect 28264 8366 28316 8372
rect 28264 8288 28316 8294
rect 28264 8230 28316 8236
rect 28276 7857 28304 8230
rect 28368 8106 28396 9862
rect 28460 9654 28488 12106
rect 28644 11626 28672 12854
rect 28632 11620 28684 11626
rect 28632 11562 28684 11568
rect 28540 10668 28592 10674
rect 28540 10610 28592 10616
rect 28448 9648 28500 9654
rect 28448 9590 28500 9596
rect 28446 9480 28502 9489
rect 28446 9415 28448 9424
rect 28500 9415 28502 9424
rect 28448 9386 28500 9392
rect 28368 8078 28488 8106
rect 28356 8016 28408 8022
rect 28356 7958 28408 7964
rect 28262 7848 28318 7857
rect 28262 7783 28318 7792
rect 28262 7304 28318 7313
rect 28262 7239 28264 7248
rect 28316 7239 28318 7248
rect 28264 7210 28316 7216
rect 28368 7002 28396 7958
rect 28356 6996 28408 7002
rect 28356 6938 28408 6944
rect 28080 6860 28132 6866
rect 28080 6802 28132 6808
rect 28368 6186 28396 6938
rect 28460 6746 28488 8078
rect 28552 7546 28580 10610
rect 28540 7540 28592 7546
rect 28540 7482 28592 7488
rect 28644 7478 28672 11562
rect 28736 8634 28764 14912
rect 28816 13932 28868 13938
rect 28816 13874 28868 13880
rect 28828 13462 28856 13874
rect 28816 13456 28868 13462
rect 28816 13398 28868 13404
rect 28816 10668 28868 10674
rect 28816 10610 28868 10616
rect 28828 10577 28856 10610
rect 28814 10568 28870 10577
rect 28814 10503 28870 10512
rect 28920 9926 28948 15966
rect 29012 15026 29040 16594
rect 29092 15088 29144 15094
rect 29092 15030 29144 15036
rect 29000 15020 29052 15026
rect 29000 14962 29052 14968
rect 29012 9994 29040 14962
rect 29104 14482 29132 15030
rect 29092 14476 29144 14482
rect 29092 14418 29144 14424
rect 29104 14074 29132 14418
rect 29092 14068 29144 14074
rect 29092 14010 29144 14016
rect 29092 12300 29144 12306
rect 29092 12242 29144 12248
rect 29000 9988 29052 9994
rect 29000 9930 29052 9936
rect 28908 9920 28960 9926
rect 28908 9862 28960 9868
rect 28908 9580 28960 9586
rect 28908 9522 28960 9528
rect 28816 9036 28868 9042
rect 28816 8978 28868 8984
rect 28724 8628 28776 8634
rect 28724 8570 28776 8576
rect 28736 8430 28764 8570
rect 28724 8424 28776 8430
rect 28724 8366 28776 8372
rect 28632 7472 28684 7478
rect 28632 7414 28684 7420
rect 28632 6860 28684 6866
rect 28632 6802 28684 6808
rect 28460 6730 28580 6746
rect 28460 6724 28592 6730
rect 28460 6718 28540 6724
rect 28540 6666 28592 6672
rect 28448 6656 28500 6662
rect 28448 6598 28500 6604
rect 28356 6180 28408 6186
rect 28356 6122 28408 6128
rect 27988 6112 28040 6118
rect 27988 6054 28040 6060
rect 27712 5840 27764 5846
rect 27710 5808 27712 5817
rect 27764 5808 27766 5817
rect 27710 5743 27766 5752
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 27804 4616 27856 4622
rect 27804 4558 27856 4564
rect 27344 4140 27396 4146
rect 27344 4082 27396 4088
rect 27528 4140 27580 4146
rect 27528 4082 27580 4088
rect 27252 3732 27304 3738
rect 27252 3674 27304 3680
rect 27264 3398 27292 3674
rect 27356 3534 27384 4082
rect 27816 3738 27844 4558
rect 27896 4140 27948 4146
rect 27896 4082 27948 4088
rect 27804 3732 27856 3738
rect 27804 3674 27856 3680
rect 27344 3528 27396 3534
rect 27344 3470 27396 3476
rect 27908 3448 27936 4082
rect 28000 3602 28028 6054
rect 28172 5024 28224 5030
rect 28172 4966 28224 4972
rect 27988 3596 28040 3602
rect 27988 3538 28040 3544
rect 27724 3420 27936 3448
rect 27988 3460 28040 3466
rect 27252 3392 27304 3398
rect 27252 3334 27304 3340
rect 27526 3088 27582 3097
rect 27526 3023 27528 3032
rect 27580 3023 27582 3032
rect 27528 2994 27580 3000
rect 27344 2984 27396 2990
rect 27344 2926 27396 2932
rect 27356 1086 27384 2926
rect 27540 2854 27568 2994
rect 27528 2848 27580 2854
rect 27528 2790 27580 2796
rect 27436 2508 27488 2514
rect 27436 2450 27488 2456
rect 27344 1080 27396 1086
rect 27344 1022 27396 1028
rect 27448 800 27476 2450
rect 27620 2372 27672 2378
rect 27620 2314 27672 2320
rect 27528 2304 27580 2310
rect 27528 2246 27580 2252
rect 27540 950 27568 2246
rect 27632 1902 27660 2314
rect 27620 1896 27672 1902
rect 27620 1838 27672 1844
rect 27528 944 27580 950
rect 27528 886 27580 892
rect 27724 800 27752 3420
rect 27988 3402 28040 3408
rect 27804 2984 27856 2990
rect 27804 2926 27856 2932
rect 27816 1154 27844 2926
rect 27804 1148 27856 1154
rect 27804 1090 27856 1096
rect 28000 800 28028 3402
rect 28184 2514 28212 4966
rect 28460 4570 28488 6598
rect 28552 6390 28580 6666
rect 28540 6384 28592 6390
rect 28540 6326 28592 6332
rect 28552 5692 28580 6326
rect 28644 6322 28672 6802
rect 28724 6656 28776 6662
rect 28722 6624 28724 6633
rect 28776 6624 28778 6633
rect 28722 6559 28778 6568
rect 28632 6316 28684 6322
rect 28632 6258 28684 6264
rect 28828 5760 28856 8978
rect 28920 8922 28948 9522
rect 29012 9042 29040 9930
rect 29104 9450 29132 12242
rect 29196 9654 29224 16934
rect 29288 11762 29316 19110
rect 29460 18828 29512 18834
rect 29460 18770 29512 18776
rect 29472 18290 29500 18770
rect 29564 18290 29592 50322
rect 29644 39364 29696 39370
rect 29644 39306 29696 39312
rect 29460 18284 29512 18290
rect 29460 18226 29512 18232
rect 29552 18284 29604 18290
rect 29552 18226 29604 18232
rect 29552 16176 29604 16182
rect 29552 16118 29604 16124
rect 29564 16017 29592 16118
rect 29550 16008 29606 16017
rect 29550 15943 29606 15952
rect 29564 15162 29592 15943
rect 29460 15156 29512 15162
rect 29460 15098 29512 15104
rect 29552 15156 29604 15162
rect 29552 15098 29604 15104
rect 29472 14890 29500 15098
rect 29460 14884 29512 14890
rect 29460 14826 29512 14832
rect 29368 14408 29420 14414
rect 29368 14350 29420 14356
rect 29380 14074 29408 14350
rect 29460 14272 29512 14278
rect 29460 14214 29512 14220
rect 29368 14068 29420 14074
rect 29368 14010 29420 14016
rect 29472 13802 29500 14214
rect 29552 13932 29604 13938
rect 29552 13874 29604 13880
rect 29460 13796 29512 13802
rect 29460 13738 29512 13744
rect 29564 12434 29592 13874
rect 29472 12406 29592 12434
rect 29276 11756 29328 11762
rect 29276 11698 29328 11704
rect 29276 11552 29328 11558
rect 29276 11494 29328 11500
rect 29368 11552 29420 11558
rect 29368 11494 29420 11500
rect 29288 10606 29316 11494
rect 29276 10600 29328 10606
rect 29276 10542 29328 10548
rect 29184 9648 29236 9654
rect 29184 9590 29236 9596
rect 29184 9512 29236 9518
rect 29184 9454 29236 9460
rect 29274 9480 29330 9489
rect 29092 9444 29144 9450
rect 29092 9386 29144 9392
rect 29000 9036 29052 9042
rect 29000 8978 29052 8984
rect 29092 9036 29144 9042
rect 29092 8978 29144 8984
rect 28920 8894 29040 8922
rect 28908 6180 28960 6186
rect 28908 6122 28960 6128
rect 28920 5846 28948 6122
rect 28908 5840 28960 5846
rect 28908 5782 28960 5788
rect 28736 5732 28856 5760
rect 28632 5704 28684 5710
rect 28552 5664 28632 5692
rect 28632 5646 28684 5652
rect 28736 5250 28764 5732
rect 28816 5636 28868 5642
rect 28868 5596 28948 5624
rect 28816 5578 28868 5584
rect 28540 5228 28592 5234
rect 28736 5222 28856 5250
rect 28592 5188 28672 5216
rect 28540 5170 28592 5176
rect 28368 4542 28488 4570
rect 28368 4282 28396 4542
rect 28540 4480 28592 4486
rect 28540 4422 28592 4428
rect 28356 4276 28408 4282
rect 28356 4218 28408 4224
rect 28262 4176 28318 4185
rect 28262 4111 28318 4120
rect 28276 3602 28304 4111
rect 28264 3596 28316 3602
rect 28264 3538 28316 3544
rect 28172 2508 28224 2514
rect 28172 2450 28224 2456
rect 28368 2446 28396 4218
rect 28448 3936 28500 3942
rect 28448 3878 28500 3884
rect 28460 3738 28488 3878
rect 28448 3732 28500 3738
rect 28448 3674 28500 3680
rect 28460 3058 28488 3674
rect 28552 3126 28580 4422
rect 28644 3942 28672 5188
rect 28724 5160 28776 5166
rect 28724 5102 28776 5108
rect 28736 4690 28764 5102
rect 28724 4684 28776 4690
rect 28724 4626 28776 4632
rect 28724 4480 28776 4486
rect 28722 4448 28724 4457
rect 28776 4448 28778 4457
rect 28722 4383 28778 4392
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28644 3534 28672 3878
rect 28828 3602 28856 5222
rect 28816 3596 28868 3602
rect 28816 3538 28868 3544
rect 28632 3528 28684 3534
rect 28632 3470 28684 3476
rect 28540 3120 28592 3126
rect 28540 3062 28592 3068
rect 28448 3052 28500 3058
rect 28448 2994 28500 3000
rect 28920 2582 28948 5596
rect 29012 5409 29040 8894
rect 29104 8566 29132 8978
rect 29196 8974 29224 9454
rect 29274 9415 29330 9424
rect 29288 9382 29316 9415
rect 29276 9376 29328 9382
rect 29276 9318 29328 9324
rect 29184 8968 29236 8974
rect 29184 8910 29236 8916
rect 29182 8800 29238 8809
rect 29182 8735 29238 8744
rect 29092 8560 29144 8566
rect 29092 8502 29144 8508
rect 29196 8498 29224 8735
rect 29184 8492 29236 8498
rect 29184 8434 29236 8440
rect 29288 8072 29316 9318
rect 29380 8090 29408 11494
rect 29472 11257 29500 12406
rect 29656 11762 29684 39306
rect 29748 35894 29776 55626
rect 29748 35866 29868 35894
rect 29736 18828 29788 18834
rect 29736 18770 29788 18776
rect 29748 18426 29776 18770
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 29736 18284 29788 18290
rect 29736 18226 29788 18232
rect 29748 17660 29776 18226
rect 29840 18193 29868 35866
rect 29932 18465 29960 60998
rect 30300 60734 30328 61678
rect 30116 60706 30328 60734
rect 30484 60722 30512 63242
rect 31022 63200 31078 63294
rect 31220 61198 31248 63294
rect 31758 63200 31814 64000
rect 32494 63322 32550 64000
rect 32494 63306 32628 63322
rect 32494 63300 32640 63306
rect 32494 63294 32588 63300
rect 32494 63200 32550 63294
rect 32588 63242 32640 63248
rect 33230 63200 33286 64000
rect 33966 63322 34022 64000
rect 33966 63306 34100 63322
rect 33324 63300 33376 63306
rect 33324 63242 33376 63248
rect 33966 63300 34112 63306
rect 33966 63294 34060 63300
rect 31772 61198 31800 63200
rect 32956 61260 33008 61266
rect 32956 61202 33008 61208
rect 31208 61192 31260 61198
rect 31208 61134 31260 61140
rect 31760 61192 31812 61198
rect 31760 61134 31812 61140
rect 31300 61056 31352 61062
rect 31300 60998 31352 61004
rect 32588 61056 32640 61062
rect 32588 60998 32640 61004
rect 30472 60716 30524 60722
rect 30012 60512 30064 60518
rect 30012 60454 30064 60460
rect 30024 60042 30052 60454
rect 30012 60036 30064 60042
rect 30012 59978 30064 59984
rect 30116 59702 30144 60706
rect 30472 60658 30524 60664
rect 30564 60716 30616 60722
rect 30564 60658 30616 60664
rect 30576 60246 30604 60658
rect 31208 60648 31260 60654
rect 31208 60590 31260 60596
rect 30932 60512 30984 60518
rect 30932 60454 30984 60460
rect 30564 60240 30616 60246
rect 30564 60182 30616 60188
rect 30748 60240 30800 60246
rect 30748 60182 30800 60188
rect 30760 60110 30788 60182
rect 30944 60110 30972 60454
rect 31220 60110 31248 60590
rect 30196 60104 30248 60110
rect 30196 60046 30248 60052
rect 30748 60104 30800 60110
rect 30748 60046 30800 60052
rect 30932 60104 30984 60110
rect 31116 60104 31168 60110
rect 30932 60046 30984 60052
rect 31114 60072 31116 60081
rect 31208 60104 31260 60110
rect 31168 60072 31170 60081
rect 30104 59696 30156 59702
rect 30104 59638 30156 59644
rect 30208 59634 30236 60046
rect 31208 60046 31260 60052
rect 31114 60007 31170 60016
rect 30472 59968 30524 59974
rect 30524 59928 30604 59956
rect 30472 59910 30524 59916
rect 30288 59696 30340 59702
rect 30288 59638 30340 59644
rect 30012 59628 30064 59634
rect 30012 59570 30064 59576
rect 30196 59628 30248 59634
rect 30196 59570 30248 59576
rect 30024 59430 30052 59570
rect 30300 59498 30328 59638
rect 30288 59492 30340 59498
rect 30288 59434 30340 59440
rect 30380 59492 30432 59498
rect 30380 59434 30432 59440
rect 30012 59424 30064 59430
rect 30012 59366 30064 59372
rect 30392 55758 30420 59434
rect 30472 55956 30524 55962
rect 30472 55898 30524 55904
rect 30484 55758 30512 55898
rect 30576 55826 30604 59928
rect 30654 59528 30710 59537
rect 30654 59463 30710 59472
rect 30668 59430 30696 59463
rect 30656 59424 30708 59430
rect 30656 59366 30708 59372
rect 30564 55820 30616 55826
rect 30564 55762 30616 55768
rect 30380 55752 30432 55758
rect 30380 55694 30432 55700
rect 30472 55752 30524 55758
rect 30472 55694 30524 55700
rect 30668 47734 30696 59366
rect 31312 47802 31340 60998
rect 32220 59968 32272 59974
rect 32218 59936 32220 59945
rect 32496 59968 32548 59974
rect 32272 59936 32274 59945
rect 32496 59910 32548 59916
rect 32218 59871 32274 59880
rect 32508 59430 32536 59910
rect 32496 59424 32548 59430
rect 32496 59366 32548 59372
rect 31300 47796 31352 47802
rect 31300 47738 31352 47744
rect 30656 47728 30708 47734
rect 30656 47670 30708 47676
rect 32220 47592 32272 47598
rect 32220 47534 32272 47540
rect 31760 43104 31812 43110
rect 31760 43046 31812 43052
rect 31116 37324 31168 37330
rect 31116 37266 31168 37272
rect 31024 33652 31076 33658
rect 31024 33594 31076 33600
rect 31036 33318 31064 33594
rect 31024 33312 31076 33318
rect 31024 33254 31076 33260
rect 30380 30184 30432 30190
rect 30380 30126 30432 30132
rect 30392 26926 30420 30126
rect 30840 29028 30892 29034
rect 30840 28970 30892 28976
rect 30380 26920 30432 26926
rect 30380 26862 30432 26868
rect 30656 20936 30708 20942
rect 30656 20878 30708 20884
rect 30748 20936 30800 20942
rect 30748 20878 30800 20884
rect 30668 20466 30696 20878
rect 30760 20602 30788 20878
rect 30748 20596 30800 20602
rect 30748 20538 30800 20544
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30208 19854 30236 20402
rect 30748 20392 30800 20398
rect 30748 20334 30800 20340
rect 30760 20262 30788 20334
rect 30748 20256 30800 20262
rect 30748 20198 30800 20204
rect 30196 19848 30248 19854
rect 30196 19790 30248 19796
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 30208 18766 30236 19790
rect 30300 19378 30328 19790
rect 30288 19372 30340 19378
rect 30288 19314 30340 19320
rect 30564 19372 30616 19378
rect 30564 19314 30616 19320
rect 30576 18970 30604 19314
rect 30564 18964 30616 18970
rect 30564 18906 30616 18912
rect 30748 18828 30800 18834
rect 30748 18770 30800 18776
rect 30196 18760 30248 18766
rect 30196 18702 30248 18708
rect 30012 18624 30064 18630
rect 30012 18566 30064 18572
rect 29918 18456 29974 18465
rect 29918 18391 29974 18400
rect 30024 18290 30052 18566
rect 30012 18284 30064 18290
rect 30012 18226 30064 18232
rect 29826 18184 29882 18193
rect 29826 18119 29882 18128
rect 29828 17808 29880 17814
rect 29826 17776 29828 17785
rect 29880 17776 29882 17785
rect 29826 17711 29882 17720
rect 30012 17672 30064 17678
rect 29748 17632 30012 17660
rect 30012 17614 30064 17620
rect 30024 16658 30052 17614
rect 30012 16652 30064 16658
rect 30012 16594 30064 16600
rect 29734 16280 29790 16289
rect 29734 16215 29790 16224
rect 29748 16046 29776 16215
rect 29736 16040 29788 16046
rect 29736 15982 29788 15988
rect 30010 15328 30066 15337
rect 30010 15263 30066 15272
rect 29736 14816 29788 14822
rect 29736 14758 29788 14764
rect 29748 14482 29776 14758
rect 29736 14476 29788 14482
rect 29736 14418 29788 14424
rect 29748 12986 29776 14418
rect 29920 14068 29972 14074
rect 29920 14010 29972 14016
rect 29828 13864 29880 13870
rect 29828 13806 29880 13812
rect 29840 13161 29868 13806
rect 29826 13152 29882 13161
rect 29826 13087 29882 13096
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 29748 12782 29776 12922
rect 29736 12776 29788 12782
rect 29736 12718 29788 12724
rect 29932 12374 29960 14010
rect 30024 12442 30052 15263
rect 30208 15094 30236 18702
rect 30760 18222 30788 18770
rect 30748 18216 30800 18222
rect 30748 18158 30800 18164
rect 30288 17536 30340 17542
rect 30288 17478 30340 17484
rect 30196 15088 30248 15094
rect 30196 15030 30248 15036
rect 30104 13320 30156 13326
rect 30104 13262 30156 13268
rect 30012 12436 30064 12442
rect 30012 12378 30064 12384
rect 29920 12368 29972 12374
rect 29920 12310 29972 12316
rect 30116 12238 30144 13262
rect 30104 12232 30156 12238
rect 29734 12200 29790 12209
rect 30104 12174 30156 12180
rect 29734 12135 29790 12144
rect 29552 11756 29604 11762
rect 29552 11698 29604 11704
rect 29644 11756 29696 11762
rect 29644 11698 29696 11704
rect 29458 11248 29514 11257
rect 29564 11218 29592 11698
rect 29644 11348 29696 11354
rect 29644 11290 29696 11296
rect 29458 11183 29514 11192
rect 29552 11212 29604 11218
rect 29552 11154 29604 11160
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 29460 10056 29512 10062
rect 29460 9998 29512 10004
rect 29196 8044 29316 8072
rect 29368 8084 29420 8090
rect 29196 7954 29224 8044
rect 29368 8026 29420 8032
rect 29184 7948 29236 7954
rect 29184 7890 29236 7896
rect 29276 7948 29328 7954
rect 29276 7890 29328 7896
rect 29288 7818 29316 7890
rect 29276 7812 29328 7818
rect 29276 7754 29328 7760
rect 29092 7744 29144 7750
rect 29092 7686 29144 7692
rect 29104 7410 29132 7686
rect 29092 7404 29144 7410
rect 29092 7346 29144 7352
rect 28998 5400 29054 5409
rect 28998 5335 29054 5344
rect 29104 5166 29132 7346
rect 29288 6322 29316 7754
rect 29380 6390 29408 8026
rect 29368 6384 29420 6390
rect 29368 6326 29420 6332
rect 29276 6316 29328 6322
rect 29276 6258 29328 6264
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 29092 5160 29144 5166
rect 29092 5102 29144 5108
rect 28998 4720 29054 4729
rect 28998 4655 29054 4664
rect 29012 4622 29040 4655
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 29104 2854 29132 5102
rect 29196 4622 29224 5170
rect 29472 4690 29500 9998
rect 29564 8838 29592 10406
rect 29552 8832 29604 8838
rect 29552 8774 29604 8780
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 29564 8265 29592 8434
rect 29550 8256 29606 8265
rect 29550 8191 29606 8200
rect 29656 7290 29684 11290
rect 29748 10130 29776 12135
rect 30300 12102 30328 17478
rect 30470 17232 30526 17241
rect 30470 17167 30526 17176
rect 30380 13864 30432 13870
rect 30380 13806 30432 13812
rect 30288 12096 30340 12102
rect 30288 12038 30340 12044
rect 29828 11892 29880 11898
rect 29828 11834 29880 11840
rect 29840 11762 29868 11834
rect 29828 11756 29880 11762
rect 29828 11698 29880 11704
rect 30300 11393 30328 12038
rect 30286 11384 30342 11393
rect 30286 11319 30342 11328
rect 30196 11076 30248 11082
rect 30196 11018 30248 11024
rect 29736 10124 29788 10130
rect 29736 10066 29788 10072
rect 29920 9988 29972 9994
rect 29920 9930 29972 9936
rect 29736 8900 29788 8906
rect 29736 8842 29788 8848
rect 29828 8900 29880 8906
rect 29828 8842 29880 8848
rect 29564 7262 29684 7290
rect 29748 7562 29776 8842
rect 29840 8362 29868 8842
rect 29932 8786 29960 9930
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 30116 9722 30144 9862
rect 30104 9716 30156 9722
rect 30104 9658 30156 9664
rect 30012 9580 30064 9586
rect 30012 9522 30064 9528
rect 30024 8945 30052 9522
rect 30116 9081 30144 9658
rect 30102 9072 30158 9081
rect 30102 9007 30158 9016
rect 30010 8936 30066 8945
rect 30010 8871 30066 8880
rect 29932 8758 30144 8786
rect 29918 8664 29974 8673
rect 29918 8599 29974 8608
rect 29932 8430 29960 8599
rect 29920 8424 29972 8430
rect 29920 8366 29972 8372
rect 29828 8356 29880 8362
rect 29828 8298 29880 8304
rect 30012 8356 30064 8362
rect 30012 8298 30064 8304
rect 30024 7886 30052 8298
rect 30012 7880 30064 7886
rect 30012 7822 30064 7828
rect 29748 7546 30052 7562
rect 29748 7540 30064 7546
rect 29748 7534 30012 7540
rect 29748 7274 29776 7534
rect 30012 7482 30064 7488
rect 29736 7268 29788 7274
rect 29460 4684 29512 4690
rect 29460 4626 29512 4632
rect 29184 4616 29236 4622
rect 29184 4558 29236 4564
rect 29564 4282 29592 7262
rect 29736 7210 29788 7216
rect 29920 7268 29972 7274
rect 29920 7210 29972 7216
rect 29644 7200 29696 7206
rect 29644 7142 29696 7148
rect 29656 5794 29684 7142
rect 29932 6186 29960 7210
rect 30012 6928 30064 6934
rect 30012 6870 30064 6876
rect 29920 6180 29972 6186
rect 29920 6122 29972 6128
rect 29656 5766 29776 5794
rect 29644 5704 29696 5710
rect 29642 5672 29644 5681
rect 29696 5672 29698 5681
rect 29642 5607 29698 5616
rect 29656 4758 29684 5607
rect 29644 4752 29696 4758
rect 29644 4694 29696 4700
rect 29552 4276 29604 4282
rect 29552 4218 29604 4224
rect 29644 4072 29696 4078
rect 29644 4014 29696 4020
rect 29092 2848 29144 2854
rect 29092 2790 29144 2796
rect 28908 2576 28960 2582
rect 28908 2518 28960 2524
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 28908 2372 28960 2378
rect 28908 2314 28960 2320
rect 28540 1080 28592 1086
rect 28540 1022 28592 1028
rect 28264 944 28316 950
rect 28264 886 28316 892
rect 28276 800 28304 886
rect 28552 800 28580 1022
rect 28816 1012 28868 1018
rect 28816 954 28868 960
rect 28828 800 28856 954
rect 28920 950 28948 2314
rect 29092 1148 29144 1154
rect 29092 1090 29144 1096
rect 28908 944 28960 950
rect 28908 886 28960 892
rect 29104 800 29132 1090
rect 29368 944 29420 950
rect 29368 886 29420 892
rect 29380 800 29408 886
rect 29656 800 29684 4014
rect 29748 3398 29776 5766
rect 29736 3392 29788 3398
rect 29736 3334 29788 3340
rect 29748 2922 29776 3334
rect 29736 2916 29788 2922
rect 29736 2858 29788 2864
rect 29932 2774 29960 6122
rect 30024 4554 30052 6870
rect 30012 4548 30064 4554
rect 30012 4490 30064 4496
rect 29840 2746 29960 2774
rect 29840 2310 29868 2746
rect 30024 2446 30052 4490
rect 30116 2922 30144 8758
rect 30208 7206 30236 11018
rect 30286 10160 30342 10169
rect 30286 10095 30342 10104
rect 30300 9994 30328 10095
rect 30288 9988 30340 9994
rect 30288 9930 30340 9936
rect 30392 9926 30420 13806
rect 30380 9920 30432 9926
rect 30380 9862 30432 9868
rect 30380 9716 30432 9722
rect 30380 9658 30432 9664
rect 30288 9580 30340 9586
rect 30288 9522 30340 9528
rect 30300 9382 30328 9522
rect 30392 9489 30420 9658
rect 30378 9480 30434 9489
rect 30378 9415 30434 9424
rect 30288 9376 30340 9382
rect 30288 9318 30340 9324
rect 30300 7954 30328 9318
rect 30484 7954 30512 17167
rect 30852 15162 30880 28970
rect 30932 20936 30984 20942
rect 30932 20878 30984 20884
rect 30944 19786 30972 20878
rect 31024 20596 31076 20602
rect 31024 20538 31076 20544
rect 31036 20058 31064 20538
rect 31128 20398 31156 37266
rect 31576 24268 31628 24274
rect 31576 24210 31628 24216
rect 31392 20936 31444 20942
rect 31392 20878 31444 20884
rect 31116 20392 31168 20398
rect 31404 20369 31432 20878
rect 31484 20392 31536 20398
rect 31116 20334 31168 20340
rect 31390 20360 31446 20369
rect 31024 20052 31076 20058
rect 31024 19994 31076 20000
rect 30932 19780 30984 19786
rect 30932 19722 30984 19728
rect 31036 17746 31064 19994
rect 31024 17740 31076 17746
rect 31024 17682 31076 17688
rect 31128 16250 31156 20334
rect 31484 20334 31536 20340
rect 31390 20295 31446 20304
rect 31404 19446 31432 20295
rect 31392 19440 31444 19446
rect 31392 19382 31444 19388
rect 31496 18834 31524 20334
rect 31392 18828 31444 18834
rect 31392 18770 31444 18776
rect 31484 18828 31536 18834
rect 31484 18770 31536 18776
rect 31404 18737 31432 18770
rect 31390 18728 31446 18737
rect 31390 18663 31446 18672
rect 31392 17536 31444 17542
rect 31392 17478 31444 17484
rect 31404 17202 31432 17478
rect 31392 17196 31444 17202
rect 31392 17138 31444 17144
rect 31206 16552 31262 16561
rect 31206 16487 31262 16496
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 31220 16182 31248 16487
rect 31300 16244 31352 16250
rect 31300 16186 31352 16192
rect 31208 16176 31260 16182
rect 31208 16118 31260 16124
rect 31220 15570 31248 16118
rect 31312 15978 31340 16186
rect 31300 15972 31352 15978
rect 31300 15914 31352 15920
rect 31208 15564 31260 15570
rect 31208 15506 31260 15512
rect 30840 15156 30892 15162
rect 30840 15098 30892 15104
rect 30564 15020 30616 15026
rect 30564 14962 30616 14968
rect 30576 13870 30604 14962
rect 30852 14074 30880 15098
rect 30932 15088 30984 15094
rect 30932 15030 30984 15036
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 30852 13870 30880 14010
rect 30564 13864 30616 13870
rect 30564 13806 30616 13812
rect 30840 13864 30892 13870
rect 30840 13806 30892 13812
rect 30944 13802 30972 15030
rect 31300 14340 31352 14346
rect 31300 14282 31352 14288
rect 31024 14272 31076 14278
rect 31024 14214 31076 14220
rect 31036 13938 31064 14214
rect 31312 14006 31340 14282
rect 31300 14000 31352 14006
rect 31300 13942 31352 13948
rect 31024 13932 31076 13938
rect 31076 13892 31248 13920
rect 31024 13874 31076 13880
rect 30932 13796 30984 13802
rect 30932 13738 30984 13744
rect 30840 13524 30892 13530
rect 30840 13466 30892 13472
rect 30748 12844 30800 12850
rect 30748 12786 30800 12792
rect 30760 12434 30788 12786
rect 30668 12406 30788 12434
rect 30668 11150 30696 12406
rect 30748 11756 30800 11762
rect 30748 11698 30800 11704
rect 30760 11558 30788 11698
rect 30748 11552 30800 11558
rect 30748 11494 30800 11500
rect 30656 11144 30708 11150
rect 30656 11086 30708 11092
rect 30656 11008 30708 11014
rect 30656 10950 30708 10956
rect 30668 10010 30696 10950
rect 30760 10130 30788 11494
rect 30748 10124 30800 10130
rect 30748 10066 30800 10072
rect 30668 9982 30788 10010
rect 30564 9920 30616 9926
rect 30564 9862 30616 9868
rect 30288 7948 30340 7954
rect 30288 7890 30340 7896
rect 30472 7948 30524 7954
rect 30472 7890 30524 7896
rect 30300 7834 30328 7890
rect 30300 7806 30420 7834
rect 30286 7712 30342 7721
rect 30286 7647 30342 7656
rect 30196 7200 30248 7206
rect 30196 7142 30248 7148
rect 30300 6730 30328 7647
rect 30392 6798 30420 7806
rect 30472 7812 30524 7818
rect 30472 7754 30524 7760
rect 30380 6792 30432 6798
rect 30380 6734 30432 6740
rect 30288 6724 30340 6730
rect 30288 6666 30340 6672
rect 30380 6180 30432 6186
rect 30380 6122 30432 6128
rect 30392 5914 30420 6122
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 30392 5710 30420 5850
rect 30380 5704 30432 5710
rect 30380 5646 30432 5652
rect 30288 4548 30340 4554
rect 30288 4490 30340 4496
rect 30300 3534 30328 4490
rect 30484 3670 30512 7754
rect 30472 3664 30524 3670
rect 30472 3606 30524 3612
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 30196 3460 30248 3466
rect 30196 3402 30248 3408
rect 30104 2916 30156 2922
rect 30104 2858 30156 2864
rect 30012 2440 30064 2446
rect 30012 2382 30064 2388
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 29828 2304 29880 2310
rect 29828 2246 29880 2252
rect 29932 800 29960 2314
rect 30208 800 30236 3402
rect 30576 2990 30604 9862
rect 30654 8936 30710 8945
rect 30654 8871 30710 8880
rect 30668 8838 30696 8871
rect 30656 8832 30708 8838
rect 30656 8774 30708 8780
rect 30656 7336 30708 7342
rect 30656 7278 30708 7284
rect 30668 7041 30696 7278
rect 30654 7032 30710 7041
rect 30654 6967 30710 6976
rect 30760 6934 30788 9982
rect 30852 8974 30880 13466
rect 30930 13424 30986 13433
rect 30930 13359 30986 13368
rect 30840 8968 30892 8974
rect 30840 8910 30892 8916
rect 30944 8566 30972 13359
rect 31116 12776 31168 12782
rect 31022 12744 31078 12753
rect 31116 12718 31168 12724
rect 31022 12679 31078 12688
rect 31036 12646 31064 12679
rect 31024 12640 31076 12646
rect 31024 12582 31076 12588
rect 31128 12374 31156 12718
rect 31024 12368 31076 12374
rect 31024 12310 31076 12316
rect 31116 12368 31168 12374
rect 31116 12310 31168 12316
rect 31036 10674 31064 12310
rect 31220 12238 31248 13892
rect 31404 13258 31432 17138
rect 31496 15094 31524 18770
rect 31484 15088 31536 15094
rect 31484 15030 31536 15036
rect 31588 13938 31616 24210
rect 31668 21072 31720 21078
rect 31668 21014 31720 21020
rect 31680 20806 31708 21014
rect 31668 20800 31720 20806
rect 31668 20742 31720 20748
rect 31666 20496 31722 20505
rect 31666 20431 31722 20440
rect 31680 19514 31708 20431
rect 31668 19508 31720 19514
rect 31668 19450 31720 19456
rect 31680 18766 31708 19450
rect 31668 18760 31720 18766
rect 31668 18702 31720 18708
rect 31772 16726 31800 43046
rect 32036 42628 32088 42634
rect 32036 42570 32088 42576
rect 31944 17672 31996 17678
rect 31944 17614 31996 17620
rect 31760 16720 31812 16726
rect 31760 16662 31812 16668
rect 31760 16108 31812 16114
rect 31760 16050 31812 16056
rect 31852 16108 31904 16114
rect 31852 16050 31904 16056
rect 31772 15502 31800 16050
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31760 14952 31812 14958
rect 31760 14894 31812 14900
rect 31772 14618 31800 14894
rect 31668 14612 31720 14618
rect 31668 14554 31720 14560
rect 31760 14612 31812 14618
rect 31760 14554 31812 14560
rect 31680 14498 31708 14554
rect 31864 14498 31892 16050
rect 31956 14929 31984 17614
rect 31942 14920 31998 14929
rect 31942 14855 31998 14864
rect 31944 14816 31996 14822
rect 31944 14758 31996 14764
rect 31680 14470 31892 14498
rect 31772 13938 31800 14470
rect 31850 14376 31906 14385
rect 31850 14311 31906 14320
rect 31576 13932 31628 13938
rect 31576 13874 31628 13880
rect 31760 13932 31812 13938
rect 31760 13874 31812 13880
rect 31864 13734 31892 14311
rect 31956 13938 31984 14758
rect 31944 13932 31996 13938
rect 31944 13874 31996 13880
rect 31852 13728 31904 13734
rect 31852 13670 31904 13676
rect 31864 13546 31892 13670
rect 31864 13518 31984 13546
rect 31956 13462 31984 13518
rect 31944 13456 31996 13462
rect 31944 13398 31996 13404
rect 31852 13388 31904 13394
rect 31772 13348 31852 13376
rect 31392 13252 31444 13258
rect 31392 13194 31444 13200
rect 31404 12238 31432 13194
rect 31484 12980 31536 12986
rect 31484 12922 31536 12928
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 31208 12232 31260 12238
rect 31208 12174 31260 12180
rect 31392 12232 31444 12238
rect 31392 12174 31444 12180
rect 31128 11898 31156 12174
rect 31300 12096 31352 12102
rect 31300 12038 31352 12044
rect 31116 11892 31168 11898
rect 31116 11834 31168 11840
rect 31208 11348 31260 11354
rect 31208 11290 31260 11296
rect 31024 10668 31076 10674
rect 31024 10610 31076 10616
rect 30932 8560 30984 8566
rect 30932 8502 30984 8508
rect 30840 8356 30892 8362
rect 30840 8298 30892 8304
rect 30748 6928 30800 6934
rect 30748 6870 30800 6876
rect 30852 6662 30880 8298
rect 31024 7404 31076 7410
rect 31024 7346 31076 7352
rect 30932 6860 30984 6866
rect 30932 6802 30984 6808
rect 30840 6656 30892 6662
rect 30840 6598 30892 6604
rect 30748 6112 30800 6118
rect 30748 6054 30800 6060
rect 30760 5846 30788 6054
rect 30748 5840 30800 5846
rect 30748 5782 30800 5788
rect 30852 5234 30880 6598
rect 30944 6322 30972 6802
rect 30932 6316 30984 6322
rect 30932 6258 30984 6264
rect 30840 5228 30892 5234
rect 30840 5170 30892 5176
rect 30746 4856 30802 4865
rect 30746 4791 30802 4800
rect 30760 4214 30788 4791
rect 30748 4208 30800 4214
rect 30748 4150 30800 4156
rect 30840 3936 30892 3942
rect 30840 3878 30892 3884
rect 30852 3058 30880 3878
rect 30944 3534 30972 6258
rect 31036 5914 31064 7346
rect 31116 7200 31168 7206
rect 31220 7177 31248 11290
rect 31312 11082 31340 12038
rect 31300 11076 31352 11082
rect 31300 11018 31352 11024
rect 31496 10520 31524 12922
rect 31576 12368 31628 12374
rect 31576 12310 31628 12316
rect 31588 12170 31616 12310
rect 31576 12164 31628 12170
rect 31576 12106 31628 12112
rect 31588 11830 31616 12106
rect 31576 11824 31628 11830
rect 31576 11766 31628 11772
rect 31668 11824 31720 11830
rect 31668 11766 31720 11772
rect 31680 11354 31708 11766
rect 31668 11348 31720 11354
rect 31668 11290 31720 11296
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 31312 10492 31524 10520
rect 31312 8634 31340 10492
rect 31680 9586 31708 11086
rect 31772 10742 31800 13348
rect 31852 13330 31904 13336
rect 31852 13252 31904 13258
rect 31852 13194 31904 13200
rect 31864 13161 31892 13194
rect 31944 13184 31996 13190
rect 31850 13152 31906 13161
rect 31944 13126 31996 13132
rect 31850 13087 31906 13096
rect 31956 11898 31984 13126
rect 31852 11892 31904 11898
rect 31852 11834 31904 11840
rect 31944 11892 31996 11898
rect 31944 11834 31996 11840
rect 31864 11150 31892 11834
rect 31942 11792 31998 11801
rect 31942 11727 31998 11736
rect 31852 11144 31904 11150
rect 31852 11086 31904 11092
rect 31760 10736 31812 10742
rect 31760 10678 31812 10684
rect 31760 10464 31812 10470
rect 31760 10406 31812 10412
rect 31668 9580 31720 9586
rect 31668 9522 31720 9528
rect 31484 9376 31536 9382
rect 31484 9318 31536 9324
rect 31392 9036 31444 9042
rect 31392 8978 31444 8984
rect 31404 8838 31432 8978
rect 31496 8974 31524 9318
rect 31574 9072 31630 9081
rect 31574 9007 31630 9016
rect 31680 9024 31708 9522
rect 31772 9466 31800 10406
rect 31852 10260 31904 10266
rect 31852 10202 31904 10208
rect 31864 9994 31892 10202
rect 31852 9988 31904 9994
rect 31852 9930 31904 9936
rect 31956 9518 31984 11727
rect 32048 11694 32076 42570
rect 32232 22094 32260 47534
rect 32312 43648 32364 43654
rect 32312 43590 32364 43596
rect 32324 43314 32352 43590
rect 32312 43308 32364 43314
rect 32312 43250 32364 43256
rect 32496 43308 32548 43314
rect 32496 43250 32548 43256
rect 32508 42770 32536 43250
rect 32496 42764 32548 42770
rect 32496 42706 32548 42712
rect 32600 24177 32628 60998
rect 32968 60110 32996 61202
rect 33244 61130 33272 63200
rect 33336 61198 33364 63242
rect 33966 63200 34022 63294
rect 34060 63242 34112 63248
rect 34702 63200 34758 64000
rect 35438 63322 35494 64000
rect 36174 63322 36230 64000
rect 36910 63322 36966 64000
rect 34796 63300 34848 63306
rect 34796 63242 34848 63248
rect 35438 63294 35940 63322
rect 33508 61668 33560 61674
rect 33508 61610 33560 61616
rect 33520 61198 33548 61610
rect 33324 61192 33376 61198
rect 33324 61134 33376 61140
rect 33508 61192 33560 61198
rect 33508 61134 33560 61140
rect 34716 61130 34744 63200
rect 34808 61198 34836 63242
rect 35438 63200 35494 63294
rect 34934 61500 35242 61509
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61435 35242 61444
rect 35912 61266 35940 63294
rect 36174 63294 36400 63322
rect 36174 63200 36230 63294
rect 35992 61396 36044 61402
rect 35992 61338 36044 61344
rect 36176 61396 36228 61402
rect 36176 61338 36228 61344
rect 35900 61260 35952 61266
rect 35900 61202 35952 61208
rect 34796 61192 34848 61198
rect 34796 61134 34848 61140
rect 36004 61130 36032 61338
rect 33232 61124 33284 61130
rect 33232 61066 33284 61072
rect 34704 61124 34756 61130
rect 34704 61066 34756 61072
rect 35900 61124 35952 61130
rect 35900 61066 35952 61072
rect 35992 61124 36044 61130
rect 35992 61066 36044 61072
rect 33508 61056 33560 61062
rect 33508 60998 33560 61004
rect 32956 60104 33008 60110
rect 32956 60046 33008 60052
rect 33048 59968 33100 59974
rect 33048 59910 33100 59916
rect 33060 56846 33088 59910
rect 33416 57044 33468 57050
rect 33416 56986 33468 56992
rect 33428 56846 33456 56986
rect 33048 56840 33100 56846
rect 33048 56782 33100 56788
rect 33416 56840 33468 56846
rect 33416 56782 33468 56788
rect 32680 56704 32732 56710
rect 32680 56646 32732 56652
rect 32692 50386 32720 56646
rect 33520 51074 33548 60998
rect 35716 60512 35768 60518
rect 35716 60454 35768 60460
rect 34934 60412 35242 60421
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60347 35242 60356
rect 34520 60104 34572 60110
rect 34520 60046 34572 60052
rect 34532 59634 34560 60046
rect 34520 59628 34572 59634
rect 34520 59570 34572 59576
rect 34532 58546 34560 59570
rect 34934 59324 35242 59333
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59259 35242 59268
rect 34520 58540 34572 58546
rect 34520 58482 34572 58488
rect 34934 58236 35242 58245
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58171 35242 58180
rect 35728 57934 35756 60454
rect 35808 58472 35860 58478
rect 35808 58414 35860 58420
rect 35820 58002 35848 58414
rect 35808 57996 35860 58002
rect 35808 57938 35860 57944
rect 35716 57928 35768 57934
rect 35716 57870 35768 57876
rect 34796 57860 34848 57866
rect 34796 57802 34848 57808
rect 33152 51046 33548 51074
rect 32680 50380 32732 50386
rect 32680 50322 32732 50328
rect 32680 43308 32732 43314
rect 32680 43250 32732 43256
rect 32692 42838 32720 43250
rect 32680 42832 32732 42838
rect 32678 42800 32680 42809
rect 32732 42800 32734 42809
rect 32678 42735 32734 42744
rect 33152 42702 33180 51046
rect 33232 50380 33284 50386
rect 33232 50322 33284 50328
rect 33048 42696 33100 42702
rect 33048 42638 33100 42644
rect 33140 42696 33192 42702
rect 33140 42638 33192 42644
rect 33060 42514 33088 42638
rect 33060 42486 33180 42514
rect 33152 42158 33180 42486
rect 33140 42152 33192 42158
rect 33140 42094 33192 42100
rect 33244 26234 33272 50322
rect 34520 47660 34572 47666
rect 34520 47602 34572 47608
rect 33784 45552 33836 45558
rect 33784 45494 33836 45500
rect 33796 43722 33824 45494
rect 34244 43920 34296 43926
rect 34244 43862 34296 43868
rect 34060 43784 34112 43790
rect 34060 43726 34112 43732
rect 33784 43716 33836 43722
rect 33784 43658 33836 43664
rect 33796 42770 33824 43658
rect 33784 42764 33836 42770
rect 33784 42706 33836 42712
rect 33876 42696 33928 42702
rect 33876 42638 33928 42644
rect 33888 42226 33916 42638
rect 33876 42220 33928 42226
rect 33876 42162 33928 42168
rect 34072 42158 34100 43726
rect 33784 42152 33836 42158
rect 33784 42094 33836 42100
rect 34060 42152 34112 42158
rect 34060 42094 34112 42100
rect 33508 39296 33560 39302
rect 33508 39238 33560 39244
rect 33520 37330 33548 39238
rect 33508 37324 33560 37330
rect 33508 37266 33560 37272
rect 33796 35494 33824 42094
rect 33784 35488 33836 35494
rect 33784 35430 33836 35436
rect 33784 29504 33836 29510
rect 33784 29446 33836 29452
rect 33152 26206 33272 26234
rect 32586 24168 32642 24177
rect 32586 24103 32642 24112
rect 32232 22066 32352 22094
rect 32220 18352 32272 18358
rect 32220 18294 32272 18300
rect 32232 18086 32260 18294
rect 32220 18080 32272 18086
rect 32220 18022 32272 18028
rect 32220 17128 32272 17134
rect 32220 17070 32272 17076
rect 32232 15910 32260 17070
rect 32324 16182 32352 22066
rect 32864 20324 32916 20330
rect 32864 20266 32916 20272
rect 32876 19922 32904 20266
rect 32864 19916 32916 19922
rect 32864 19858 32916 19864
rect 32496 19372 32548 19378
rect 32496 19314 32548 19320
rect 32402 18864 32458 18873
rect 32402 18799 32458 18808
rect 32416 18766 32444 18799
rect 32404 18760 32456 18766
rect 32404 18702 32456 18708
rect 32416 18358 32444 18702
rect 32404 18352 32456 18358
rect 32404 18294 32456 18300
rect 32404 18216 32456 18222
rect 32404 18158 32456 18164
rect 32416 17218 32444 18158
rect 32508 17746 32536 19314
rect 32588 18216 32640 18222
rect 32586 18184 32588 18193
rect 32680 18216 32732 18222
rect 32640 18184 32642 18193
rect 32680 18158 32732 18164
rect 32772 18216 32824 18222
rect 32772 18158 32824 18164
rect 32586 18119 32642 18128
rect 32692 18086 32720 18158
rect 32680 18080 32732 18086
rect 32680 18022 32732 18028
rect 32496 17740 32548 17746
rect 32496 17682 32548 17688
rect 32416 17190 32628 17218
rect 32600 17134 32628 17190
rect 32692 17134 32720 18022
rect 32784 17882 32812 18158
rect 32772 17876 32824 17882
rect 32772 17818 32824 17824
rect 32772 17536 32824 17542
rect 32772 17478 32824 17484
rect 32784 17202 32812 17478
rect 32876 17202 32904 19858
rect 32956 18692 33008 18698
rect 32956 18634 33008 18640
rect 32968 18290 32996 18634
rect 32956 18284 33008 18290
rect 32956 18226 33008 18232
rect 32772 17196 32824 17202
rect 32772 17138 32824 17144
rect 32864 17196 32916 17202
rect 32864 17138 32916 17144
rect 32588 17128 32640 17134
rect 32588 17070 32640 17076
rect 32680 17128 32732 17134
rect 32680 17070 32732 17076
rect 32404 16516 32456 16522
rect 32404 16458 32456 16464
rect 32312 16176 32364 16182
rect 32312 16118 32364 16124
rect 32220 15904 32272 15910
rect 32220 15846 32272 15852
rect 32128 15020 32180 15026
rect 32128 14962 32180 14968
rect 32140 14618 32168 14962
rect 32128 14612 32180 14618
rect 32128 14554 32180 14560
rect 32036 11688 32088 11694
rect 32036 11630 32088 11636
rect 32034 10432 32090 10441
rect 32034 10367 32090 10376
rect 32048 9722 32076 10367
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32140 9722 32168 9998
rect 32036 9716 32088 9722
rect 32036 9658 32088 9664
rect 32128 9716 32180 9722
rect 32128 9658 32180 9664
rect 31944 9512 31996 9518
rect 31772 9438 31892 9466
rect 31944 9454 31996 9460
rect 31864 9110 31892 9438
rect 32126 9208 32182 9217
rect 32126 9143 32182 9152
rect 31852 9104 31904 9110
rect 31852 9046 31904 9052
rect 31484 8968 31536 8974
rect 31484 8910 31536 8916
rect 31392 8832 31444 8838
rect 31392 8774 31444 8780
rect 31484 8832 31536 8838
rect 31588 8820 31616 9007
rect 31680 8996 31800 9024
rect 31668 8900 31720 8906
rect 31668 8842 31720 8848
rect 31536 8792 31616 8820
rect 31484 8774 31536 8780
rect 31496 8634 31524 8774
rect 31300 8628 31352 8634
rect 31300 8570 31352 8576
rect 31484 8628 31536 8634
rect 31484 8570 31536 8576
rect 31576 8492 31628 8498
rect 31576 8434 31628 8440
rect 31390 8256 31446 8265
rect 31390 8191 31446 8200
rect 31300 7472 31352 7478
rect 31300 7414 31352 7420
rect 31116 7142 31168 7148
rect 31206 7168 31262 7177
rect 31128 6322 31156 7142
rect 31206 7103 31262 7112
rect 31206 6760 31262 6769
rect 31206 6695 31208 6704
rect 31260 6695 31262 6704
rect 31208 6666 31260 6672
rect 31116 6316 31168 6322
rect 31116 6258 31168 6264
rect 31024 5908 31076 5914
rect 31024 5850 31076 5856
rect 31312 5778 31340 7414
rect 31404 6202 31432 8191
rect 31484 7336 31536 7342
rect 31484 7278 31536 7284
rect 31496 6934 31524 7278
rect 31484 6928 31536 6934
rect 31484 6870 31536 6876
rect 31404 6174 31524 6202
rect 31392 6112 31444 6118
rect 31392 6054 31444 6060
rect 31300 5772 31352 5778
rect 31300 5714 31352 5720
rect 31116 4208 31168 4214
rect 31116 4150 31168 4156
rect 30932 3528 30984 3534
rect 30932 3470 30984 3476
rect 31024 3392 31076 3398
rect 31024 3334 31076 3340
rect 31036 3233 31064 3334
rect 31022 3224 31078 3233
rect 31022 3159 31078 3168
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 30564 2984 30616 2990
rect 30564 2926 30616 2932
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 30472 2644 30524 2650
rect 30472 2586 30524 2592
rect 30288 2576 30340 2582
rect 30484 2530 30512 2586
rect 30340 2524 30512 2530
rect 30288 2518 30512 2524
rect 30300 2502 30512 2518
rect 30472 2372 30524 2378
rect 30472 2314 30524 2320
rect 30484 800 30512 2314
rect 30760 800 30788 2926
rect 31128 2446 31156 4150
rect 31312 3738 31340 5714
rect 31404 5710 31432 6054
rect 31392 5704 31444 5710
rect 31392 5646 31444 5652
rect 31496 4593 31524 6174
rect 31482 4584 31538 4593
rect 31482 4519 31538 4528
rect 31588 4026 31616 8434
rect 31680 8265 31708 8842
rect 31772 8362 31800 8996
rect 32140 8974 32168 9143
rect 31852 8968 31904 8974
rect 31852 8910 31904 8916
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 31864 8566 31892 8910
rect 31944 8628 31996 8634
rect 31944 8570 31996 8576
rect 31852 8560 31904 8566
rect 31852 8502 31904 8508
rect 31760 8356 31812 8362
rect 31760 8298 31812 8304
rect 31666 8256 31722 8265
rect 31666 8191 31722 8200
rect 31668 8084 31720 8090
rect 31668 8026 31720 8032
rect 31680 7886 31708 8026
rect 31668 7880 31720 7886
rect 31668 7822 31720 7828
rect 31668 7744 31720 7750
rect 31668 7686 31720 7692
rect 31680 7002 31708 7686
rect 31668 6996 31720 7002
rect 31668 6938 31720 6944
rect 31760 6724 31812 6730
rect 31760 6666 31812 6672
rect 31496 3998 31616 4026
rect 31496 3913 31524 3998
rect 31576 3936 31628 3942
rect 31482 3904 31538 3913
rect 31576 3878 31628 3884
rect 31482 3839 31538 3848
rect 31300 3732 31352 3738
rect 31300 3674 31352 3680
rect 31312 3602 31340 3674
rect 31300 3596 31352 3602
rect 31300 3538 31352 3544
rect 31312 3126 31340 3538
rect 31588 3534 31616 3878
rect 31772 3777 31800 6666
rect 31864 5234 31892 8502
rect 31956 6662 31984 8570
rect 31944 6656 31996 6662
rect 31944 6598 31996 6604
rect 31852 5228 31904 5234
rect 31852 5170 31904 5176
rect 32128 4004 32180 4010
rect 32128 3946 32180 3952
rect 31758 3768 31814 3777
rect 31758 3703 31814 3712
rect 31576 3528 31628 3534
rect 31576 3470 31628 3476
rect 31300 3120 31352 3126
rect 31300 3062 31352 3068
rect 31576 2984 31628 2990
rect 31576 2926 31628 2932
rect 31116 2440 31168 2446
rect 31116 2382 31168 2388
rect 31024 2372 31076 2378
rect 31024 2314 31076 2320
rect 31036 800 31064 2314
rect 31300 944 31352 950
rect 31300 886 31352 892
rect 31312 800 31340 886
rect 31588 800 31616 2926
rect 32140 2582 32168 3946
rect 32128 2576 32180 2582
rect 32128 2518 32180 2524
rect 32232 2310 32260 15846
rect 32312 15020 32364 15026
rect 32312 14962 32364 14968
rect 32324 12918 32352 14962
rect 32416 13326 32444 16458
rect 32496 16448 32548 16454
rect 32496 16390 32548 16396
rect 32508 14226 32536 16390
rect 32600 15994 32628 17070
rect 32772 16720 32824 16726
rect 32772 16662 32824 16668
rect 32600 15966 32720 15994
rect 32692 15502 32720 15966
rect 32680 15496 32732 15502
rect 32680 15438 32732 15444
rect 32692 15042 32720 15438
rect 32600 15014 32720 15042
rect 32600 14346 32628 15014
rect 32680 14816 32732 14822
rect 32680 14758 32732 14764
rect 32692 14414 32720 14758
rect 32680 14408 32732 14414
rect 32680 14350 32732 14356
rect 32588 14340 32640 14346
rect 32588 14282 32640 14288
rect 32508 14198 32720 14226
rect 32496 13932 32548 13938
rect 32496 13874 32548 13880
rect 32404 13320 32456 13326
rect 32404 13262 32456 13268
rect 32312 12912 32364 12918
rect 32312 12854 32364 12860
rect 32404 12776 32456 12782
rect 32404 12718 32456 12724
rect 32416 12434 32444 12718
rect 32508 12714 32536 13874
rect 32586 13560 32642 13569
rect 32586 13495 32588 13504
rect 32640 13495 32642 13504
rect 32588 13466 32640 13472
rect 32588 13184 32640 13190
rect 32588 13126 32640 13132
rect 32600 12850 32628 13126
rect 32588 12844 32640 12850
rect 32588 12786 32640 12792
rect 32496 12708 32548 12714
rect 32496 12650 32548 12656
rect 32416 12406 32536 12434
rect 32312 11892 32364 11898
rect 32312 11834 32364 11840
rect 32324 10470 32352 11834
rect 32508 11286 32536 12406
rect 32404 11280 32456 11286
rect 32404 11222 32456 11228
rect 32496 11280 32548 11286
rect 32496 11222 32548 11228
rect 32312 10464 32364 10470
rect 32312 10406 32364 10412
rect 32416 10062 32444 11222
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32404 10056 32456 10062
rect 32404 9998 32456 10004
rect 32508 9994 32536 11086
rect 32692 10606 32720 14198
rect 32784 12850 32812 16662
rect 32876 16658 32904 17138
rect 32864 16652 32916 16658
rect 32864 16594 32916 16600
rect 32876 15026 32904 16594
rect 32956 15972 33008 15978
rect 32956 15914 33008 15920
rect 32968 15162 32996 15914
rect 32956 15156 33008 15162
rect 33008 15116 33088 15144
rect 32956 15098 33008 15104
rect 32864 15020 32916 15026
rect 32864 14962 32916 14968
rect 32956 14544 33008 14550
rect 32956 14486 33008 14492
rect 32968 14414 32996 14486
rect 32956 14408 33008 14414
rect 32956 14350 33008 14356
rect 32864 14340 32916 14346
rect 32864 14282 32916 14288
rect 32876 14074 32904 14282
rect 32864 14068 32916 14074
rect 32864 14010 32916 14016
rect 33060 13326 33088 15116
rect 33048 13320 33100 13326
rect 33048 13262 33100 13268
rect 32772 12844 32824 12850
rect 32772 12786 32824 12792
rect 33060 12782 33088 13262
rect 33048 12776 33100 12782
rect 33048 12718 33100 12724
rect 32772 12368 32824 12374
rect 32772 12310 32824 12316
rect 32588 10600 32640 10606
rect 32588 10542 32640 10548
rect 32680 10600 32732 10606
rect 32680 10542 32732 10548
rect 32496 9988 32548 9994
rect 32496 9930 32548 9936
rect 32312 9920 32364 9926
rect 32312 9862 32364 9868
rect 32324 8294 32352 9862
rect 32404 8900 32456 8906
rect 32404 8842 32456 8848
rect 32416 8809 32444 8842
rect 32402 8800 32458 8809
rect 32402 8735 32458 8744
rect 32312 8288 32364 8294
rect 32312 8230 32364 8236
rect 32508 2446 32536 9930
rect 32600 9586 32628 10542
rect 32784 10452 32812 12310
rect 32864 12096 32916 12102
rect 32864 12038 32916 12044
rect 32876 11762 32904 12038
rect 33152 11762 33180 26206
rect 33796 23050 33824 29446
rect 34256 27606 34284 43862
rect 34244 27600 34296 27606
rect 34244 27542 34296 27548
rect 34060 25832 34112 25838
rect 34060 25774 34112 25780
rect 33784 23044 33836 23050
rect 33784 22986 33836 22992
rect 33784 22772 33836 22778
rect 33784 22714 33836 22720
rect 33324 21344 33376 21350
rect 33324 21286 33376 21292
rect 33336 20398 33364 21286
rect 33796 20641 33824 22714
rect 33782 20632 33838 20641
rect 33782 20567 33838 20576
rect 33416 20460 33468 20466
rect 33416 20402 33468 20408
rect 33600 20460 33652 20466
rect 33600 20402 33652 20408
rect 33324 20392 33376 20398
rect 33324 20334 33376 20340
rect 33232 17536 33284 17542
rect 33232 17478 33284 17484
rect 33244 16590 33272 17478
rect 33232 16584 33284 16590
rect 33232 16526 33284 16532
rect 33232 12776 33284 12782
rect 33232 12718 33284 12724
rect 32864 11756 32916 11762
rect 32864 11698 32916 11704
rect 32956 11756 33008 11762
rect 32956 11698 33008 11704
rect 33140 11756 33192 11762
rect 33140 11698 33192 11704
rect 32864 11076 32916 11082
rect 32864 11018 32916 11024
rect 32692 10424 32812 10452
rect 32588 9580 32640 9586
rect 32588 9522 32640 9528
rect 32600 8974 32628 9522
rect 32588 8968 32640 8974
rect 32588 8910 32640 8916
rect 32692 8906 32720 10424
rect 32772 9580 32824 9586
rect 32772 9522 32824 9528
rect 32680 8900 32732 8906
rect 32680 8842 32732 8848
rect 32588 6724 32640 6730
rect 32588 6666 32640 6672
rect 32600 4078 32628 6666
rect 32784 5914 32812 9522
rect 32876 8809 32904 11018
rect 32968 10810 32996 11698
rect 33140 11280 33192 11286
rect 33140 11222 33192 11228
rect 33048 11144 33100 11150
rect 33048 11086 33100 11092
rect 32956 10804 33008 10810
rect 32956 10746 33008 10752
rect 33060 10554 33088 11086
rect 33152 10674 33180 11222
rect 33140 10668 33192 10674
rect 33140 10610 33192 10616
rect 33060 10526 33180 10554
rect 33152 9722 33180 10526
rect 33140 9716 33192 9722
rect 33140 9658 33192 9664
rect 33244 9568 33272 12718
rect 33336 11082 33364 20334
rect 33428 19514 33456 20402
rect 33612 19854 33640 20402
rect 33600 19848 33652 19854
rect 33600 19790 33652 19796
rect 33416 19508 33468 19514
rect 33416 19450 33468 19456
rect 33796 17678 33824 20567
rect 33968 19712 34020 19718
rect 33968 19654 34020 19660
rect 33980 19514 34008 19654
rect 34072 19514 34100 25774
rect 34532 22094 34560 47602
rect 34704 44192 34756 44198
rect 34704 44134 34756 44140
rect 34716 33590 34744 44134
rect 34704 33584 34756 33590
rect 34704 33526 34756 33532
rect 34808 30802 34836 57802
rect 35440 57792 35492 57798
rect 35440 57734 35492 57740
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 35452 45082 35480 57734
rect 35440 45076 35492 45082
rect 35440 45018 35492 45024
rect 35256 45008 35308 45014
rect 35256 44950 35308 44956
rect 35268 44878 35296 44950
rect 35072 44872 35124 44878
rect 35072 44814 35124 44820
rect 35256 44872 35308 44878
rect 35256 44814 35308 44820
rect 35084 44198 35112 44814
rect 35072 44192 35124 44198
rect 35072 44134 35124 44140
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 35912 43722 35940 61066
rect 36084 61056 36136 61062
rect 36084 60998 36136 61004
rect 35900 43716 35952 43722
rect 35900 43658 35952 43664
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35900 33856 35952 33862
rect 35900 33798 35952 33804
rect 35912 33522 35940 33798
rect 36096 33590 36124 60998
rect 36188 60858 36216 61338
rect 36176 60852 36228 60858
rect 36176 60794 36228 60800
rect 36372 60790 36400 63294
rect 36910 63294 37320 63322
rect 36910 63200 36966 63294
rect 37292 61198 37320 63294
rect 37646 63200 37702 64000
rect 38382 63322 38438 64000
rect 39118 63322 39174 64000
rect 39854 63322 39910 64000
rect 40590 63322 40646 64000
rect 41326 63322 41382 64000
rect 38382 63294 38792 63322
rect 38382 63200 38438 63294
rect 37660 61198 37688 63200
rect 38764 61198 38792 63294
rect 39118 63306 39252 63322
rect 39118 63300 39264 63306
rect 39118 63294 39212 63300
rect 39118 63200 39174 63294
rect 39212 63242 39264 63248
rect 39854 63294 40080 63322
rect 40590 63306 40724 63322
rect 39854 63200 39910 63294
rect 37280 61192 37332 61198
rect 37280 61134 37332 61140
rect 37648 61192 37700 61198
rect 37648 61134 37700 61140
rect 38752 61192 38804 61198
rect 38752 61134 38804 61140
rect 40052 61130 40080 63294
rect 40132 63300 40184 63306
rect 40132 63242 40184 63248
rect 40590 63300 40736 63306
rect 40590 63294 40684 63300
rect 40144 61198 40172 63242
rect 40590 63200 40646 63294
rect 40684 63242 40736 63248
rect 41326 63294 41552 63322
rect 41326 63200 41382 63294
rect 40132 61192 40184 61198
rect 40132 61134 40184 61140
rect 38200 61124 38252 61130
rect 38200 61066 38252 61072
rect 40040 61124 40092 61130
rect 40040 61066 40092 61072
rect 41420 61124 41472 61130
rect 41420 61066 41472 61072
rect 36360 60784 36412 60790
rect 36360 60726 36412 60732
rect 38212 58546 38240 61066
rect 39120 61056 39172 61062
rect 39120 60998 39172 61004
rect 40224 61056 40276 61062
rect 40224 60998 40276 61004
rect 40316 61056 40368 61062
rect 40316 60998 40368 61004
rect 38844 59152 38896 59158
rect 38844 59094 38896 59100
rect 38856 58546 38884 59094
rect 37924 58540 37976 58546
rect 37924 58482 37976 58488
rect 38200 58540 38252 58546
rect 38200 58482 38252 58488
rect 38292 58540 38344 58546
rect 38292 58482 38344 58488
rect 38476 58540 38528 58546
rect 38476 58482 38528 58488
rect 38844 58540 38896 58546
rect 38844 58482 38896 58488
rect 36912 58404 36964 58410
rect 36912 58346 36964 58352
rect 36268 57928 36320 57934
rect 36268 57870 36320 57876
rect 36280 56982 36308 57870
rect 36268 56976 36320 56982
rect 36268 56918 36320 56924
rect 36544 50380 36596 50386
rect 36544 50322 36596 50328
rect 36360 46368 36412 46374
rect 36360 46310 36412 46316
rect 36372 45490 36400 46310
rect 36360 45484 36412 45490
rect 36360 45426 36412 45432
rect 36556 33862 36584 50322
rect 36636 45484 36688 45490
rect 36636 45426 36688 45432
rect 36544 33856 36596 33862
rect 36544 33798 36596 33804
rect 36084 33584 36136 33590
rect 36084 33526 36136 33532
rect 35900 33516 35952 33522
rect 35900 33458 35952 33464
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 36360 31136 36412 31142
rect 36360 31078 36412 31084
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34796 30796 34848 30802
rect 34796 30738 34848 30744
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35440 27600 35492 27606
rect 35440 27542 35492 27548
rect 34612 27328 34664 27334
rect 34612 27270 34664 27276
rect 34624 23526 34652 27270
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34612 23520 34664 23526
rect 34612 23462 34664 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34532 22066 34652 22094
rect 34334 19816 34390 19825
rect 34334 19751 34390 19760
rect 34348 19718 34376 19751
rect 34336 19712 34388 19718
rect 34336 19654 34388 19660
rect 33968 19508 34020 19514
rect 33968 19450 34020 19456
rect 34060 19508 34112 19514
rect 34060 19450 34112 19456
rect 33980 19378 34008 19450
rect 33968 19372 34020 19378
rect 33968 19314 34020 19320
rect 34072 18358 34100 19450
rect 34060 18352 34112 18358
rect 34060 18294 34112 18300
rect 33876 18216 33928 18222
rect 33876 18158 33928 18164
rect 33888 17746 33916 18158
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 33876 17740 33928 17746
rect 33876 17682 33928 17688
rect 33784 17672 33836 17678
rect 33784 17614 33836 17620
rect 33692 17604 33744 17610
rect 33692 17546 33744 17552
rect 33704 17270 33732 17546
rect 33876 17536 33928 17542
rect 33876 17478 33928 17484
rect 33692 17264 33744 17270
rect 33692 17206 33744 17212
rect 33416 17128 33468 17134
rect 33416 17070 33468 17076
rect 33508 17128 33560 17134
rect 33508 17070 33560 17076
rect 33428 11354 33456 17070
rect 33520 16998 33548 17070
rect 33508 16992 33560 16998
rect 33508 16934 33560 16940
rect 33888 16538 33916 17478
rect 33980 17270 34008 18022
rect 34060 17740 34112 17746
rect 34060 17682 34112 17688
rect 33968 17264 34020 17270
rect 33968 17206 34020 17212
rect 33888 16510 34008 16538
rect 33980 16454 34008 16510
rect 33968 16448 34020 16454
rect 33968 16390 34020 16396
rect 33600 14612 33652 14618
rect 33600 14554 33652 14560
rect 33612 14414 33640 14554
rect 33600 14408 33652 14414
rect 33600 14350 33652 14356
rect 33508 13728 33560 13734
rect 33508 13670 33560 13676
rect 33416 11348 33468 11354
rect 33416 11290 33468 11296
rect 33520 11150 33548 13670
rect 33600 13456 33652 13462
rect 33600 13398 33652 13404
rect 33612 12434 33640 13398
rect 33784 12844 33836 12850
rect 33784 12786 33836 12792
rect 33612 12406 33732 12434
rect 33600 11824 33652 11830
rect 33600 11766 33652 11772
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 33324 11076 33376 11082
rect 33324 11018 33376 11024
rect 33324 10668 33376 10674
rect 33324 10610 33376 10616
rect 33416 10668 33468 10674
rect 33416 10610 33468 10616
rect 33508 10668 33560 10674
rect 33508 10610 33560 10616
rect 33336 9722 33364 10610
rect 33428 10441 33456 10610
rect 33414 10432 33470 10441
rect 33414 10367 33470 10376
rect 33324 9716 33376 9722
rect 33324 9658 33376 9664
rect 33060 9540 33272 9568
rect 33416 9580 33468 9586
rect 32956 9376 33008 9382
rect 32956 9318 33008 9324
rect 32968 9110 32996 9318
rect 32956 9104 33008 9110
rect 32956 9046 33008 9052
rect 32862 8800 32918 8809
rect 32862 8735 32918 8744
rect 32876 8634 32904 8735
rect 32864 8628 32916 8634
rect 32864 8570 32916 8576
rect 33060 8537 33088 9540
rect 33416 9522 33468 9528
rect 33140 9104 33192 9110
rect 33140 9046 33192 9052
rect 33046 8528 33102 8537
rect 32864 8492 32916 8498
rect 33046 8463 33048 8472
rect 32864 8434 32916 8440
rect 33100 8463 33102 8472
rect 33048 8434 33100 8440
rect 32876 8090 32904 8434
rect 32864 8084 32916 8090
rect 32864 8026 32916 8032
rect 32772 5908 32824 5914
rect 32772 5850 32824 5856
rect 32876 5370 32904 8026
rect 33152 7818 33180 9046
rect 33428 8974 33456 9522
rect 33520 9081 33548 10610
rect 33612 10266 33640 11766
rect 33600 10260 33652 10266
rect 33600 10202 33652 10208
rect 33600 10056 33652 10062
rect 33600 9998 33652 10004
rect 33506 9072 33562 9081
rect 33506 9007 33562 9016
rect 33416 8968 33468 8974
rect 33416 8910 33468 8916
rect 33232 8832 33284 8838
rect 33232 8774 33284 8780
rect 33244 7886 33272 8774
rect 33324 8628 33376 8634
rect 33324 8570 33376 8576
rect 33232 7880 33284 7886
rect 33232 7822 33284 7828
rect 33140 7812 33192 7818
rect 33140 7754 33192 7760
rect 33048 7744 33100 7750
rect 33048 7686 33100 7692
rect 33060 6458 33088 7686
rect 33140 6656 33192 6662
rect 33140 6598 33192 6604
rect 33152 6458 33180 6598
rect 33048 6452 33100 6458
rect 33048 6394 33100 6400
rect 33140 6452 33192 6458
rect 33140 6394 33192 6400
rect 32956 6112 33008 6118
rect 32956 6054 33008 6060
rect 32864 5364 32916 5370
rect 32864 5306 32916 5312
rect 32968 5001 32996 6054
rect 33048 5908 33100 5914
rect 33048 5850 33100 5856
rect 32954 4992 33010 5001
rect 32954 4927 33010 4936
rect 32864 4684 32916 4690
rect 32864 4626 32916 4632
rect 32876 4078 32904 4626
rect 32968 4622 32996 4927
rect 32956 4616 33008 4622
rect 32956 4558 33008 4564
rect 33060 4185 33088 5850
rect 33336 5681 33364 8570
rect 33428 7886 33456 8910
rect 33416 7880 33468 7886
rect 33416 7822 33468 7828
rect 33612 7721 33640 9998
rect 33598 7712 33654 7721
rect 33598 7647 33654 7656
rect 33704 6798 33732 12406
rect 33796 12306 33824 12786
rect 33784 12300 33836 12306
rect 33784 12242 33836 12248
rect 33796 11762 33824 12242
rect 33784 11756 33836 11762
rect 33784 11698 33836 11704
rect 33784 11076 33836 11082
rect 33784 11018 33836 11024
rect 33796 6866 33824 11018
rect 33876 10668 33928 10674
rect 33876 10610 33928 10616
rect 33888 10062 33916 10610
rect 33876 10056 33928 10062
rect 33876 9998 33928 10004
rect 33876 9172 33928 9178
rect 33980 9160 34008 16390
rect 34072 16289 34100 17682
rect 34426 17096 34482 17105
rect 34426 17031 34482 17040
rect 34058 16280 34114 16289
rect 34058 16215 34114 16224
rect 34060 15564 34112 15570
rect 34060 15506 34112 15512
rect 33928 9132 34008 9160
rect 33876 9114 33928 9120
rect 33968 8900 34020 8906
rect 33968 8842 34020 8848
rect 33980 8809 34008 8842
rect 33966 8800 34022 8809
rect 33888 8758 33966 8786
rect 33888 8498 33916 8758
rect 33966 8735 34022 8744
rect 33876 8492 33928 8498
rect 33876 8434 33928 8440
rect 33968 8492 34020 8498
rect 33968 8434 34020 8440
rect 33980 8090 34008 8434
rect 33968 8084 34020 8090
rect 33968 8026 34020 8032
rect 33784 6860 33836 6866
rect 33784 6802 33836 6808
rect 33692 6792 33744 6798
rect 33692 6734 33744 6740
rect 33796 6390 33824 6802
rect 33784 6384 33836 6390
rect 33784 6326 33836 6332
rect 33322 5672 33378 5681
rect 33322 5607 33378 5616
rect 33140 5092 33192 5098
rect 33140 5034 33192 5040
rect 33152 4554 33180 5034
rect 33140 4548 33192 4554
rect 33140 4490 33192 4496
rect 33336 4282 33364 5607
rect 33508 4820 33560 4826
rect 33508 4762 33560 4768
rect 33520 4486 33548 4762
rect 33796 4554 33824 6326
rect 34072 5710 34100 15506
rect 34440 15162 34468 17031
rect 34428 15156 34480 15162
rect 34428 15098 34480 15104
rect 34520 13728 34572 13734
rect 34520 13670 34572 13676
rect 34532 12918 34560 13670
rect 34520 12912 34572 12918
rect 34520 12854 34572 12860
rect 34336 12164 34388 12170
rect 34336 12106 34388 12112
rect 34152 11348 34204 11354
rect 34152 11290 34204 11296
rect 34164 9625 34192 11290
rect 34348 10810 34376 12106
rect 34518 11248 34574 11257
rect 34518 11183 34574 11192
rect 34428 11076 34480 11082
rect 34428 11018 34480 11024
rect 34336 10804 34388 10810
rect 34336 10746 34388 10752
rect 34244 10668 34296 10674
rect 34244 10610 34296 10616
rect 34256 10266 34284 10610
rect 34348 10441 34376 10746
rect 34334 10432 34390 10441
rect 34334 10367 34390 10376
rect 34244 10260 34296 10266
rect 34244 10202 34296 10208
rect 34440 10198 34468 11018
rect 34428 10192 34480 10198
rect 34428 10134 34480 10140
rect 34336 9648 34388 9654
rect 34150 9616 34206 9625
rect 34336 9590 34388 9596
rect 34150 9551 34206 9560
rect 34244 9512 34296 9518
rect 34244 9454 34296 9460
rect 34256 8974 34284 9454
rect 34152 8968 34204 8974
rect 34150 8936 34152 8945
rect 34244 8968 34296 8974
rect 34204 8936 34206 8945
rect 34244 8910 34296 8916
rect 34150 8871 34206 8880
rect 34348 8498 34376 9590
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 34336 8492 34388 8498
rect 34336 8434 34388 8440
rect 34164 8401 34192 8434
rect 34150 8392 34206 8401
rect 34150 8327 34206 8336
rect 34336 8356 34388 8362
rect 34336 8298 34388 8304
rect 34060 5704 34112 5710
rect 34060 5646 34112 5652
rect 34072 4554 34100 5646
rect 34244 5568 34296 5574
rect 34244 5510 34296 5516
rect 34256 5234 34284 5510
rect 34244 5228 34296 5234
rect 34244 5170 34296 5176
rect 34348 5098 34376 8298
rect 34532 7750 34560 11183
rect 34624 10810 34652 22066
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 34808 20942 34836 21490
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 20936 34848 20942
rect 34796 20878 34848 20884
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35348 18216 35400 18222
rect 35348 18158 35400 18164
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34796 17672 34848 17678
rect 34796 17614 34848 17620
rect 34808 16998 34836 17614
rect 34796 16992 34848 16998
rect 34796 16934 34848 16940
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35360 15570 35388 18158
rect 35348 15564 35400 15570
rect 35348 15506 35400 15512
rect 34704 15360 34756 15366
rect 34704 15302 34756 15308
rect 34716 15026 34744 15302
rect 34704 15020 34756 15026
rect 34704 14962 34756 14968
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34704 14000 34756 14006
rect 34704 13942 34756 13948
rect 34612 10804 34664 10810
rect 34612 10746 34664 10752
rect 34716 9674 34744 13942
rect 35360 13870 35388 15506
rect 34796 13864 34848 13870
rect 34796 13806 34848 13812
rect 35348 13864 35400 13870
rect 35348 13806 35400 13812
rect 34808 12986 34836 13806
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34796 12980 34848 12986
rect 34796 12922 34848 12928
rect 35256 12980 35308 12986
rect 35256 12922 35308 12928
rect 34796 12844 34848 12850
rect 34796 12786 34848 12792
rect 34808 11121 34836 12786
rect 35268 12753 35296 12922
rect 35254 12744 35310 12753
rect 35254 12679 35310 12688
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35348 12232 35400 12238
rect 35348 12174 35400 12180
rect 35360 11898 35388 12174
rect 35348 11892 35400 11898
rect 35348 11834 35400 11840
rect 35348 11756 35400 11762
rect 35348 11698 35400 11704
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35360 11354 35388 11698
rect 35348 11348 35400 11354
rect 35348 11290 35400 11296
rect 34794 11112 34850 11121
rect 34794 11047 34850 11056
rect 35348 10804 35400 10810
rect 35348 10746 35400 10752
rect 35164 10668 35216 10674
rect 35164 10610 35216 10616
rect 35176 10470 35204 10610
rect 35164 10464 35216 10470
rect 35164 10406 35216 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35256 9988 35308 9994
rect 35256 9930 35308 9936
rect 35268 9897 35296 9930
rect 35254 9888 35310 9897
rect 35254 9823 35310 9832
rect 34716 9646 34836 9674
rect 34808 9500 34836 9646
rect 34716 9472 34836 9500
rect 34520 7744 34572 7750
rect 34520 7686 34572 7692
rect 34428 7404 34480 7410
rect 34428 7346 34480 7352
rect 34440 7002 34468 7346
rect 34428 6996 34480 7002
rect 34428 6938 34480 6944
rect 34532 6322 34560 7686
rect 34520 6316 34572 6322
rect 34520 6258 34572 6264
rect 34428 5228 34480 5234
rect 34428 5170 34480 5176
rect 34336 5092 34388 5098
rect 34336 5034 34388 5040
rect 33784 4548 33836 4554
rect 33784 4490 33836 4496
rect 34060 4548 34112 4554
rect 34060 4490 34112 4496
rect 33508 4480 33560 4486
rect 33508 4422 33560 4428
rect 33600 4480 33652 4486
rect 33600 4422 33652 4428
rect 33324 4276 33376 4282
rect 33324 4218 33376 4224
rect 33046 4176 33102 4185
rect 33046 4111 33102 4120
rect 32588 4072 32640 4078
rect 32588 4014 32640 4020
rect 32864 4072 32916 4078
rect 32864 4014 32916 4020
rect 33140 4072 33192 4078
rect 33140 4014 33192 4020
rect 32600 3398 32628 4014
rect 33152 3890 33180 4014
rect 32692 3862 33180 3890
rect 32588 3392 32640 3398
rect 32588 3334 32640 3340
rect 32496 2440 32548 2446
rect 32496 2382 32548 2388
rect 32588 2372 32640 2378
rect 32588 2314 32640 2320
rect 32220 2304 32272 2310
rect 32220 2246 32272 2252
rect 32404 1216 32456 1222
rect 32404 1158 32456 1164
rect 32128 1080 32180 1086
rect 32128 1022 32180 1028
rect 31852 1012 31904 1018
rect 31852 954 31904 960
rect 31864 800 31892 954
rect 32140 800 32168 1022
rect 32416 800 32444 1158
rect 32600 950 32628 2314
rect 32588 944 32640 950
rect 32588 886 32640 892
rect 32692 800 32720 3862
rect 33336 3738 33364 4218
rect 33324 3732 33376 3738
rect 33324 3674 33376 3680
rect 33416 3596 33468 3602
rect 33416 3538 33468 3544
rect 33232 3460 33284 3466
rect 33232 3402 33284 3408
rect 32956 944 33008 950
rect 32956 886 33008 892
rect 32968 800 32996 886
rect 33244 800 33272 3402
rect 33428 898 33456 3538
rect 33612 2990 33640 4422
rect 34244 4276 34296 4282
rect 34244 4218 34296 4224
rect 34256 3194 34284 4218
rect 34348 3194 34376 5034
rect 34440 4554 34468 5170
rect 34612 5092 34664 5098
rect 34612 5034 34664 5040
rect 34520 4616 34572 4622
rect 34520 4558 34572 4564
rect 34428 4548 34480 4554
rect 34428 4490 34480 4496
rect 34244 3188 34296 3194
rect 34244 3130 34296 3136
rect 34336 3188 34388 3194
rect 34336 3130 34388 3136
rect 34532 3058 34560 4558
rect 34624 4214 34652 5034
rect 34612 4208 34664 4214
rect 34716 4185 34744 9472
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35360 7886 35388 10746
rect 35452 10674 35480 27542
rect 36176 24268 36228 24274
rect 36176 24210 36228 24216
rect 35532 24200 35584 24206
rect 35532 24142 35584 24148
rect 35544 12238 35572 24142
rect 35624 20936 35676 20942
rect 35624 20878 35676 20884
rect 35636 15502 35664 20878
rect 35716 20800 35768 20806
rect 35716 20742 35768 20748
rect 35992 20800 36044 20806
rect 35992 20742 36044 20748
rect 35728 20534 35756 20742
rect 35716 20528 35768 20534
rect 35716 20470 35768 20476
rect 35900 20460 35952 20466
rect 35900 20402 35952 20408
rect 35912 19514 35940 20402
rect 36004 20262 36032 20742
rect 36084 20528 36136 20534
rect 36084 20470 36136 20476
rect 35992 20256 36044 20262
rect 35992 20198 36044 20204
rect 36096 19786 36124 20470
rect 36084 19780 36136 19786
rect 36084 19722 36136 19728
rect 36188 19718 36216 24210
rect 36176 19712 36228 19718
rect 36176 19654 36228 19660
rect 36268 19712 36320 19718
rect 36268 19654 36320 19660
rect 35900 19508 35952 19514
rect 35900 19450 35952 19456
rect 36188 16522 36216 19654
rect 36280 19446 36308 19654
rect 36268 19440 36320 19446
rect 36268 19382 36320 19388
rect 36372 19378 36400 31078
rect 36648 22166 36676 45426
rect 36924 45354 36952 58346
rect 37936 58342 37964 58482
rect 38304 58410 38332 58482
rect 38292 58404 38344 58410
rect 38292 58346 38344 58352
rect 37556 58336 37608 58342
rect 37556 58278 37608 58284
rect 37924 58336 37976 58342
rect 37924 58278 37976 58284
rect 37372 45484 37424 45490
rect 37372 45426 37424 45432
rect 36912 45348 36964 45354
rect 36912 45290 36964 45296
rect 37280 42696 37332 42702
rect 37280 42638 37332 42644
rect 37292 42362 37320 42638
rect 37384 42634 37412 45426
rect 37372 42628 37424 42634
rect 37372 42570 37424 42576
rect 37280 42356 37332 42362
rect 37280 42298 37332 42304
rect 37384 35290 37412 42570
rect 37372 35284 37424 35290
rect 37372 35226 37424 35232
rect 37384 35018 37412 35226
rect 37372 35012 37424 35018
rect 37372 34954 37424 34960
rect 37568 32434 37596 58278
rect 38488 45490 38516 58482
rect 38016 45484 38068 45490
rect 38016 45426 38068 45432
rect 38476 45484 38528 45490
rect 38476 45426 38528 45432
rect 37832 33312 37884 33318
rect 37832 33254 37884 33260
rect 37556 32428 37608 32434
rect 37556 32370 37608 32376
rect 36636 22160 36688 22166
rect 36636 22102 36688 22108
rect 37844 22094 37872 33254
rect 37752 22066 37872 22094
rect 38028 22094 38056 45426
rect 38488 33658 38516 45426
rect 39132 36650 39160 60998
rect 40236 60858 40264 60998
rect 40224 60852 40276 60858
rect 40224 60794 40276 60800
rect 40040 58472 40092 58478
rect 40040 58414 40092 58420
rect 40052 55758 40080 58414
rect 40040 55752 40092 55758
rect 40040 55694 40092 55700
rect 40132 53712 40184 53718
rect 40132 53654 40184 53660
rect 39304 42560 39356 42566
rect 39304 42502 39356 42508
rect 39120 36644 39172 36650
rect 39120 36586 39172 36592
rect 38476 33652 38528 33658
rect 38476 33594 38528 33600
rect 39316 25838 39344 42502
rect 39396 42356 39448 42362
rect 39396 42298 39448 42304
rect 39304 25832 39356 25838
rect 39304 25774 39356 25780
rect 38844 24608 38896 24614
rect 38844 24550 38896 24556
rect 38856 22094 38884 24550
rect 38028 22066 38148 22094
rect 38856 22066 39068 22094
rect 36544 21004 36596 21010
rect 36544 20946 36596 20952
rect 36360 19372 36412 19378
rect 36360 19314 36412 19320
rect 35808 16516 35860 16522
rect 35808 16458 35860 16464
rect 36176 16516 36228 16522
rect 36176 16458 36228 16464
rect 35820 16114 35848 16458
rect 36268 16448 36320 16454
rect 36268 16390 36320 16396
rect 35808 16108 35860 16114
rect 35808 16050 35860 16056
rect 36280 15570 36308 16390
rect 36268 15564 36320 15570
rect 36268 15506 36320 15512
rect 35624 15496 35676 15502
rect 35624 15438 35676 15444
rect 35624 15360 35676 15366
rect 35624 15302 35676 15308
rect 35636 14822 35664 15302
rect 35624 14816 35676 14822
rect 35624 14758 35676 14764
rect 35532 12232 35584 12238
rect 35636 12220 35664 14758
rect 36084 14340 36136 14346
rect 36084 14282 36136 14288
rect 35716 13864 35768 13870
rect 35716 13806 35768 13812
rect 35728 12322 35756 13806
rect 36096 13394 36124 14282
rect 36372 14074 36400 19314
rect 36556 19310 36584 20946
rect 37096 20800 37148 20806
rect 37096 20742 37148 20748
rect 37108 20602 37136 20742
rect 37096 20596 37148 20602
rect 37096 20538 37148 20544
rect 37280 20596 37332 20602
rect 37280 20538 37332 20544
rect 37188 20324 37240 20330
rect 37188 20266 37240 20272
rect 37096 20256 37148 20262
rect 37096 20198 37148 20204
rect 36544 19304 36596 19310
rect 36544 19246 36596 19252
rect 37108 18766 37136 20198
rect 37200 19854 37228 20266
rect 37188 19848 37240 19854
rect 37188 19790 37240 19796
rect 37096 18760 37148 18766
rect 37096 18702 37148 18708
rect 37096 18624 37148 18630
rect 37096 18566 37148 18572
rect 36912 17604 36964 17610
rect 36912 17546 36964 17552
rect 36924 16998 36952 17546
rect 36912 16992 36964 16998
rect 36912 16934 36964 16940
rect 36924 16658 36952 16934
rect 36728 16652 36780 16658
rect 36728 16594 36780 16600
rect 36912 16652 36964 16658
rect 36912 16594 36964 16600
rect 36544 16584 36596 16590
rect 36544 16526 36596 16532
rect 36452 15904 36504 15910
rect 36452 15846 36504 15852
rect 36464 15638 36492 15846
rect 36452 15632 36504 15638
rect 36452 15574 36504 15580
rect 36556 15502 36584 16526
rect 36740 16250 36768 16594
rect 36728 16244 36780 16250
rect 36728 16186 36780 16192
rect 36544 15496 36596 15502
rect 36544 15438 36596 15444
rect 36556 15094 36584 15438
rect 36740 15366 36768 16186
rect 37108 15910 37136 18566
rect 37200 17882 37228 19790
rect 37188 17876 37240 17882
rect 37188 17818 37240 17824
rect 37200 16658 37228 17818
rect 37188 16652 37240 16658
rect 37188 16594 37240 16600
rect 37096 15904 37148 15910
rect 37096 15846 37148 15852
rect 36728 15360 36780 15366
rect 37292 15337 37320 20538
rect 37372 19916 37424 19922
rect 37372 19858 37424 19864
rect 37384 18834 37412 19858
rect 37372 18828 37424 18834
rect 37372 18770 37424 18776
rect 37556 16040 37608 16046
rect 37556 15982 37608 15988
rect 37568 15570 37596 15982
rect 37556 15564 37608 15570
rect 37556 15506 37608 15512
rect 36728 15302 36780 15308
rect 37278 15328 37334 15337
rect 37278 15263 37334 15272
rect 36544 15088 36596 15094
rect 36544 15030 36596 15036
rect 37372 14408 37424 14414
rect 37372 14350 37424 14356
rect 37556 14408 37608 14414
rect 37556 14350 37608 14356
rect 37384 14074 37412 14350
rect 36360 14068 36412 14074
rect 36360 14010 36412 14016
rect 37372 14068 37424 14074
rect 37372 14010 37424 14016
rect 37568 14006 37596 14350
rect 37556 14000 37608 14006
rect 37002 13968 37058 13977
rect 36728 13932 36780 13938
rect 37556 13942 37608 13948
rect 37002 13903 37058 13912
rect 36728 13874 36780 13880
rect 35992 13388 36044 13394
rect 35992 13330 36044 13336
rect 36084 13388 36136 13394
rect 36084 13330 36136 13336
rect 35808 13252 35860 13258
rect 35808 13194 35860 13200
rect 35820 12442 35848 13194
rect 36004 12782 36032 13330
rect 36096 12918 36124 13330
rect 36452 13320 36504 13326
rect 36452 13262 36504 13268
rect 36084 12912 36136 12918
rect 36084 12854 36136 12860
rect 35992 12776 36044 12782
rect 35992 12718 36044 12724
rect 36464 12714 36492 13262
rect 36636 13184 36688 13190
rect 36636 13126 36688 13132
rect 36452 12708 36504 12714
rect 36452 12650 36504 12656
rect 35900 12640 35952 12646
rect 35900 12582 35952 12588
rect 36176 12640 36228 12646
rect 36176 12582 36228 12588
rect 35808 12436 35860 12442
rect 35808 12378 35860 12384
rect 35728 12294 35848 12322
rect 35636 12192 35756 12220
rect 35532 12174 35584 12180
rect 35624 11892 35676 11898
rect 35624 11834 35676 11840
rect 35532 11348 35584 11354
rect 35532 11290 35584 11296
rect 35440 10668 35492 10674
rect 35440 10610 35492 10616
rect 35544 10470 35572 11290
rect 35532 10464 35584 10470
rect 35532 10406 35584 10412
rect 35440 9988 35492 9994
rect 35440 9930 35492 9936
rect 35452 8566 35480 9930
rect 35440 8560 35492 8566
rect 35440 8502 35492 8508
rect 35348 7880 35400 7886
rect 35348 7822 35400 7828
rect 35532 7540 35584 7546
rect 35532 7482 35584 7488
rect 34796 7404 34848 7410
rect 34796 7346 34848 7352
rect 34808 6730 34836 7346
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34796 6724 34848 6730
rect 34796 6666 34848 6672
rect 35256 6656 35308 6662
rect 35256 6598 35308 6604
rect 35348 6656 35400 6662
rect 35348 6598 35400 6604
rect 35268 6458 35296 6598
rect 35256 6452 35308 6458
rect 35256 6394 35308 6400
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35164 5636 35216 5642
rect 35164 5578 35216 5584
rect 35176 5273 35204 5578
rect 35360 5370 35388 6598
rect 35544 6390 35572 7482
rect 35532 6384 35584 6390
rect 35532 6326 35584 6332
rect 35636 5914 35664 11834
rect 35728 10826 35756 12192
rect 35820 11218 35848 12294
rect 35912 11218 35940 12582
rect 35992 11552 36044 11558
rect 35992 11494 36044 11500
rect 35808 11212 35860 11218
rect 35808 11154 35860 11160
rect 35900 11212 35952 11218
rect 35900 11154 35952 11160
rect 35820 11098 35848 11154
rect 35820 11070 35940 11098
rect 36004 11082 36032 11494
rect 35912 11014 35940 11070
rect 35992 11076 36044 11082
rect 35992 11018 36044 11024
rect 35900 11008 35952 11014
rect 35900 10950 35952 10956
rect 35728 10798 35940 10826
rect 36188 10810 36216 12582
rect 36648 12306 36676 13126
rect 36636 12300 36688 12306
rect 36636 12242 36688 12248
rect 36636 11552 36688 11558
rect 36636 11494 36688 11500
rect 35716 10464 35768 10470
rect 35912 10452 35940 10798
rect 36176 10804 36228 10810
rect 36176 10746 36228 10752
rect 36544 10532 36596 10538
rect 36544 10474 36596 10480
rect 35716 10406 35768 10412
rect 35820 10424 35940 10452
rect 35728 10062 35756 10406
rect 35716 10056 35768 10062
rect 35716 9998 35768 10004
rect 35820 9110 35848 10424
rect 36084 10260 36136 10266
rect 36084 10202 36136 10208
rect 35900 10056 35952 10062
rect 35900 9998 35952 10004
rect 35912 9761 35940 9998
rect 35898 9752 35954 9761
rect 35898 9687 35954 9696
rect 35992 9580 36044 9586
rect 35992 9522 36044 9528
rect 35900 9376 35952 9382
rect 35900 9318 35952 9324
rect 35808 9104 35860 9110
rect 35808 9046 35860 9052
rect 35912 8974 35940 9318
rect 36004 9217 36032 9522
rect 35990 9208 36046 9217
rect 35990 9143 36046 9152
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 35900 8968 35952 8974
rect 36096 8945 36124 10202
rect 36556 9722 36584 10474
rect 36452 9716 36504 9722
rect 36452 9658 36504 9664
rect 36544 9716 36596 9722
rect 36544 9658 36596 9664
rect 36176 9580 36228 9586
rect 36176 9522 36228 9528
rect 35900 8910 35952 8916
rect 36082 8936 36138 8945
rect 35820 8634 35848 8910
rect 36082 8871 36138 8880
rect 35808 8628 35860 8634
rect 35808 8570 35860 8576
rect 35714 8528 35770 8537
rect 35714 8463 35770 8472
rect 35728 8430 35756 8463
rect 35716 8424 35768 8430
rect 35716 8366 35768 8372
rect 35808 8424 35860 8430
rect 35808 8366 35860 8372
rect 35820 8090 35848 8366
rect 35808 8084 35860 8090
rect 35808 8026 35860 8032
rect 36188 7993 36216 9522
rect 36268 9376 36320 9382
rect 36268 9318 36320 9324
rect 36280 9042 36308 9318
rect 36268 9036 36320 9042
rect 36268 8978 36320 8984
rect 36360 8968 36412 8974
rect 36360 8910 36412 8916
rect 36372 8566 36400 8910
rect 36360 8560 36412 8566
rect 36360 8502 36412 8508
rect 36268 8288 36320 8294
rect 36268 8230 36320 8236
rect 36174 7984 36230 7993
rect 36174 7919 36230 7928
rect 36084 7880 36136 7886
rect 36084 7822 36136 7828
rect 36096 7478 36124 7822
rect 36084 7472 36136 7478
rect 36084 7414 36136 7420
rect 36084 6316 36136 6322
rect 36084 6258 36136 6264
rect 35532 5908 35584 5914
rect 35532 5850 35584 5856
rect 35624 5908 35676 5914
rect 35624 5850 35676 5856
rect 35820 5902 36032 5930
rect 35544 5794 35572 5850
rect 35820 5794 35848 5902
rect 35544 5766 35848 5794
rect 36004 5778 36032 5902
rect 35440 5704 35492 5710
rect 35492 5664 35572 5692
rect 35440 5646 35492 5652
rect 35348 5364 35400 5370
rect 35348 5306 35400 5312
rect 35162 5264 35218 5273
rect 35162 5199 35218 5208
rect 34980 5160 35032 5166
rect 35348 5160 35400 5166
rect 35032 5108 35348 5114
rect 34980 5102 35400 5108
rect 34992 5086 35388 5102
rect 35440 5092 35492 5098
rect 35440 5034 35492 5040
rect 34796 5024 34848 5030
rect 34796 4966 34848 4972
rect 34612 4150 34664 4156
rect 34702 4176 34758 4185
rect 34702 4111 34758 4120
rect 34612 4072 34664 4078
rect 34612 4014 34664 4020
rect 34704 4072 34756 4078
rect 34704 4014 34756 4020
rect 34624 3602 34652 4014
rect 34612 3596 34664 3602
rect 34612 3538 34664 3544
rect 34520 3052 34572 3058
rect 34520 2994 34572 3000
rect 33600 2984 33652 2990
rect 34716 2938 34744 4014
rect 34808 3534 34836 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35348 4548 35400 4554
rect 35348 4490 35400 4496
rect 35360 4146 35388 4490
rect 35348 4140 35400 4146
rect 35348 4082 35400 4088
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 33600 2926 33652 2932
rect 34532 2910 34744 2938
rect 33508 2372 33560 2378
rect 33508 2314 33560 2320
rect 33520 1018 33548 2314
rect 33784 1148 33836 1154
rect 33784 1090 33836 1096
rect 33508 1012 33560 1018
rect 33508 954 33560 960
rect 33428 870 33548 898
rect 33520 800 33548 870
rect 33796 800 33824 1090
rect 34060 944 34112 950
rect 34532 898 34560 2910
rect 34808 2774 34836 3334
rect 35452 3058 35480 5034
rect 35440 3052 35492 3058
rect 35440 2994 35492 3000
rect 35544 2774 35572 5664
rect 35820 5574 35848 5766
rect 35900 5772 35952 5778
rect 35900 5714 35952 5720
rect 35992 5772 36044 5778
rect 35992 5714 36044 5720
rect 35808 5568 35860 5574
rect 35808 5510 35860 5516
rect 35716 5160 35768 5166
rect 35716 5102 35768 5108
rect 35624 4072 35676 4078
rect 35624 4014 35676 4020
rect 35636 3398 35664 4014
rect 35624 3392 35676 3398
rect 35624 3334 35676 3340
rect 35624 2984 35676 2990
rect 35624 2926 35676 2932
rect 34716 2746 34836 2774
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34716 2122 34744 2746
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35452 2746 35572 2774
rect 34888 2440 34940 2446
rect 34888 2382 34940 2388
rect 34060 886 34112 892
rect 34072 800 34100 886
rect 34348 870 34560 898
rect 34624 2094 34744 2122
rect 34348 800 34376 870
rect 34624 800 34652 2094
rect 34900 2038 34928 2382
rect 35164 2372 35216 2378
rect 35164 2314 35216 2320
rect 34888 2032 34940 2038
rect 34888 1974 34940 1980
rect 35176 1086 35204 2314
rect 35452 2310 35480 2746
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 35164 1080 35216 1086
rect 35164 1022 35216 1028
rect 35636 1018 35664 2926
rect 35624 1012 35676 1018
rect 35624 954 35676 960
rect 34900 870 35020 898
rect 34900 800 34928 870
rect 4526 0 4582 800
rect 4802 0 4858 800
rect 5078 0 5134 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 34992 202 35020 870
rect 35176 870 35296 898
rect 35176 800 35204 870
rect 34980 196 35032 202
rect 34980 138 35032 144
rect 35162 0 35218 800
rect 35268 406 35296 870
rect 35452 870 35572 898
rect 35452 800 35480 870
rect 35256 400 35308 406
rect 35256 342 35308 348
rect 35438 0 35494 800
rect 35544 134 35572 870
rect 35728 800 35756 5102
rect 35912 4146 35940 5714
rect 35992 5568 36044 5574
rect 35992 5510 36044 5516
rect 36004 5302 36032 5510
rect 35992 5296 36044 5302
rect 35992 5238 36044 5244
rect 35992 5024 36044 5030
rect 35992 4966 36044 4972
rect 36004 4554 36032 4966
rect 35992 4548 36044 4554
rect 35992 4490 36044 4496
rect 35900 4140 35952 4146
rect 35900 4082 35952 4088
rect 35898 4040 35954 4049
rect 35898 3975 35954 3984
rect 35912 3534 35940 3975
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36096 2774 36124 6258
rect 36280 5778 36308 8230
rect 36360 7744 36412 7750
rect 36360 7686 36412 7692
rect 36268 5772 36320 5778
rect 36268 5714 36320 5720
rect 36268 5636 36320 5642
rect 36268 5578 36320 5584
rect 36174 5264 36230 5273
rect 36280 5234 36308 5578
rect 36372 5574 36400 7686
rect 36464 6458 36492 9658
rect 36544 9444 36596 9450
rect 36544 9386 36596 9392
rect 36556 8634 36584 9386
rect 36544 8628 36596 8634
rect 36544 8570 36596 8576
rect 36648 8514 36676 11494
rect 36740 9042 36768 13874
rect 37016 12434 37044 13903
rect 37280 13728 37332 13734
rect 37280 13670 37332 13676
rect 37292 12850 37320 13670
rect 37280 12844 37332 12850
rect 37280 12786 37332 12792
rect 37292 12434 37320 12786
rect 37752 12434 37780 22066
rect 37832 19168 37884 19174
rect 37832 19110 37884 19116
rect 37844 18737 37872 19110
rect 37830 18728 37886 18737
rect 37830 18663 37886 18672
rect 37924 15156 37976 15162
rect 37924 15098 37976 15104
rect 37936 14550 37964 15098
rect 38016 14612 38068 14618
rect 38016 14554 38068 14560
rect 37924 14544 37976 14550
rect 37924 14486 37976 14492
rect 37936 14074 37964 14486
rect 37924 14068 37976 14074
rect 37924 14010 37976 14016
rect 38028 13938 38056 14554
rect 38016 13932 38068 13938
rect 38016 13874 38068 13880
rect 38016 13524 38068 13530
rect 38016 13466 38068 13472
rect 38028 12918 38056 13466
rect 38016 12912 38068 12918
rect 38016 12854 38068 12860
rect 38028 12442 38056 12854
rect 38016 12436 38068 12442
rect 37016 12406 37136 12434
rect 37292 12406 37412 12434
rect 37752 12406 37872 12434
rect 36820 11212 36872 11218
rect 36820 11154 36872 11160
rect 36728 9036 36780 9042
rect 36728 8978 36780 8984
rect 36556 8486 36676 8514
rect 36728 8492 36780 8498
rect 36556 8294 36584 8486
rect 36728 8434 36780 8440
rect 36636 8424 36688 8430
rect 36636 8366 36688 8372
rect 36544 8288 36596 8294
rect 36544 8230 36596 8236
rect 36542 7984 36598 7993
rect 36542 7919 36598 7928
rect 36556 7750 36584 7919
rect 36544 7744 36596 7750
rect 36544 7686 36596 7692
rect 36556 7478 36584 7686
rect 36544 7472 36596 7478
rect 36544 7414 36596 7420
rect 36452 6452 36504 6458
rect 36452 6394 36504 6400
rect 36360 5568 36412 5574
rect 36360 5510 36412 5516
rect 36174 5199 36230 5208
rect 36268 5228 36320 5234
rect 36188 3058 36216 5199
rect 36268 5170 36320 5176
rect 36372 4826 36400 5510
rect 36360 4820 36412 4826
rect 36360 4762 36412 4768
rect 36358 4720 36414 4729
rect 36358 4655 36414 4664
rect 36372 4554 36400 4655
rect 36360 4548 36412 4554
rect 36360 4490 36412 4496
rect 36268 4480 36320 4486
rect 36268 4422 36320 4428
rect 36176 3052 36228 3058
rect 36176 2994 36228 3000
rect 36004 2746 36124 2774
rect 36004 800 36032 2746
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 36096 1222 36124 2314
rect 36084 1216 36136 1222
rect 36084 1158 36136 1164
rect 36280 800 36308 4422
rect 36450 4176 36506 4185
rect 36450 4111 36506 4120
rect 36464 1034 36492 4111
rect 36648 3738 36676 8366
rect 36740 7546 36768 8434
rect 36832 7698 36860 11154
rect 36912 8288 36964 8294
rect 36912 8230 36964 8236
rect 36924 7886 36952 8230
rect 36912 7880 36964 7886
rect 36912 7822 36964 7828
rect 37004 7812 37056 7818
rect 37004 7754 37056 7760
rect 36832 7670 36952 7698
rect 36728 7540 36780 7546
rect 36728 7482 36780 7488
rect 36728 7404 36780 7410
rect 36728 7346 36780 7352
rect 36740 6254 36768 7346
rect 36820 7336 36872 7342
rect 36820 7278 36872 7284
rect 36832 6866 36860 7278
rect 36820 6860 36872 6866
rect 36820 6802 36872 6808
rect 36728 6248 36780 6254
rect 36728 6190 36780 6196
rect 36832 5778 36860 6802
rect 36924 6390 36952 7670
rect 37016 7478 37044 7754
rect 37004 7472 37056 7478
rect 37004 7414 37056 7420
rect 36912 6384 36964 6390
rect 36912 6326 36964 6332
rect 37108 5778 37136 12406
rect 37384 11082 37412 12406
rect 37372 11076 37424 11082
rect 37372 11018 37424 11024
rect 37280 9920 37332 9926
rect 37280 9862 37332 9868
rect 37188 8968 37240 8974
rect 37188 8910 37240 8916
rect 37200 6225 37228 8910
rect 37186 6216 37242 6225
rect 37186 6151 37242 6160
rect 36820 5772 36872 5778
rect 36820 5714 36872 5720
rect 37096 5772 37148 5778
rect 37096 5714 37148 5720
rect 36728 5636 36780 5642
rect 36728 5578 36780 5584
rect 36740 4486 36768 5578
rect 36820 5568 36872 5574
rect 36820 5510 36872 5516
rect 36728 4480 36780 4486
rect 36728 4422 36780 4428
rect 36636 3732 36688 3738
rect 36636 3674 36688 3680
rect 36544 2984 36596 2990
rect 36544 2926 36596 2932
rect 36556 1154 36584 2926
rect 36544 1148 36596 1154
rect 36544 1090 36596 1096
rect 36464 1006 36584 1034
rect 36556 800 36584 1006
rect 36832 800 36860 5510
rect 37004 5160 37056 5166
rect 37004 5102 37056 5108
rect 36912 4752 36964 4758
rect 36912 4694 36964 4700
rect 36924 3534 36952 4694
rect 37016 4622 37044 5102
rect 37004 4616 37056 4622
rect 37004 4558 37056 4564
rect 37016 3602 37044 4558
rect 37094 4040 37150 4049
rect 37094 3975 37150 3984
rect 37004 3596 37056 3602
rect 37004 3538 37056 3544
rect 36912 3528 36964 3534
rect 36912 3470 36964 3476
rect 36924 2990 36952 3470
rect 36912 2984 36964 2990
rect 36912 2926 36964 2932
rect 37108 800 37136 3975
rect 37292 3058 37320 9862
rect 37384 8566 37412 11018
rect 37556 10736 37608 10742
rect 37556 10678 37608 10684
rect 37568 9489 37596 10678
rect 37738 10160 37794 10169
rect 37738 10095 37794 10104
rect 37752 9586 37780 10095
rect 37648 9580 37700 9586
rect 37648 9522 37700 9528
rect 37740 9580 37792 9586
rect 37740 9522 37792 9528
rect 37554 9480 37610 9489
rect 37554 9415 37610 9424
rect 37556 9376 37608 9382
rect 37462 9344 37518 9353
rect 37556 9318 37608 9324
rect 37462 9279 37518 9288
rect 37476 8974 37504 9279
rect 37464 8968 37516 8974
rect 37464 8910 37516 8916
rect 37372 8560 37424 8566
rect 37372 8502 37424 8508
rect 37384 8294 37412 8502
rect 37568 8498 37596 9318
rect 37556 8492 37608 8498
rect 37556 8434 37608 8440
rect 37372 8288 37424 8294
rect 37372 8230 37424 8236
rect 37556 7812 37608 7818
rect 37556 7754 37608 7760
rect 37372 4820 37424 4826
rect 37372 4762 37424 4768
rect 37384 4282 37412 4762
rect 37372 4276 37424 4282
rect 37372 4218 37424 4224
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 37464 2848 37516 2854
rect 37464 2790 37516 2796
rect 37476 2360 37504 2790
rect 37384 2332 37504 2360
rect 37384 800 37412 2332
rect 37568 1358 37596 7754
rect 37660 5914 37688 9522
rect 37740 9444 37792 9450
rect 37740 9386 37792 9392
rect 37752 9178 37780 9386
rect 37740 9172 37792 9178
rect 37740 9114 37792 9120
rect 37844 9042 37872 12406
rect 38016 12378 38068 12384
rect 37924 12096 37976 12102
rect 37924 12038 37976 12044
rect 37936 9586 37964 12038
rect 38120 11218 38148 22066
rect 39040 21554 39068 22066
rect 39028 21548 39080 21554
rect 39028 21490 39080 21496
rect 38568 21344 38620 21350
rect 38568 21286 38620 21292
rect 38476 21140 38528 21146
rect 38476 21082 38528 21088
rect 38488 20942 38516 21082
rect 38580 20942 38608 21286
rect 38476 20936 38528 20942
rect 38476 20878 38528 20884
rect 38568 20936 38620 20942
rect 38568 20878 38620 20884
rect 38384 20392 38436 20398
rect 38488 20380 38516 20878
rect 38752 20800 38804 20806
rect 38752 20742 38804 20748
rect 38764 20466 38792 20742
rect 38752 20460 38804 20466
rect 38752 20402 38804 20408
rect 38436 20352 38516 20380
rect 38384 20334 38436 20340
rect 38200 19712 38252 19718
rect 38200 19654 38252 19660
rect 38212 15910 38240 19654
rect 38844 18760 38896 18766
rect 38844 18702 38896 18708
rect 38856 18306 38884 18702
rect 38660 18284 38712 18290
rect 38660 18226 38712 18232
rect 38764 18278 38884 18306
rect 38672 17610 38700 18226
rect 38764 17814 38792 18278
rect 38844 18216 38896 18222
rect 38844 18158 38896 18164
rect 38856 17882 38884 18158
rect 38844 17876 38896 17882
rect 38844 17818 38896 17824
rect 38936 17876 38988 17882
rect 38936 17818 38988 17824
rect 38752 17808 38804 17814
rect 38752 17750 38804 17756
rect 38660 17604 38712 17610
rect 38660 17546 38712 17552
rect 38948 17542 38976 17818
rect 38936 17536 38988 17542
rect 38936 17478 38988 17484
rect 38292 17332 38344 17338
rect 38292 17274 38344 17280
rect 38304 16590 38332 17274
rect 38844 17128 38896 17134
rect 38844 17070 38896 17076
rect 39040 17082 39068 21490
rect 39212 21480 39264 21486
rect 39212 21422 39264 21428
rect 39224 19378 39252 21422
rect 39212 19372 39264 19378
rect 39212 19314 39264 19320
rect 39120 18624 39172 18630
rect 39120 18566 39172 18572
rect 39132 18290 39160 18566
rect 39120 18284 39172 18290
rect 39120 18226 39172 18232
rect 39224 17746 39252 19314
rect 39212 17740 39264 17746
rect 39212 17682 39264 17688
rect 39210 17640 39266 17649
rect 39210 17575 39212 17584
rect 39264 17575 39266 17584
rect 39212 17546 39264 17552
rect 39224 17270 39252 17546
rect 39212 17264 39264 17270
rect 39212 17206 39264 17212
rect 38292 16584 38344 16590
rect 38292 16526 38344 16532
rect 38856 16454 38884 17070
rect 39040 17054 39252 17082
rect 38844 16448 38896 16454
rect 38844 16390 38896 16396
rect 38200 15904 38252 15910
rect 38200 15846 38252 15852
rect 38212 11665 38240 15846
rect 38752 14952 38804 14958
rect 38752 14894 38804 14900
rect 38660 13932 38712 13938
rect 38660 13874 38712 13880
rect 38292 13320 38344 13326
rect 38292 13262 38344 13268
rect 38198 11656 38254 11665
rect 38198 11591 38254 11600
rect 38108 11212 38160 11218
rect 38108 11154 38160 11160
rect 38304 10554 38332 13262
rect 38672 12850 38700 13874
rect 38764 13870 38792 14894
rect 38752 13864 38804 13870
rect 38752 13806 38804 13812
rect 38764 13326 38792 13806
rect 38856 13462 38884 16390
rect 38936 14816 38988 14822
rect 38936 14758 38988 14764
rect 39120 14816 39172 14822
rect 39120 14758 39172 14764
rect 38948 13938 38976 14758
rect 39028 14340 39080 14346
rect 39028 14282 39080 14288
rect 39040 14074 39068 14282
rect 39132 14278 39160 14758
rect 39120 14272 39172 14278
rect 39120 14214 39172 14220
rect 39028 14068 39080 14074
rect 39028 14010 39080 14016
rect 38936 13932 38988 13938
rect 38936 13874 38988 13880
rect 38844 13456 38896 13462
rect 38844 13398 38896 13404
rect 38752 13320 38804 13326
rect 38752 13262 38804 13268
rect 39120 13320 39172 13326
rect 39120 13262 39172 13268
rect 38660 12844 38712 12850
rect 38660 12786 38712 12792
rect 38384 12436 38436 12442
rect 39132 12434 39160 13262
rect 38384 12378 38436 12384
rect 39040 12406 39160 12434
rect 38396 12102 38424 12378
rect 38384 12096 38436 12102
rect 38384 12038 38436 12044
rect 38752 11756 38804 11762
rect 38752 11698 38804 11704
rect 38476 11144 38528 11150
rect 38528 11104 38608 11132
rect 38476 11086 38528 11092
rect 38384 11076 38436 11082
rect 38384 11018 38436 11024
rect 38396 10792 38424 11018
rect 38396 10764 38516 10792
rect 38384 10668 38436 10674
rect 38384 10610 38436 10616
rect 38396 10577 38424 10610
rect 38120 10526 38332 10554
rect 38382 10568 38438 10577
rect 38016 10464 38068 10470
rect 38016 10406 38068 10412
rect 38028 10169 38056 10406
rect 38014 10160 38070 10169
rect 38014 10095 38070 10104
rect 38120 9654 38148 10526
rect 38382 10503 38438 10512
rect 38488 10418 38516 10764
rect 38212 10390 38516 10418
rect 38212 10198 38240 10390
rect 38200 10192 38252 10198
rect 38580 10169 38608 11104
rect 38658 10976 38714 10985
rect 38658 10911 38714 10920
rect 38200 10134 38252 10140
rect 38290 10160 38346 10169
rect 38108 9648 38160 9654
rect 38014 9616 38070 9625
rect 37924 9580 37976 9586
rect 38108 9590 38160 9596
rect 38014 9551 38070 9560
rect 37924 9522 37976 9528
rect 37922 9480 37978 9489
rect 37922 9415 37978 9424
rect 37832 9036 37884 9042
rect 37832 8978 37884 8984
rect 37936 8480 37964 9415
rect 38028 9178 38056 9551
rect 38016 9172 38068 9178
rect 38016 9114 38068 9120
rect 38108 9036 38160 9042
rect 38108 8978 38160 8984
rect 38120 8498 38148 8978
rect 38212 8906 38240 10134
rect 38290 10095 38346 10104
rect 38566 10160 38622 10169
rect 38566 10095 38622 10104
rect 38304 10062 38332 10095
rect 38292 10056 38344 10062
rect 38292 9998 38344 10004
rect 38672 9994 38700 10911
rect 38660 9988 38712 9994
rect 38660 9930 38712 9936
rect 38292 9920 38344 9926
rect 38384 9920 38436 9926
rect 38292 9862 38344 9868
rect 38382 9888 38384 9897
rect 38436 9888 38438 9897
rect 38304 9738 38332 9862
rect 38382 9823 38438 9832
rect 38566 9888 38622 9897
rect 38566 9823 38622 9832
rect 38304 9710 38516 9738
rect 38384 9648 38436 9654
rect 38384 9590 38436 9596
rect 38290 9208 38346 9217
rect 38290 9143 38346 9152
rect 38304 9110 38332 9143
rect 38292 9104 38344 9110
rect 38292 9046 38344 9052
rect 38200 8900 38252 8906
rect 38200 8842 38252 8848
rect 37844 8452 37964 8480
rect 38108 8492 38160 8498
rect 37740 8356 37792 8362
rect 37740 8298 37792 8304
rect 37648 5908 37700 5914
rect 37648 5850 37700 5856
rect 37752 5098 37780 8298
rect 37740 5092 37792 5098
rect 37740 5034 37792 5040
rect 37752 4622 37780 5034
rect 37844 4758 37872 8452
rect 38108 8434 38160 8440
rect 38292 8492 38344 8498
rect 38292 8434 38344 8440
rect 38108 7880 38160 7886
rect 38108 7822 38160 7828
rect 38200 7880 38252 7886
rect 38200 7822 38252 7828
rect 38120 7546 38148 7822
rect 38108 7540 38160 7546
rect 38108 7482 38160 7488
rect 38212 6186 38240 7822
rect 38304 7818 38332 8434
rect 38292 7812 38344 7818
rect 38292 7754 38344 7760
rect 38396 7750 38424 9590
rect 38384 7744 38436 7750
rect 38384 7686 38436 7692
rect 38396 7410 38424 7686
rect 38384 7404 38436 7410
rect 38384 7346 38436 7352
rect 38488 6474 38516 9710
rect 38580 8974 38608 9823
rect 38660 9104 38712 9110
rect 38660 9046 38712 9052
rect 38568 8968 38620 8974
rect 38568 8910 38620 8916
rect 38580 8809 38608 8910
rect 38566 8800 38622 8809
rect 38566 8735 38622 8744
rect 38672 8362 38700 9046
rect 38660 8356 38712 8362
rect 38660 8298 38712 8304
rect 38488 6446 38608 6474
rect 38476 6316 38528 6322
rect 38476 6258 38528 6264
rect 38200 6180 38252 6186
rect 38200 6122 38252 6128
rect 38016 5228 38068 5234
rect 38016 5170 38068 5176
rect 38028 4758 38056 5170
rect 37832 4752 37884 4758
rect 37832 4694 37884 4700
rect 38016 4752 38068 4758
rect 38016 4694 38068 4700
rect 37740 4616 37792 4622
rect 37740 4558 37792 4564
rect 37832 4616 37884 4622
rect 37832 4558 37884 4564
rect 37844 4282 37872 4558
rect 38016 4480 38068 4486
rect 38016 4422 38068 4428
rect 37832 4276 37884 4282
rect 37832 4218 37884 4224
rect 37740 4208 37792 4214
rect 37740 4150 37792 4156
rect 37752 3369 37780 4150
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 37844 3777 37872 4082
rect 37830 3768 37886 3777
rect 37830 3703 37886 3712
rect 38028 3602 38056 4422
rect 38212 4298 38240 6122
rect 38382 5808 38438 5817
rect 38382 5743 38384 5752
rect 38436 5743 38438 5752
rect 38384 5714 38436 5720
rect 38108 4276 38160 4282
rect 38212 4270 38332 4298
rect 38108 4218 38160 4224
rect 38016 3596 38068 3602
rect 38016 3538 38068 3544
rect 37924 3392 37976 3398
rect 37738 3360 37794 3369
rect 37924 3334 37976 3340
rect 37738 3295 37794 3304
rect 37648 3188 37700 3194
rect 37648 3130 37700 3136
rect 37556 1352 37608 1358
rect 37556 1294 37608 1300
rect 37660 800 37688 3130
rect 37936 3126 37964 3334
rect 37924 3120 37976 3126
rect 37924 3062 37976 3068
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 37752 950 37780 2314
rect 38120 2122 38148 4218
rect 38200 4208 38252 4214
rect 38198 4176 38200 4185
rect 38252 4176 38254 4185
rect 38198 4111 38254 4120
rect 38198 4040 38254 4049
rect 38198 3975 38200 3984
rect 38252 3975 38254 3984
rect 38200 3946 38252 3952
rect 38304 3777 38332 4270
rect 38290 3768 38346 3777
rect 38200 3732 38252 3738
rect 38290 3703 38346 3712
rect 38200 3674 38252 3680
rect 37936 2094 38148 2122
rect 37740 944 37792 950
rect 37740 886 37792 892
rect 37936 800 37964 2094
rect 38212 800 38240 3674
rect 38304 3670 38332 3703
rect 38292 3664 38344 3670
rect 38292 3606 38344 3612
rect 38488 800 38516 6258
rect 38580 3126 38608 6446
rect 38660 5024 38712 5030
rect 38660 4966 38712 4972
rect 38568 3120 38620 3126
rect 38568 3062 38620 3068
rect 38672 3058 38700 4966
rect 38660 3052 38712 3058
rect 38660 2994 38712 3000
rect 38660 2916 38712 2922
rect 38660 2858 38712 2864
rect 38672 2514 38700 2858
rect 38660 2508 38712 2514
rect 38660 2450 38712 2456
rect 38660 2372 38712 2378
rect 38660 2314 38712 2320
rect 35532 128 35584 134
rect 35532 70 35584 76
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38672 202 38700 2314
rect 38764 1358 38792 11698
rect 38844 11212 38896 11218
rect 38844 11154 38896 11160
rect 38856 6458 38884 11154
rect 39040 11082 39068 12406
rect 39224 11286 39252 17054
rect 39304 15156 39356 15162
rect 39304 15098 39356 15104
rect 39212 11280 39264 11286
rect 39212 11222 39264 11228
rect 39028 11076 39080 11082
rect 39028 11018 39080 11024
rect 38936 8832 38988 8838
rect 38936 8774 38988 8780
rect 38948 8634 38976 8774
rect 38936 8628 38988 8634
rect 38936 8570 38988 8576
rect 38936 8492 38988 8498
rect 38936 8434 38988 8440
rect 38844 6452 38896 6458
rect 38844 6394 38896 6400
rect 38948 5658 38976 8434
rect 39040 7954 39068 11018
rect 39316 10130 39344 15098
rect 39408 11082 39436 42298
rect 39948 36712 40000 36718
rect 39948 36654 40000 36660
rect 39960 35562 39988 36654
rect 39948 35556 40000 35562
rect 39948 35498 40000 35504
rect 40040 35080 40092 35086
rect 40040 35022 40092 35028
rect 40052 34474 40080 35022
rect 40040 34468 40092 34474
rect 40040 34410 40092 34416
rect 40040 34196 40092 34202
rect 40040 34138 40092 34144
rect 40052 33522 40080 34138
rect 40040 33516 40092 33522
rect 40040 33458 40092 33464
rect 39764 24336 39816 24342
rect 39764 24278 39816 24284
rect 39488 22976 39540 22982
rect 39488 22918 39540 22924
rect 39396 11076 39448 11082
rect 39396 11018 39448 11024
rect 39304 10124 39356 10130
rect 39304 10066 39356 10072
rect 39120 9988 39172 9994
rect 39120 9930 39172 9936
rect 39132 8673 39160 9930
rect 39396 9444 39448 9450
rect 39396 9386 39448 9392
rect 39118 8664 39174 8673
rect 39118 8599 39174 8608
rect 39302 8664 39358 8673
rect 39302 8599 39358 8608
rect 39212 8492 39264 8498
rect 39212 8434 39264 8440
rect 39224 8090 39252 8434
rect 39316 8430 39344 8599
rect 39304 8424 39356 8430
rect 39304 8366 39356 8372
rect 39212 8084 39264 8090
rect 39212 8026 39264 8032
rect 39028 7948 39080 7954
rect 39028 7890 39080 7896
rect 39028 6996 39080 7002
rect 39028 6938 39080 6944
rect 38856 5642 38976 5658
rect 38844 5636 38976 5642
rect 38896 5630 38976 5636
rect 38844 5578 38896 5584
rect 38856 5030 38884 5578
rect 38936 5568 38988 5574
rect 38936 5510 38988 5516
rect 38844 5024 38896 5030
rect 38844 4966 38896 4972
rect 38856 4826 38884 4966
rect 38844 4820 38896 4826
rect 38844 4762 38896 4768
rect 38948 4622 38976 5510
rect 38936 4616 38988 4622
rect 38936 4558 38988 4564
rect 39040 4554 39068 6938
rect 39120 5228 39172 5234
rect 39120 5170 39172 5176
rect 39212 5228 39264 5234
rect 39212 5170 39264 5176
rect 39132 4826 39160 5170
rect 39120 4820 39172 4826
rect 39120 4762 39172 4768
rect 39120 4684 39172 4690
rect 39120 4626 39172 4632
rect 39028 4548 39080 4554
rect 39028 4490 39080 4496
rect 38844 4480 38896 4486
rect 38844 4422 38896 4428
rect 38856 3534 38884 4422
rect 39028 3664 39080 3670
rect 39028 3606 39080 3612
rect 38844 3528 38896 3534
rect 38844 3470 38896 3476
rect 38844 3392 38896 3398
rect 38844 3334 38896 3340
rect 38856 2922 38884 3334
rect 38936 2984 38988 2990
rect 38936 2926 38988 2932
rect 38844 2916 38896 2922
rect 38844 2858 38896 2864
rect 38844 2372 38896 2378
rect 38844 2314 38896 2320
rect 38752 1352 38804 1358
rect 38752 1294 38804 1300
rect 38752 1216 38804 1222
rect 38752 1158 38804 1164
rect 38764 800 38792 1158
rect 38660 196 38712 202
rect 38660 138 38712 144
rect 38750 0 38806 800
rect 38856 134 38884 2314
rect 38948 406 38976 2926
rect 39040 800 39068 3606
rect 39132 3466 39160 4626
rect 39120 3460 39172 3466
rect 39120 3402 39172 3408
rect 39132 2446 39160 3402
rect 39120 2440 39172 2446
rect 39120 2382 39172 2388
rect 39224 1222 39252 5170
rect 39408 4146 39436 9386
rect 39396 4140 39448 4146
rect 39396 4082 39448 4088
rect 39396 3460 39448 3466
rect 39396 3402 39448 3408
rect 39408 3194 39436 3402
rect 39396 3188 39448 3194
rect 39396 3130 39448 3136
rect 39304 3052 39356 3058
rect 39304 2994 39356 3000
rect 39212 1216 39264 1222
rect 39212 1158 39264 1164
rect 39316 800 39344 2994
rect 39500 2582 39528 22918
rect 39580 22160 39632 22166
rect 39580 22102 39632 22108
rect 39592 5370 39620 22102
rect 39672 20324 39724 20330
rect 39672 20266 39724 20272
rect 39684 12986 39712 20266
rect 39672 12980 39724 12986
rect 39672 12922 39724 12928
rect 39672 12844 39724 12850
rect 39672 12786 39724 12792
rect 39684 8566 39712 12786
rect 39672 8560 39724 8566
rect 39672 8502 39724 8508
rect 39580 5364 39632 5370
rect 39580 5306 39632 5312
rect 39776 3194 39804 24278
rect 40052 21570 40080 33458
rect 39960 21542 40080 21570
rect 39960 20482 39988 21542
rect 40040 21412 40092 21418
rect 40040 21354 40092 21360
rect 40052 20602 40080 21354
rect 40040 20596 40092 20602
rect 40040 20538 40092 20544
rect 39960 20454 40080 20482
rect 40052 19310 40080 20454
rect 40040 19304 40092 19310
rect 40040 19246 40092 19252
rect 40052 19145 40080 19246
rect 40038 19136 40094 19145
rect 40038 19071 40094 19080
rect 39856 17740 39908 17746
rect 39856 17682 39908 17688
rect 39868 4078 39896 17682
rect 39948 17128 40000 17134
rect 39948 17070 40000 17076
rect 39960 11014 39988 17070
rect 40040 16652 40092 16658
rect 40040 16594 40092 16600
rect 40052 16250 40080 16594
rect 40144 16250 40172 53654
rect 40328 35086 40356 60998
rect 40960 60512 41012 60518
rect 40960 60454 41012 60460
rect 40972 60110 41000 60454
rect 41432 60330 41460 61066
rect 41524 60790 41552 63294
rect 41604 63300 41656 63306
rect 41604 63242 41656 63248
rect 41616 61198 41644 63242
rect 42062 63200 42118 64000
rect 42798 63200 42854 64000
rect 43534 63200 43590 64000
rect 44270 63322 44326 64000
rect 45006 63322 45062 64000
rect 44270 63294 44588 63322
rect 44270 63200 44326 63294
rect 41788 61668 41840 61674
rect 41788 61610 41840 61616
rect 41604 61192 41656 61198
rect 41604 61134 41656 61140
rect 41696 61056 41748 61062
rect 41696 60998 41748 61004
rect 41512 60784 41564 60790
rect 41512 60726 41564 60732
rect 41156 60302 41460 60330
rect 41156 60246 41184 60302
rect 41144 60240 41196 60246
rect 41144 60182 41196 60188
rect 41236 60240 41288 60246
rect 41236 60182 41288 60188
rect 41604 60240 41656 60246
rect 41604 60182 41656 60188
rect 40960 60104 41012 60110
rect 40960 60046 41012 60052
rect 40868 60036 40920 60042
rect 40868 59978 40920 59984
rect 40880 59498 40908 59978
rect 40868 59492 40920 59498
rect 40868 59434 40920 59440
rect 40776 50448 40828 50454
rect 40776 50390 40828 50396
rect 40408 47796 40460 47802
rect 40408 47738 40460 47744
rect 40316 35080 40368 35086
rect 40316 35022 40368 35028
rect 40316 29640 40368 29646
rect 40316 29582 40368 29588
rect 40224 19848 40276 19854
rect 40224 19790 40276 19796
rect 40236 17746 40264 19790
rect 40224 17740 40276 17746
rect 40224 17682 40276 17688
rect 40224 16992 40276 16998
rect 40224 16934 40276 16940
rect 40236 16697 40264 16934
rect 40222 16688 40278 16697
rect 40222 16623 40278 16632
rect 40040 16244 40092 16250
rect 40040 16186 40092 16192
rect 40132 16244 40184 16250
rect 40132 16186 40184 16192
rect 40040 15020 40092 15026
rect 40040 14962 40092 14968
rect 40052 14278 40080 14962
rect 40040 14272 40092 14278
rect 40040 14214 40092 14220
rect 40038 12336 40094 12345
rect 40038 12271 40094 12280
rect 40052 12238 40080 12271
rect 40040 12232 40092 12238
rect 40040 12174 40092 12180
rect 40224 11076 40276 11082
rect 40224 11018 40276 11024
rect 39948 11008 40000 11014
rect 39948 10950 40000 10956
rect 39960 10198 39988 10950
rect 40040 10600 40092 10606
rect 40040 10542 40092 10548
rect 39948 10192 40000 10198
rect 39948 10134 40000 10140
rect 40052 9042 40080 10542
rect 40040 9036 40092 9042
rect 40040 8978 40092 8984
rect 40132 8968 40184 8974
rect 40132 8910 40184 8916
rect 39948 8492 40000 8498
rect 40000 8452 40080 8480
rect 39948 8434 40000 8440
rect 40052 8294 40080 8452
rect 40144 8362 40172 8910
rect 40132 8356 40184 8362
rect 40132 8298 40184 8304
rect 40040 8288 40092 8294
rect 40040 8230 40092 8236
rect 39946 8120 40002 8129
rect 39946 8055 40002 8064
rect 39960 8022 39988 8055
rect 39948 8016 40000 8022
rect 39948 7958 40000 7964
rect 40040 8016 40092 8022
rect 40040 7958 40092 7964
rect 40052 6866 40080 7958
rect 40130 6896 40186 6905
rect 40040 6860 40092 6866
rect 40130 6831 40186 6840
rect 40040 6802 40092 6808
rect 40052 5778 40080 6802
rect 40040 5772 40092 5778
rect 40040 5714 40092 5720
rect 40040 4616 40092 4622
rect 40040 4558 40092 4564
rect 39856 4072 39908 4078
rect 39856 4014 39908 4020
rect 39764 3188 39816 3194
rect 39764 3130 39816 3136
rect 40052 2854 40080 4558
rect 40144 4146 40172 6831
rect 40236 4826 40264 11018
rect 40224 4820 40276 4826
rect 40224 4762 40276 4768
rect 40224 4616 40276 4622
rect 40224 4558 40276 4564
rect 40132 4140 40184 4146
rect 40132 4082 40184 4088
rect 40236 3670 40264 4558
rect 40224 3664 40276 3670
rect 40224 3606 40276 3612
rect 40328 3194 40356 29582
rect 40420 12238 40448 47738
rect 40592 35692 40644 35698
rect 40592 35634 40644 35640
rect 40604 35494 40632 35634
rect 40592 35488 40644 35494
rect 40592 35430 40644 35436
rect 40500 35080 40552 35086
rect 40500 35022 40552 35028
rect 40512 34202 40540 35022
rect 40500 34196 40552 34202
rect 40500 34138 40552 34144
rect 40684 30932 40736 30938
rect 40684 30874 40736 30880
rect 40696 30258 40724 30874
rect 40592 30252 40644 30258
rect 40592 30194 40644 30200
rect 40684 30252 40736 30258
rect 40684 30194 40736 30200
rect 40500 19780 40552 19786
rect 40500 19722 40552 19728
rect 40512 19514 40540 19722
rect 40500 19508 40552 19514
rect 40500 19450 40552 19456
rect 40500 19304 40552 19310
rect 40500 19246 40552 19252
rect 40512 18834 40540 19246
rect 40500 18828 40552 18834
rect 40500 18770 40552 18776
rect 40500 18624 40552 18630
rect 40500 18566 40552 18572
rect 40512 17678 40540 18566
rect 40500 17672 40552 17678
rect 40500 17614 40552 17620
rect 40500 16448 40552 16454
rect 40500 16390 40552 16396
rect 40512 16182 40540 16390
rect 40500 16176 40552 16182
rect 40500 16118 40552 16124
rect 40500 13932 40552 13938
rect 40500 13874 40552 13880
rect 40408 12232 40460 12238
rect 40408 12174 40460 12180
rect 40512 11082 40540 13874
rect 40500 11076 40552 11082
rect 40500 11018 40552 11024
rect 40604 9466 40632 30194
rect 40684 20596 40736 20602
rect 40684 20538 40736 20544
rect 40696 19786 40724 20538
rect 40684 19780 40736 19786
rect 40684 19722 40736 19728
rect 40684 16720 40736 16726
rect 40684 16662 40736 16668
rect 40696 16590 40724 16662
rect 40684 16584 40736 16590
rect 40684 16526 40736 16532
rect 40788 14929 40816 50390
rect 40880 36650 40908 59434
rect 41144 58880 41196 58886
rect 41144 58822 41196 58828
rect 41156 57050 41184 58822
rect 41144 57044 41196 57050
rect 41144 56986 41196 56992
rect 41248 56352 41276 60182
rect 41616 60110 41644 60182
rect 41604 60104 41656 60110
rect 41604 60046 41656 60052
rect 41616 59090 41644 60046
rect 41604 59084 41656 59090
rect 41604 59026 41656 59032
rect 41512 59016 41564 59022
rect 41512 58958 41564 58964
rect 41420 56772 41472 56778
rect 41420 56714 41472 56720
rect 41156 56324 41276 56352
rect 41052 55276 41104 55282
rect 41052 55218 41104 55224
rect 41064 53650 41092 55218
rect 41052 53644 41104 53650
rect 41052 53586 41104 53592
rect 41156 51814 41184 56324
rect 41432 56302 41460 56714
rect 41524 56370 41552 58958
rect 41616 58410 41644 59026
rect 41604 58404 41656 58410
rect 41604 58346 41656 58352
rect 41512 56364 41564 56370
rect 41512 56306 41564 56312
rect 41420 56296 41472 56302
rect 41420 56238 41472 56244
rect 41236 56228 41288 56234
rect 41236 56170 41288 56176
rect 41248 55282 41276 56170
rect 41328 56160 41380 56166
rect 41328 56102 41380 56108
rect 41236 55276 41288 55282
rect 41236 55218 41288 55224
rect 41248 53582 41276 55218
rect 41340 55214 41368 56102
rect 41524 55418 41552 56306
rect 41616 56234 41644 58346
rect 41604 56228 41656 56234
rect 41604 56170 41656 56176
rect 41512 55412 41564 55418
rect 41512 55354 41564 55360
rect 41340 55186 41552 55214
rect 41236 53576 41288 53582
rect 41236 53518 41288 53524
rect 41144 51808 41196 51814
rect 41144 51750 41196 51756
rect 41420 40724 41472 40730
rect 41420 40666 41472 40672
rect 40868 36644 40920 36650
rect 40868 36586 40920 36592
rect 41328 19508 41380 19514
rect 41328 19450 41380 19456
rect 40960 19168 41012 19174
rect 40960 19110 41012 19116
rect 40972 18766 41000 19110
rect 41236 18828 41288 18834
rect 41236 18770 41288 18776
rect 40960 18760 41012 18766
rect 40960 18702 41012 18708
rect 41144 18624 41196 18630
rect 41144 18566 41196 18572
rect 40960 18216 41012 18222
rect 40960 18158 41012 18164
rect 41156 18170 41184 18566
rect 41248 18358 41276 18770
rect 41236 18352 41288 18358
rect 41236 18294 41288 18300
rect 40972 17202 41000 18158
rect 41156 18142 41276 18170
rect 41248 17814 41276 18142
rect 41236 17808 41288 17814
rect 41236 17750 41288 17756
rect 41144 17264 41196 17270
rect 41144 17206 41196 17212
rect 40960 17196 41012 17202
rect 40960 17138 41012 17144
rect 40868 17128 40920 17134
rect 40868 17070 40920 17076
rect 40880 15978 40908 17070
rect 41156 16794 41184 17206
rect 41144 16788 41196 16794
rect 41144 16730 41196 16736
rect 40960 16584 41012 16590
rect 40960 16526 41012 16532
rect 41052 16584 41104 16590
rect 41052 16526 41104 16532
rect 40972 16250 41000 16526
rect 41064 16250 41092 16526
rect 40960 16244 41012 16250
rect 40960 16186 41012 16192
rect 41052 16244 41104 16250
rect 41052 16186 41104 16192
rect 40868 15972 40920 15978
rect 40868 15914 40920 15920
rect 41248 15858 41276 17750
rect 41340 17134 41368 19450
rect 41328 17128 41380 17134
rect 41328 17070 41380 17076
rect 41328 16720 41380 16726
rect 41328 16662 41380 16668
rect 40972 15830 41276 15858
rect 40868 15088 40920 15094
rect 40868 15030 40920 15036
rect 40774 14920 40830 14929
rect 40774 14855 40830 14864
rect 40880 14822 40908 15030
rect 40868 14816 40920 14822
rect 40868 14758 40920 14764
rect 40684 14408 40736 14414
rect 40684 14350 40736 14356
rect 40696 10810 40724 14350
rect 40774 14240 40830 14249
rect 40774 14175 40830 14184
rect 40684 10804 40736 10810
rect 40684 10746 40736 10752
rect 40696 10606 40724 10746
rect 40684 10600 40736 10606
rect 40684 10542 40736 10548
rect 40604 9438 40724 9466
rect 40592 9376 40644 9382
rect 40592 9318 40644 9324
rect 40406 8936 40462 8945
rect 40406 8871 40462 8880
rect 40420 4010 40448 8871
rect 40604 8634 40632 9318
rect 40592 8628 40644 8634
rect 40592 8570 40644 8576
rect 40500 5228 40552 5234
rect 40500 5170 40552 5176
rect 40408 4004 40460 4010
rect 40408 3946 40460 3952
rect 40408 3664 40460 3670
rect 40406 3632 40408 3641
rect 40460 3632 40462 3641
rect 40406 3567 40462 3576
rect 40316 3188 40368 3194
rect 40316 3130 40368 3136
rect 40132 3052 40184 3058
rect 40132 2994 40184 3000
rect 40040 2848 40092 2854
rect 40040 2790 40092 2796
rect 39488 2576 39540 2582
rect 39488 2518 39540 2524
rect 39856 1284 39908 1290
rect 39856 1226 39908 1232
rect 39580 944 39632 950
rect 39580 886 39632 892
rect 39592 800 39620 886
rect 39868 800 39896 1226
rect 40144 800 40172 2994
rect 40512 2666 40540 5170
rect 40592 5160 40644 5166
rect 40592 5102 40644 5108
rect 40604 3602 40632 5102
rect 40696 4826 40724 9438
rect 40788 7750 40816 14175
rect 40868 12708 40920 12714
rect 40868 12650 40920 12656
rect 40880 12170 40908 12650
rect 40868 12164 40920 12170
rect 40868 12106 40920 12112
rect 40972 11801 41000 15830
rect 41340 15586 41368 16662
rect 41156 15558 41368 15586
rect 41052 15496 41104 15502
rect 41052 15438 41104 15444
rect 41064 12434 41092 15438
rect 41156 12714 41184 15558
rect 41340 15502 41368 15558
rect 41432 15502 41460 40666
rect 41524 19122 41552 55186
rect 41708 35834 41736 60998
rect 41800 59634 41828 61610
rect 42076 61198 42104 63200
rect 42812 61198 42840 63200
rect 43548 63170 43576 63200
rect 43536 63164 43588 63170
rect 43536 63106 43588 63112
rect 44364 63164 44416 63170
rect 44364 63106 44416 63112
rect 44376 61198 44404 63106
rect 44560 61198 44588 63294
rect 45006 63294 45600 63322
rect 45006 63200 45062 63294
rect 45572 61198 45600 63294
rect 45742 63200 45798 64000
rect 46478 63322 46534 64000
rect 46478 63294 46704 63322
rect 46478 63200 46534 63294
rect 45756 61198 45784 63200
rect 42064 61192 42116 61198
rect 42064 61134 42116 61140
rect 42800 61192 42852 61198
rect 42800 61134 42852 61140
rect 44364 61192 44416 61198
rect 44364 61134 44416 61140
rect 44548 61192 44600 61198
rect 44548 61134 44600 61140
rect 45560 61192 45612 61198
rect 45560 61134 45612 61140
rect 45744 61192 45796 61198
rect 45744 61134 45796 61140
rect 42984 61124 43036 61130
rect 42984 61066 43036 61072
rect 44824 61124 44876 61130
rect 44824 61066 44876 61072
rect 42248 60580 42300 60586
rect 42248 60522 42300 60528
rect 42260 60178 42288 60522
rect 42248 60172 42300 60178
rect 42248 60114 42300 60120
rect 42708 60172 42760 60178
rect 42708 60114 42760 60120
rect 42432 60104 42484 60110
rect 42432 60046 42484 60052
rect 42064 60036 42116 60042
rect 42064 59978 42116 59984
rect 41788 59628 41840 59634
rect 41788 59570 41840 59576
rect 42076 59401 42104 59978
rect 42444 59974 42472 60046
rect 42432 59968 42484 59974
rect 42432 59910 42484 59916
rect 42444 59702 42472 59910
rect 42432 59696 42484 59702
rect 42432 59638 42484 59644
rect 42720 59650 42748 60114
rect 42720 59622 42840 59650
rect 42812 59566 42840 59622
rect 42708 59560 42760 59566
rect 42708 59502 42760 59508
rect 42800 59560 42852 59566
rect 42800 59502 42852 59508
rect 42062 59392 42118 59401
rect 42062 59327 42118 59336
rect 42616 58336 42668 58342
rect 42616 58278 42668 58284
rect 42064 55276 42116 55282
rect 42064 55218 42116 55224
rect 41696 35828 41748 35834
rect 41696 35770 41748 35776
rect 41972 22432 42024 22438
rect 41972 22374 42024 22380
rect 41880 21004 41932 21010
rect 41880 20946 41932 20952
rect 41892 20806 41920 20946
rect 41984 20942 42012 22374
rect 41972 20936 42024 20942
rect 41972 20878 42024 20884
rect 41604 20800 41656 20806
rect 41604 20742 41656 20748
rect 41880 20800 41932 20806
rect 41880 20742 41932 20748
rect 41616 20466 41644 20742
rect 41604 20460 41656 20466
rect 41604 20402 41656 20408
rect 41696 20392 41748 20398
rect 41696 20334 41748 20340
rect 41708 19378 41736 20334
rect 41788 20256 41840 20262
rect 41788 20198 41840 20204
rect 41880 20256 41932 20262
rect 41880 20198 41932 20204
rect 41800 19786 41828 20198
rect 41788 19780 41840 19786
rect 41788 19722 41840 19728
rect 41892 19378 41920 20198
rect 41696 19372 41748 19378
rect 41696 19314 41748 19320
rect 41880 19372 41932 19378
rect 41880 19314 41932 19320
rect 41984 19258 42012 20878
rect 41892 19230 42012 19258
rect 41524 19094 41644 19122
rect 41512 18352 41564 18358
rect 41512 18294 41564 18300
rect 41524 16697 41552 18294
rect 41510 16688 41566 16697
rect 41510 16623 41566 16632
rect 41616 16046 41644 19094
rect 41696 16448 41748 16454
rect 41748 16396 41828 16402
rect 41696 16390 41828 16396
rect 41708 16374 41828 16390
rect 41800 16182 41828 16374
rect 41788 16176 41840 16182
rect 41788 16118 41840 16124
rect 41696 16108 41748 16114
rect 41696 16050 41748 16056
rect 41604 16040 41656 16046
rect 41604 15982 41656 15988
rect 41512 15972 41564 15978
rect 41512 15914 41564 15920
rect 41236 15496 41288 15502
rect 41236 15438 41288 15444
rect 41328 15496 41380 15502
rect 41328 15438 41380 15444
rect 41420 15496 41472 15502
rect 41420 15438 41472 15444
rect 41144 12708 41196 12714
rect 41144 12650 41196 12656
rect 41064 12406 41184 12434
rect 41156 12238 41184 12406
rect 41144 12232 41196 12238
rect 41142 12200 41144 12209
rect 41196 12200 41198 12209
rect 41142 12135 41198 12144
rect 41144 12096 41196 12102
rect 41144 12038 41196 12044
rect 41050 11928 41106 11937
rect 41050 11863 41106 11872
rect 41064 11830 41092 11863
rect 41052 11824 41104 11830
rect 40958 11792 41014 11801
rect 41052 11766 41104 11772
rect 41156 11762 41184 12038
rect 40958 11727 41014 11736
rect 41144 11756 41196 11762
rect 41144 11698 41196 11704
rect 40960 11076 41012 11082
rect 40960 11018 41012 11024
rect 41052 11076 41104 11082
rect 41052 11018 41104 11024
rect 40776 7744 40828 7750
rect 40776 7686 40828 7692
rect 40684 4820 40736 4826
rect 40684 4762 40736 4768
rect 40868 4548 40920 4554
rect 40868 4490 40920 4496
rect 40880 3738 40908 4490
rect 40868 3732 40920 3738
rect 40868 3674 40920 3680
rect 40592 3596 40644 3602
rect 40592 3538 40644 3544
rect 40776 3528 40828 3534
rect 40776 3470 40828 3476
rect 40788 2990 40816 3470
rect 40776 2984 40828 2990
rect 40776 2926 40828 2932
rect 40420 2638 40540 2666
rect 40420 800 40448 2638
rect 40972 2106 41000 11018
rect 41064 4690 41092 11018
rect 41248 5098 41276 15438
rect 41524 15162 41552 15914
rect 41708 15706 41736 16050
rect 41696 15700 41748 15706
rect 41696 15642 41748 15648
rect 41604 15496 41656 15502
rect 41604 15438 41656 15444
rect 41512 15156 41564 15162
rect 41512 15098 41564 15104
rect 41616 15026 41644 15438
rect 41512 15020 41564 15026
rect 41512 14962 41564 14968
rect 41604 15020 41656 15026
rect 41604 14962 41656 14968
rect 41524 14929 41552 14962
rect 41510 14920 41566 14929
rect 41510 14855 41566 14864
rect 41512 14272 41564 14278
rect 41512 14214 41564 14220
rect 41328 14000 41380 14006
rect 41524 13954 41552 14214
rect 41328 13942 41380 13948
rect 41340 13734 41368 13942
rect 41432 13926 41552 13954
rect 41432 13870 41460 13926
rect 41420 13864 41472 13870
rect 41420 13806 41472 13812
rect 41328 13728 41380 13734
rect 41328 13670 41380 13676
rect 41616 12764 41644 14962
rect 41786 13968 41842 13977
rect 41696 13932 41748 13938
rect 41786 13903 41788 13912
rect 41696 13874 41748 13880
rect 41840 13903 41842 13912
rect 41788 13874 41840 13880
rect 41708 13394 41736 13874
rect 41696 13388 41748 13394
rect 41696 13330 41748 13336
rect 41616 12736 41736 12764
rect 41420 12708 41472 12714
rect 41420 12650 41472 12656
rect 41432 12238 41460 12650
rect 41708 12374 41736 12736
rect 41604 12368 41656 12374
rect 41510 12336 41566 12345
rect 41604 12310 41656 12316
rect 41696 12368 41748 12374
rect 41696 12310 41748 12316
rect 41510 12271 41566 12280
rect 41524 12238 41552 12271
rect 41328 12232 41380 12238
rect 41328 12174 41380 12180
rect 41420 12232 41472 12238
rect 41420 12174 41472 12180
rect 41512 12232 41564 12238
rect 41512 12174 41564 12180
rect 41340 11801 41368 12174
rect 41326 11792 41382 11801
rect 41326 11727 41382 11736
rect 41510 11792 41566 11801
rect 41510 11727 41566 11736
rect 41328 11688 41380 11694
rect 41328 11630 41380 11636
rect 41340 11354 41368 11630
rect 41328 11348 41380 11354
rect 41328 11290 41380 11296
rect 41328 10668 41380 10674
rect 41328 10610 41380 10616
rect 41340 10266 41368 10610
rect 41328 10260 41380 10266
rect 41328 10202 41380 10208
rect 41420 9580 41472 9586
rect 41420 9522 41472 9528
rect 41432 9178 41460 9522
rect 41420 9172 41472 9178
rect 41420 9114 41472 9120
rect 41524 7206 41552 11727
rect 41616 11098 41644 12310
rect 41788 12096 41840 12102
rect 41788 12038 41840 12044
rect 41800 11218 41828 12038
rect 41788 11212 41840 11218
rect 41788 11154 41840 11160
rect 41616 11070 41736 11098
rect 41604 10464 41656 10470
rect 41604 10406 41656 10412
rect 41512 7200 41564 7206
rect 41512 7142 41564 7148
rect 41420 5636 41472 5642
rect 41420 5578 41472 5584
rect 41236 5092 41288 5098
rect 41236 5034 41288 5040
rect 41144 5024 41196 5030
rect 41144 4966 41196 4972
rect 41052 4684 41104 4690
rect 41052 4626 41104 4632
rect 41052 3732 41104 3738
rect 41052 3674 41104 3680
rect 41064 3126 41092 3674
rect 41156 3534 41184 4966
rect 41326 3904 41382 3913
rect 41326 3839 41382 3848
rect 41340 3602 41368 3839
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 41144 3528 41196 3534
rect 41144 3470 41196 3476
rect 41236 3528 41288 3534
rect 41236 3470 41288 3476
rect 41052 3120 41104 3126
rect 41052 3062 41104 3068
rect 41248 2922 41276 3470
rect 41236 2916 41288 2922
rect 41236 2858 41288 2864
rect 41432 2802 41460 5578
rect 41616 4146 41644 10406
rect 41708 5409 41736 11070
rect 41788 10464 41840 10470
rect 41788 10406 41840 10412
rect 41800 10130 41828 10406
rect 41788 10124 41840 10130
rect 41788 10066 41840 10072
rect 41892 9994 41920 19230
rect 42076 16590 42104 55218
rect 42248 21480 42300 21486
rect 42248 21422 42300 21428
rect 42340 21480 42392 21486
rect 42340 21422 42392 21428
rect 42260 21010 42288 21422
rect 42352 21146 42380 21422
rect 42340 21140 42392 21146
rect 42340 21082 42392 21088
rect 42248 21004 42300 21010
rect 42248 20946 42300 20952
rect 42352 19394 42380 21082
rect 42260 19366 42380 19394
rect 41972 16584 42024 16590
rect 41972 16526 42024 16532
rect 42064 16584 42116 16590
rect 42064 16526 42116 16532
rect 41984 15162 42012 16526
rect 42064 16108 42116 16114
rect 42064 16050 42116 16056
rect 42076 15706 42104 16050
rect 42064 15700 42116 15706
rect 42064 15642 42116 15648
rect 42064 15564 42116 15570
rect 42064 15506 42116 15512
rect 41972 15156 42024 15162
rect 41972 15098 42024 15104
rect 41972 14408 42024 14414
rect 41972 14350 42024 14356
rect 41984 13258 42012 14350
rect 41972 13252 42024 13258
rect 41972 13194 42024 13200
rect 41984 12714 42012 13194
rect 41972 12708 42024 12714
rect 41972 12650 42024 12656
rect 41972 11824 42024 11830
rect 41972 11766 42024 11772
rect 41984 11150 42012 11766
rect 41972 11144 42024 11150
rect 41972 11086 42024 11092
rect 41880 9988 41932 9994
rect 41880 9930 41932 9936
rect 41694 5400 41750 5409
rect 41694 5335 41750 5344
rect 41880 5228 41932 5234
rect 41880 5170 41932 5176
rect 41604 4140 41656 4146
rect 41604 4082 41656 4088
rect 41786 4040 41842 4049
rect 41696 4004 41748 4010
rect 41786 3975 41842 3984
rect 41696 3946 41748 3952
rect 41708 3738 41736 3946
rect 41696 3732 41748 3738
rect 41696 3674 41748 3680
rect 41800 3194 41828 3975
rect 41788 3188 41840 3194
rect 41788 3130 41840 3136
rect 41512 3052 41564 3058
rect 41512 2994 41564 3000
rect 41248 2774 41460 2802
rect 41052 2372 41104 2378
rect 41052 2314 41104 2320
rect 40960 2100 41012 2106
rect 40960 2042 41012 2048
rect 40960 1216 41012 1222
rect 40960 1158 41012 1164
rect 40684 1012 40736 1018
rect 40684 954 40736 960
rect 40696 800 40724 954
rect 40972 800 41000 1158
rect 41064 950 41092 2314
rect 41052 944 41104 950
rect 41052 886 41104 892
rect 41248 800 41276 2774
rect 41524 800 41552 2994
rect 41892 2774 41920 5170
rect 42076 4282 42104 15506
rect 42260 15162 42288 19366
rect 42340 19304 42392 19310
rect 42340 19246 42392 19252
rect 42248 15156 42300 15162
rect 42248 15098 42300 15104
rect 42260 14414 42288 15098
rect 42352 14414 42380 19246
rect 42524 18760 42576 18766
rect 42524 18702 42576 18708
rect 42430 18456 42486 18465
rect 42430 18391 42486 18400
rect 42444 18290 42472 18391
rect 42432 18284 42484 18290
rect 42432 18226 42484 18232
rect 42430 18184 42486 18193
rect 42430 18119 42486 18128
rect 42444 18086 42472 18119
rect 42536 18086 42564 18702
rect 42432 18080 42484 18086
rect 42432 18022 42484 18028
rect 42524 18080 42576 18086
rect 42524 18022 42576 18028
rect 42432 16108 42484 16114
rect 42432 16050 42484 16056
rect 42248 14408 42300 14414
rect 42248 14350 42300 14356
rect 42340 14408 42392 14414
rect 42340 14350 42392 14356
rect 42156 12776 42208 12782
rect 42156 12718 42208 12724
rect 42064 4276 42116 4282
rect 42064 4218 42116 4224
rect 42064 4140 42116 4146
rect 42064 4082 42116 4088
rect 41800 2746 41920 2774
rect 41800 800 41828 2746
rect 42076 800 42104 4082
rect 42168 3670 42196 12718
rect 42246 11928 42302 11937
rect 42246 11863 42248 11872
rect 42300 11863 42302 11872
rect 42248 11834 42300 11840
rect 42248 11756 42300 11762
rect 42248 11698 42300 11704
rect 42340 11756 42392 11762
rect 42340 11698 42392 11704
rect 42260 11218 42288 11698
rect 42248 11212 42300 11218
rect 42248 11154 42300 11160
rect 42352 11082 42380 11698
rect 42340 11076 42392 11082
rect 42340 11018 42392 11024
rect 42340 10124 42392 10130
rect 42340 10066 42392 10072
rect 42352 8673 42380 10066
rect 42338 8664 42394 8673
rect 42338 8599 42394 8608
rect 42156 3664 42208 3670
rect 42156 3606 42208 3612
rect 42444 2106 42472 16050
rect 42524 13728 42576 13734
rect 42524 13670 42576 13676
rect 42536 13326 42564 13670
rect 42524 13320 42576 13326
rect 42524 13262 42576 13268
rect 42524 13184 42576 13190
rect 42524 13126 42576 13132
rect 42536 11082 42564 13126
rect 42628 11354 42656 58278
rect 42720 56681 42748 59502
rect 42706 56672 42762 56681
rect 42706 56607 42762 56616
rect 42996 36922 43024 61066
rect 44180 60512 44232 60518
rect 44180 60454 44232 60460
rect 43260 57044 43312 57050
rect 43260 56986 43312 56992
rect 43076 49088 43128 49094
rect 43076 49030 43128 49036
rect 42984 36916 43036 36922
rect 42984 36858 43036 36864
rect 42892 24404 42944 24410
rect 42892 24346 42944 24352
rect 42708 20800 42760 20806
rect 42708 20742 42760 20748
rect 42720 19990 42748 20742
rect 42800 20460 42852 20466
rect 42800 20402 42852 20408
rect 42812 20058 42840 20402
rect 42800 20052 42852 20058
rect 42800 19994 42852 20000
rect 42708 19984 42760 19990
rect 42904 19938 42932 24346
rect 42984 21344 43036 21350
rect 42984 21286 43036 21292
rect 42708 19926 42760 19932
rect 42812 19910 42932 19938
rect 42706 19136 42762 19145
rect 42706 19071 42762 19080
rect 42720 18766 42748 19071
rect 42812 18816 42840 19910
rect 42892 19848 42944 19854
rect 42892 19790 42944 19796
rect 42904 19378 42932 19790
rect 42996 19786 43024 21286
rect 42984 19780 43036 19786
rect 42984 19722 43036 19728
rect 42892 19372 42944 19378
rect 42892 19314 42944 19320
rect 42812 18788 43024 18816
rect 42708 18760 42760 18766
rect 42708 18702 42760 18708
rect 42890 18728 42946 18737
rect 42800 18692 42852 18698
rect 42890 18663 42892 18672
rect 42800 18634 42852 18640
rect 42944 18663 42946 18672
rect 42892 18634 42944 18640
rect 42708 18624 42760 18630
rect 42708 18566 42760 18572
rect 42720 16454 42748 18566
rect 42812 16658 42840 18634
rect 42890 18592 42946 18601
rect 42890 18527 42946 18536
rect 42904 18358 42932 18527
rect 42892 18352 42944 18358
rect 42892 18294 42944 18300
rect 42996 18290 43024 18788
rect 42984 18284 43036 18290
rect 42984 18226 43036 18232
rect 42892 18216 42944 18222
rect 42892 18158 42944 18164
rect 42800 16652 42852 16658
rect 42800 16594 42852 16600
rect 42708 16448 42760 16454
rect 42708 16390 42760 16396
rect 42708 16176 42760 16182
rect 42760 16136 42840 16164
rect 42708 16118 42760 16124
rect 42812 15858 42840 16136
rect 42904 16046 42932 18158
rect 42996 16114 43024 18226
rect 43088 16182 43116 49030
rect 43168 18624 43220 18630
rect 43168 18566 43220 18572
rect 43180 18426 43208 18566
rect 43168 18420 43220 18426
rect 43168 18362 43220 18368
rect 43076 16176 43128 16182
rect 43076 16118 43128 16124
rect 42984 16108 43036 16114
rect 42984 16050 43036 16056
rect 42892 16040 42944 16046
rect 42892 15982 42944 15988
rect 42812 15830 42932 15858
rect 42708 15088 42760 15094
rect 42708 15030 42760 15036
rect 42720 14822 42748 15030
rect 42800 15020 42852 15026
rect 42800 14962 42852 14968
rect 42708 14816 42760 14822
rect 42708 14758 42760 14764
rect 42708 14408 42760 14414
rect 42708 14350 42760 14356
rect 42720 13326 42748 14350
rect 42708 13320 42760 13326
rect 42708 13262 42760 13268
rect 42720 12850 42748 13262
rect 42812 12986 42840 14962
rect 42800 12980 42852 12986
rect 42800 12922 42852 12928
rect 42708 12844 42760 12850
rect 42708 12786 42760 12792
rect 42616 11348 42668 11354
rect 42616 11290 42668 11296
rect 42524 11076 42576 11082
rect 42524 11018 42576 11024
rect 42536 5137 42564 11018
rect 42720 10130 42748 12786
rect 42812 12646 42840 12922
rect 42904 12730 42932 15830
rect 42996 15502 43024 16050
rect 42984 15496 43036 15502
rect 42984 15438 43036 15444
rect 42984 14816 43036 14822
rect 42984 14758 43036 14764
rect 42996 14482 43024 14758
rect 43272 14634 43300 56986
rect 44192 55350 44220 60454
rect 44180 55344 44232 55350
rect 44180 55286 44232 55292
rect 44836 53514 44864 61066
rect 45376 61056 45428 61062
rect 45376 60998 45428 61004
rect 44824 53508 44876 53514
rect 44824 53450 44876 53456
rect 45388 53106 45416 60998
rect 46676 60790 46704 63294
rect 47214 63200 47270 64000
rect 47950 63322 48006 64000
rect 47950 63294 48360 63322
rect 47950 63200 48006 63294
rect 46848 61600 46900 61606
rect 46848 61542 46900 61548
rect 46860 61402 46888 61542
rect 46848 61396 46900 61402
rect 46848 61338 46900 61344
rect 47228 61198 47256 63200
rect 48332 61198 48360 63294
rect 48686 63200 48742 64000
rect 49422 63322 49478 64000
rect 49422 63294 49832 63322
rect 49422 63200 49478 63294
rect 48700 61198 48728 63200
rect 49424 61736 49476 61742
rect 49424 61678 49476 61684
rect 49436 61402 49464 61678
rect 49424 61396 49476 61402
rect 49424 61338 49476 61344
rect 49804 61198 49832 63294
rect 50158 63200 50214 64000
rect 50894 63322 50950 64000
rect 50894 63294 51304 63322
rect 50894 63200 50950 63294
rect 47216 61192 47268 61198
rect 47216 61134 47268 61140
rect 48320 61192 48372 61198
rect 48320 61134 48372 61140
rect 48688 61192 48740 61198
rect 48688 61134 48740 61140
rect 49792 61192 49844 61198
rect 49792 61134 49844 61140
rect 49700 61124 49752 61130
rect 49700 61066 49752 61072
rect 46848 61056 46900 61062
rect 46848 60998 46900 61004
rect 46664 60784 46716 60790
rect 46664 60726 46716 60732
rect 46860 56370 46888 60998
rect 49712 58546 49740 61066
rect 50068 61056 50120 61062
rect 50068 60998 50120 61004
rect 49700 58540 49752 58546
rect 49700 58482 49752 58488
rect 46848 56364 46900 56370
rect 46848 56306 46900 56312
rect 45376 53100 45428 53106
rect 45376 53042 45428 53048
rect 50080 51074 50108 60998
rect 50172 60790 50200 63200
rect 51276 61198 51304 63294
rect 51630 63200 51686 64000
rect 52366 63322 52422 64000
rect 53102 63322 53158 64000
rect 53838 63322 53894 64000
rect 54574 63322 54630 64000
rect 55310 63322 55366 64000
rect 52366 63294 52684 63322
rect 52366 63200 52422 63294
rect 51644 61198 51672 63200
rect 51264 61192 51316 61198
rect 51264 61134 51316 61140
rect 51632 61192 51684 61198
rect 51632 61134 51684 61140
rect 50620 61056 50672 61062
rect 50620 60998 50672 61004
rect 50294 60956 50602 60965
rect 50294 60954 50300 60956
rect 50356 60954 50380 60956
rect 50436 60954 50460 60956
rect 50516 60954 50540 60956
rect 50596 60954 50602 60956
rect 50356 60902 50358 60954
rect 50538 60902 50540 60954
rect 50294 60900 50300 60902
rect 50356 60900 50380 60902
rect 50436 60900 50460 60902
rect 50516 60900 50540 60902
rect 50596 60900 50602 60902
rect 50294 60891 50602 60900
rect 50160 60784 50212 60790
rect 50160 60726 50212 60732
rect 50436 60512 50488 60518
rect 50436 60454 50488 60460
rect 50448 60178 50476 60454
rect 50436 60172 50488 60178
rect 50436 60114 50488 60120
rect 50294 59868 50602 59877
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59803 50602 59812
rect 50632 59090 50660 60998
rect 52656 60790 52684 63294
rect 53102 63294 53236 63322
rect 53102 63200 53158 63294
rect 53208 61198 53236 63294
rect 53838 63294 54156 63322
rect 53838 63200 53894 63294
rect 54128 61198 54156 63294
rect 54574 63294 54708 63322
rect 54574 63200 54630 63294
rect 53196 61192 53248 61198
rect 53196 61134 53248 61140
rect 54116 61192 54168 61198
rect 54116 61134 54168 61140
rect 53472 61124 53524 61130
rect 53472 61066 53524 61072
rect 52644 60784 52696 60790
rect 52644 60726 52696 60732
rect 53104 60512 53156 60518
rect 53104 60454 53156 60460
rect 53116 59634 53144 60454
rect 53104 59628 53156 59634
rect 53104 59570 53156 59576
rect 50620 59084 50672 59090
rect 50620 59026 50672 59032
rect 50294 58780 50602 58789
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58715 50602 58724
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50080 51046 50200 51074
rect 44088 47728 44140 47734
rect 44088 47670 44140 47676
rect 43352 29640 43404 29646
rect 43352 29582 43404 29588
rect 43364 20874 43392 29582
rect 43720 21548 43772 21554
rect 43720 21490 43772 21496
rect 43352 20868 43404 20874
rect 43352 20810 43404 20816
rect 43628 20800 43680 20806
rect 43628 20742 43680 20748
rect 43352 20392 43404 20398
rect 43352 20334 43404 20340
rect 43364 19514 43392 20334
rect 43444 20052 43496 20058
rect 43444 19994 43496 20000
rect 43352 19508 43404 19514
rect 43352 19450 43404 19456
rect 43456 18630 43484 19994
rect 43640 19446 43668 20742
rect 43732 20466 43760 21490
rect 43812 20868 43864 20874
rect 43812 20810 43864 20816
rect 43720 20460 43772 20466
rect 43720 20402 43772 20408
rect 43628 19440 43680 19446
rect 43628 19382 43680 19388
rect 43640 18698 43668 19382
rect 43720 18964 43772 18970
rect 43720 18906 43772 18912
rect 43732 18766 43760 18906
rect 43720 18760 43772 18766
rect 43720 18702 43772 18708
rect 43628 18692 43680 18698
rect 43628 18634 43680 18640
rect 43444 18624 43496 18630
rect 43444 18566 43496 18572
rect 43442 18456 43498 18465
rect 43442 18391 43498 18400
rect 43456 18086 43484 18391
rect 43640 18358 43668 18634
rect 43628 18352 43680 18358
rect 43628 18294 43680 18300
rect 43444 18080 43496 18086
rect 43444 18022 43496 18028
rect 43444 16516 43496 16522
rect 43444 16458 43496 16464
rect 43180 14606 43300 14634
rect 42984 14476 43036 14482
rect 42984 14418 43036 14424
rect 42996 14226 43024 14418
rect 42996 14198 43116 14226
rect 42984 14068 43036 14074
rect 42984 14010 43036 14016
rect 42996 12850 43024 14010
rect 43088 13938 43116 14198
rect 43076 13932 43128 13938
rect 43076 13874 43128 13880
rect 43180 13410 43208 14606
rect 43260 14476 43312 14482
rect 43260 14418 43312 14424
rect 43272 13530 43300 14418
rect 43352 13864 43404 13870
rect 43352 13806 43404 13812
rect 43260 13524 43312 13530
rect 43260 13466 43312 13472
rect 43180 13382 43300 13410
rect 42984 12844 43036 12850
rect 42984 12786 43036 12792
rect 42904 12702 43208 12730
rect 42800 12640 42852 12646
rect 42800 12582 42852 12588
rect 43076 12640 43128 12646
rect 43076 12582 43128 12588
rect 42984 11144 43036 11150
rect 42984 11086 43036 11092
rect 42708 10124 42760 10130
rect 42708 10066 42760 10072
rect 42708 9104 42760 9110
rect 42708 9046 42760 9052
rect 42720 8566 42748 9046
rect 42708 8560 42760 8566
rect 42708 8502 42760 8508
rect 42720 7886 42748 8502
rect 42708 7880 42760 7886
rect 42708 7822 42760 7828
rect 42706 5536 42762 5545
rect 42706 5471 42762 5480
rect 42522 5128 42578 5137
rect 42522 5063 42578 5072
rect 42720 4622 42748 5471
rect 42892 5228 42944 5234
rect 42892 5170 42944 5176
rect 42708 4616 42760 4622
rect 42708 4558 42760 4564
rect 42616 4072 42668 4078
rect 42616 4014 42668 4020
rect 42628 3233 42656 4014
rect 42708 3732 42760 3738
rect 42708 3674 42760 3680
rect 42614 3224 42670 3233
rect 42614 3159 42670 3168
rect 42616 3120 42668 3126
rect 42614 3088 42616 3097
rect 42668 3088 42670 3097
rect 42614 3023 42670 3032
rect 42432 2100 42484 2106
rect 42432 2042 42484 2048
rect 42720 2038 42748 3674
rect 42708 2032 42760 2038
rect 42708 1974 42760 1980
rect 42616 1080 42668 1086
rect 42616 1022 42668 1028
rect 42340 944 42392 950
rect 42340 886 42392 892
rect 42352 800 42380 886
rect 42628 800 42656 1022
rect 42904 800 42932 5170
rect 42996 4554 43024 11086
rect 43088 6662 43116 12582
rect 43076 6656 43128 6662
rect 43076 6598 43128 6604
rect 43180 5370 43208 12702
rect 43272 11218 43300 13382
rect 43364 12986 43392 13806
rect 43352 12980 43404 12986
rect 43352 12922 43404 12928
rect 43456 12434 43484 16458
rect 43534 13968 43590 13977
rect 43534 13903 43590 13912
rect 43548 13870 43576 13903
rect 43536 13864 43588 13870
rect 43536 13806 43588 13812
rect 43456 12406 43576 12434
rect 43444 12300 43496 12306
rect 43444 12242 43496 12248
rect 43456 11694 43484 12242
rect 43444 11688 43496 11694
rect 43444 11630 43496 11636
rect 43260 11212 43312 11218
rect 43260 11154 43312 11160
rect 43260 6384 43312 6390
rect 43260 6326 43312 6332
rect 43168 5364 43220 5370
rect 43168 5306 43220 5312
rect 43076 5024 43128 5030
rect 43076 4966 43128 4972
rect 43088 4622 43116 4966
rect 43272 4758 43300 6326
rect 43444 6248 43496 6254
rect 43444 6190 43496 6196
rect 43456 6118 43484 6190
rect 43444 6112 43496 6118
rect 43444 6054 43496 6060
rect 43260 4752 43312 4758
rect 43260 4694 43312 4700
rect 43076 4616 43128 4622
rect 43076 4558 43128 4564
rect 43444 4616 43496 4622
rect 43444 4558 43496 4564
rect 42984 4548 43036 4554
rect 42984 4490 43036 4496
rect 42996 4146 43024 4490
rect 43352 4480 43404 4486
rect 43352 4422 43404 4428
rect 43364 4282 43392 4422
rect 43352 4276 43404 4282
rect 43352 4218 43404 4224
rect 42984 4140 43036 4146
rect 42984 4082 43036 4088
rect 42996 3398 43024 4082
rect 43456 4078 43484 4558
rect 43076 4072 43128 4078
rect 43076 4014 43128 4020
rect 43444 4072 43496 4078
rect 43444 4014 43496 4020
rect 42984 3392 43036 3398
rect 42984 3334 43036 3340
rect 42996 3058 43024 3334
rect 42984 3052 43036 3058
rect 42984 2994 43036 3000
rect 43088 2854 43116 4014
rect 43456 3534 43484 4014
rect 43444 3528 43496 3534
rect 43444 3470 43496 3476
rect 43168 3120 43220 3126
rect 43168 3062 43220 3068
rect 43076 2848 43128 2854
rect 43076 2790 43128 2796
rect 43180 800 43208 3062
rect 43260 3052 43312 3058
rect 43260 2994 43312 3000
rect 43272 2774 43300 2994
rect 43456 2990 43484 3470
rect 43444 2984 43496 2990
rect 43444 2926 43496 2932
rect 43272 2746 43392 2774
rect 43364 2446 43392 2746
rect 43352 2440 43404 2446
rect 43352 2382 43404 2388
rect 43548 2310 43576 12406
rect 43720 8900 43772 8906
rect 43720 8842 43772 8848
rect 43628 8560 43680 8566
rect 43628 8502 43680 8508
rect 43640 8362 43668 8502
rect 43628 8356 43680 8362
rect 43628 8298 43680 8304
rect 43640 7886 43668 8298
rect 43732 8090 43760 8842
rect 43824 8498 43852 20810
rect 43904 20460 43956 20466
rect 43904 20402 43956 20408
rect 43996 20460 44048 20466
rect 43996 20402 44048 20408
rect 43916 18970 43944 20402
rect 44008 20262 44036 20402
rect 43996 20256 44048 20262
rect 43996 20198 44048 20204
rect 43904 18964 43956 18970
rect 43904 18906 43956 18912
rect 43996 14272 44048 14278
rect 43996 14214 44048 14220
rect 44008 14074 44036 14214
rect 43996 14068 44048 14074
rect 43996 14010 44048 14016
rect 43996 11688 44048 11694
rect 43996 11630 44048 11636
rect 44008 10713 44036 11630
rect 43994 10704 44050 10713
rect 43994 10639 44050 10648
rect 43904 9580 43956 9586
rect 43904 9522 43956 9528
rect 43996 9580 44048 9586
rect 43996 9522 44048 9528
rect 43916 9110 43944 9522
rect 43904 9104 43956 9110
rect 43904 9046 43956 9052
rect 44008 8922 44036 9522
rect 43916 8894 44036 8922
rect 43916 8838 43944 8894
rect 43904 8832 43956 8838
rect 43904 8774 43956 8780
rect 43812 8492 43864 8498
rect 43812 8434 43864 8440
rect 43720 8084 43772 8090
rect 43720 8026 43772 8032
rect 43916 7954 43944 8774
rect 43904 7948 43956 7954
rect 43904 7890 43956 7896
rect 43628 7880 43680 7886
rect 43628 7822 43680 7828
rect 43996 7880 44048 7886
rect 43996 7822 44048 7828
rect 44008 7410 44036 7822
rect 43996 7404 44048 7410
rect 43996 7346 44048 7352
rect 43904 5364 43956 5370
rect 43904 5306 43956 5312
rect 43916 4622 43944 5306
rect 43904 4616 43956 4622
rect 43904 4558 43956 4564
rect 43996 4616 44048 4622
rect 43996 4558 44048 4564
rect 44008 4434 44036 4558
rect 43916 4406 44036 4434
rect 43628 3936 43680 3942
rect 43628 3878 43680 3884
rect 43640 3058 43668 3878
rect 43718 3632 43774 3641
rect 43718 3567 43774 3576
rect 43732 3534 43760 3567
rect 43720 3528 43772 3534
rect 43720 3470 43772 3476
rect 43916 3466 43944 4406
rect 43996 4072 44048 4078
rect 43996 4014 44048 4020
rect 43904 3460 43956 3466
rect 43904 3402 43956 3408
rect 43720 3392 43772 3398
rect 43720 3334 43772 3340
rect 43628 3052 43680 3058
rect 43628 2994 43680 3000
rect 43536 2304 43588 2310
rect 43536 2246 43588 2252
rect 43444 1148 43496 1154
rect 43444 1090 43496 1096
rect 43456 800 43484 1090
rect 43732 800 43760 3334
rect 43812 3052 43864 3058
rect 43812 2994 43864 3000
rect 43824 1290 43852 2994
rect 43904 2984 43956 2990
rect 43904 2926 43956 2932
rect 43916 2446 43944 2926
rect 43904 2440 43956 2446
rect 43904 2382 43956 2388
rect 43812 1284 43864 1290
rect 43812 1226 43864 1232
rect 44008 800 44036 4014
rect 44100 2650 44128 47670
rect 45744 44872 45796 44878
rect 45744 44814 45796 44820
rect 44364 34468 44416 34474
rect 44364 34410 44416 34416
rect 44180 18284 44232 18290
rect 44180 18226 44232 18232
rect 44192 16998 44220 18226
rect 44180 16992 44232 16998
rect 44180 16934 44232 16940
rect 44272 16652 44324 16658
rect 44272 16594 44324 16600
rect 44180 16108 44232 16114
rect 44180 16050 44232 16056
rect 44192 15434 44220 16050
rect 44180 15428 44232 15434
rect 44180 15370 44232 15376
rect 44192 11626 44220 15370
rect 44284 14822 44312 16594
rect 44272 14816 44324 14822
rect 44272 14758 44324 14764
rect 44180 11620 44232 11626
rect 44180 11562 44232 11568
rect 44192 10674 44220 11562
rect 44180 10668 44232 10674
rect 44180 10610 44232 10616
rect 44180 10056 44232 10062
rect 44180 9998 44232 10004
rect 44272 10056 44324 10062
rect 44272 9998 44324 10004
rect 44192 8906 44220 9998
rect 44284 9722 44312 9998
rect 44272 9716 44324 9722
rect 44272 9658 44324 9664
rect 44180 8900 44232 8906
rect 44180 8842 44232 8848
rect 44192 8634 44220 8842
rect 44180 8628 44232 8634
rect 44180 8570 44232 8576
rect 44180 5228 44232 5234
rect 44180 5170 44232 5176
rect 44192 3398 44220 5170
rect 44272 4140 44324 4146
rect 44272 4082 44324 4088
rect 44284 3738 44312 4082
rect 44272 3732 44324 3738
rect 44272 3674 44324 3680
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44376 3194 44404 34410
rect 45756 26234 45784 44814
rect 50068 41472 50120 41478
rect 50068 41414 50120 41420
rect 46848 38344 46900 38350
rect 46848 38286 46900 38292
rect 46480 30252 46532 30258
rect 46480 30194 46532 30200
rect 45664 26206 45784 26234
rect 44732 25764 44784 25770
rect 44732 25706 44784 25712
rect 44744 22094 44772 25706
rect 44652 22066 44772 22094
rect 44456 20596 44508 20602
rect 44456 20538 44508 20544
rect 44468 13734 44496 20538
rect 44548 14272 44600 14278
rect 44548 14214 44600 14220
rect 44456 13728 44508 13734
rect 44456 13670 44508 13676
rect 44468 11082 44496 13670
rect 44560 13394 44588 14214
rect 44548 13388 44600 13394
rect 44548 13330 44600 13336
rect 44456 11076 44508 11082
rect 44508 11036 44588 11064
rect 44456 11018 44508 11024
rect 44456 9648 44508 9654
rect 44456 9590 44508 9596
rect 44468 8974 44496 9590
rect 44560 8974 44588 11036
rect 44456 8968 44508 8974
rect 44456 8910 44508 8916
rect 44548 8968 44600 8974
rect 44548 8910 44600 8916
rect 44548 8492 44600 8498
rect 44548 8434 44600 8440
rect 44560 7478 44588 8434
rect 44548 7472 44600 7478
rect 44548 7414 44600 7420
rect 44548 5228 44600 5234
rect 44548 5170 44600 5176
rect 44456 4548 44508 4554
rect 44456 4490 44508 4496
rect 44364 3188 44416 3194
rect 44364 3130 44416 3136
rect 44468 2774 44496 4490
rect 44284 2746 44496 2774
rect 44088 2644 44140 2650
rect 44088 2586 44140 2592
rect 44180 2644 44232 2650
rect 44180 2586 44232 2592
rect 44192 2553 44220 2586
rect 44178 2544 44234 2553
rect 44178 2479 44234 2488
rect 44088 2440 44140 2446
rect 44088 2382 44140 2388
rect 44100 2106 44128 2382
rect 44088 2100 44140 2106
rect 44088 2042 44140 2048
rect 44284 800 44312 2746
rect 44560 800 44588 5170
rect 44652 3194 44680 22066
rect 45560 20936 45612 20942
rect 45560 20878 45612 20884
rect 44732 20528 44784 20534
rect 44732 20470 44784 20476
rect 44744 20058 44772 20470
rect 45376 20256 45428 20262
rect 45376 20198 45428 20204
rect 44732 20052 44784 20058
rect 44732 19994 44784 20000
rect 45388 19854 45416 20198
rect 45468 19916 45520 19922
rect 45468 19858 45520 19864
rect 45376 19848 45428 19854
rect 45376 19790 45428 19796
rect 45388 18766 45416 19790
rect 45480 19378 45508 19858
rect 45572 19718 45600 20878
rect 45560 19712 45612 19718
rect 45560 19654 45612 19660
rect 45468 19372 45520 19378
rect 45468 19314 45520 19320
rect 45376 18760 45428 18766
rect 45376 18702 45428 18708
rect 44732 18352 44784 18358
rect 44732 18294 44784 18300
rect 44744 8498 44772 18294
rect 45480 16250 45508 19314
rect 45560 16448 45612 16454
rect 45560 16390 45612 16396
rect 45468 16244 45520 16250
rect 45468 16186 45520 16192
rect 45284 15700 45336 15706
rect 45284 15642 45336 15648
rect 45192 10804 45244 10810
rect 45192 10746 45244 10752
rect 44824 10668 44876 10674
rect 44824 10610 44876 10616
rect 44836 9994 44864 10610
rect 44824 9988 44876 9994
rect 44824 9930 44876 9936
rect 45204 9586 45232 10746
rect 45100 9580 45152 9586
rect 45100 9522 45152 9528
rect 45192 9580 45244 9586
rect 45192 9522 45244 9528
rect 44916 9104 44968 9110
rect 44916 9046 44968 9052
rect 44928 8566 44956 9046
rect 44916 8560 44968 8566
rect 44916 8502 44968 8508
rect 44732 8492 44784 8498
rect 44732 8434 44784 8440
rect 44744 7886 44772 8434
rect 44732 7880 44784 7886
rect 44732 7822 44784 7828
rect 45112 7818 45140 9522
rect 45100 7812 45152 7818
rect 45100 7754 45152 7760
rect 45112 7342 45140 7754
rect 45100 7336 45152 7342
rect 45100 7278 45152 7284
rect 45008 5024 45060 5030
rect 45008 4966 45060 4972
rect 44824 4208 44876 4214
rect 44824 4150 44876 4156
rect 44732 3460 44784 3466
rect 44732 3402 44784 3408
rect 44640 3188 44692 3194
rect 44640 3130 44692 3136
rect 44744 1086 44772 3402
rect 44732 1080 44784 1086
rect 44732 1022 44784 1028
rect 44836 800 44864 4150
rect 44916 4140 44968 4146
rect 44916 4082 44968 4088
rect 44928 3126 44956 4082
rect 45020 3670 45048 4966
rect 45192 3936 45244 3942
rect 45192 3878 45244 3884
rect 45008 3664 45060 3670
rect 45008 3606 45060 3612
rect 45100 3664 45152 3670
rect 45100 3606 45152 3612
rect 44916 3120 44968 3126
rect 44916 3062 44968 3068
rect 45008 3052 45060 3058
rect 45008 2994 45060 3000
rect 45020 1222 45048 2994
rect 45008 1216 45060 1222
rect 45008 1158 45060 1164
rect 45112 800 45140 3606
rect 45204 2378 45232 3878
rect 45296 2990 45324 15642
rect 45468 11620 45520 11626
rect 45468 11562 45520 11568
rect 45480 11218 45508 11562
rect 45468 11212 45520 11218
rect 45468 11154 45520 11160
rect 45468 9920 45520 9926
rect 45468 9862 45520 9868
rect 45480 9654 45508 9862
rect 45468 9648 45520 9654
rect 45468 9590 45520 9596
rect 45376 8424 45428 8430
rect 45376 8366 45428 8372
rect 45388 7410 45416 8366
rect 45376 7404 45428 7410
rect 45376 7346 45428 7352
rect 45468 7200 45520 7206
rect 45468 7142 45520 7148
rect 45480 4758 45508 7142
rect 45468 4752 45520 4758
rect 45468 4694 45520 4700
rect 45572 3738 45600 16390
rect 45664 12434 45692 26206
rect 46296 19848 46348 19854
rect 46296 19790 46348 19796
rect 45928 19712 45980 19718
rect 45928 19654 45980 19660
rect 45940 19514 45968 19654
rect 45928 19508 45980 19514
rect 45928 19450 45980 19456
rect 45744 19372 45796 19378
rect 45744 19314 45796 19320
rect 45756 18970 45784 19314
rect 46308 18970 46336 19790
rect 45744 18964 45796 18970
rect 45744 18906 45796 18912
rect 46296 18964 46348 18970
rect 46296 18906 46348 18912
rect 46020 18760 46072 18766
rect 46020 18702 46072 18708
rect 46032 18426 46060 18702
rect 46112 18624 46164 18630
rect 46112 18566 46164 18572
rect 46020 18420 46072 18426
rect 46020 18362 46072 18368
rect 46124 18358 46152 18566
rect 46112 18352 46164 18358
rect 46112 18294 46164 18300
rect 45926 16688 45982 16697
rect 45926 16623 45982 16632
rect 45664 12406 45784 12434
rect 45652 5228 45704 5234
rect 45652 5170 45704 5176
rect 45560 3732 45612 3738
rect 45560 3674 45612 3680
rect 45376 3460 45428 3466
rect 45376 3402 45428 3408
rect 45284 2984 45336 2990
rect 45284 2926 45336 2932
rect 45192 2372 45244 2378
rect 45192 2314 45244 2320
rect 45284 2372 45336 2378
rect 45284 2314 45336 2320
rect 45296 1018 45324 2314
rect 45284 1012 45336 1018
rect 45284 954 45336 960
rect 45388 800 45416 3402
rect 45664 800 45692 5170
rect 45756 2774 45784 12406
rect 45940 8514 45968 16623
rect 46388 16516 46440 16522
rect 46388 16458 46440 16464
rect 46400 16250 46428 16458
rect 46388 16244 46440 16250
rect 46388 16186 46440 16192
rect 46204 14884 46256 14890
rect 46204 14826 46256 14832
rect 46216 14006 46244 14826
rect 46204 14000 46256 14006
rect 46204 13942 46256 13948
rect 46296 12436 46348 12442
rect 46296 12378 46348 12384
rect 46308 11762 46336 12378
rect 46388 12096 46440 12102
rect 46388 12038 46440 12044
rect 46296 11756 46348 11762
rect 46296 11698 46348 11704
rect 46204 11552 46256 11558
rect 46204 11494 46256 11500
rect 46296 11552 46348 11558
rect 46296 11494 46348 11500
rect 46216 11354 46244 11494
rect 46204 11348 46256 11354
rect 46204 11290 46256 11296
rect 46308 11082 46336 11494
rect 46296 11076 46348 11082
rect 46296 11018 46348 11024
rect 46400 10198 46428 12038
rect 46388 10192 46440 10198
rect 46388 10134 46440 10140
rect 46112 10056 46164 10062
rect 46112 9998 46164 10004
rect 46124 8974 46152 9998
rect 46296 9920 46348 9926
rect 46296 9862 46348 9868
rect 46204 9376 46256 9382
rect 46204 9318 46256 9324
rect 46112 8968 46164 8974
rect 46112 8910 46164 8916
rect 46124 8634 46152 8910
rect 46216 8634 46244 9318
rect 46308 8974 46336 9862
rect 46296 8968 46348 8974
rect 46296 8910 46348 8916
rect 46112 8628 46164 8634
rect 46112 8570 46164 8576
rect 46204 8628 46256 8634
rect 46204 8570 46256 8576
rect 46308 8514 46336 8910
rect 46400 8616 46428 10134
rect 46492 9382 46520 30194
rect 46756 20460 46808 20466
rect 46756 20402 46808 20408
rect 46572 18760 46624 18766
rect 46572 18702 46624 18708
rect 46664 18760 46716 18766
rect 46664 18702 46716 18708
rect 46584 18222 46612 18702
rect 46572 18216 46624 18222
rect 46572 18158 46624 18164
rect 46572 16448 46624 16454
rect 46572 16390 46624 16396
rect 46584 16250 46612 16390
rect 46572 16244 46624 16250
rect 46572 16186 46624 16192
rect 46584 16153 46612 16186
rect 46570 16144 46626 16153
rect 46570 16079 46626 16088
rect 46572 13320 46624 13326
rect 46572 13262 46624 13268
rect 46584 10130 46612 13262
rect 46676 11082 46704 18702
rect 46768 16658 46796 20402
rect 46860 19514 46888 38286
rect 47676 35624 47728 35630
rect 47676 35566 47728 35572
rect 47584 34536 47636 34542
rect 47584 34478 47636 34484
rect 47492 31204 47544 31210
rect 47492 31146 47544 31152
rect 47400 28416 47452 28422
rect 47400 28358 47452 28364
rect 47032 25696 47084 25702
rect 47032 25638 47084 25644
rect 46940 20392 46992 20398
rect 46940 20334 46992 20340
rect 46952 19514 46980 20334
rect 46848 19508 46900 19514
rect 46848 19450 46900 19456
rect 46940 19508 46992 19514
rect 46940 19450 46992 19456
rect 46860 18358 46888 19450
rect 46952 18630 46980 19450
rect 46940 18624 46992 18630
rect 46940 18566 46992 18572
rect 46848 18352 46900 18358
rect 46848 18294 46900 18300
rect 46952 17610 46980 18566
rect 46940 17604 46992 17610
rect 46940 17546 46992 17552
rect 46756 16652 46808 16658
rect 46756 16594 46808 16600
rect 46768 11778 46796 16594
rect 46848 15904 46900 15910
rect 46848 15846 46900 15852
rect 46860 14890 46888 15846
rect 46848 14884 46900 14890
rect 46848 14826 46900 14832
rect 46860 12102 46888 14826
rect 46848 12096 46900 12102
rect 46848 12038 46900 12044
rect 46860 11914 46888 12038
rect 46860 11886 46980 11914
rect 46768 11750 46888 11778
rect 46756 11688 46808 11694
rect 46756 11630 46808 11636
rect 46768 11286 46796 11630
rect 46756 11280 46808 11286
rect 46756 11222 46808 11228
rect 46664 11076 46716 11082
rect 46664 11018 46716 11024
rect 46572 10124 46624 10130
rect 46572 10066 46624 10072
rect 46584 9722 46612 10066
rect 46572 9716 46624 9722
rect 46572 9658 46624 9664
rect 46480 9376 46532 9382
rect 46480 9318 46532 9324
rect 46676 8838 46704 11018
rect 46754 9072 46810 9081
rect 46754 9007 46810 9016
rect 46664 8832 46716 8838
rect 46664 8774 46716 8780
rect 46400 8588 46520 8616
rect 45940 8486 46152 8514
rect 46124 8430 46152 8486
rect 46216 8486 46336 8514
rect 46388 8492 46440 8498
rect 46112 8424 46164 8430
rect 46112 8366 46164 8372
rect 46124 7886 46152 8366
rect 46112 7880 46164 7886
rect 46112 7822 46164 7828
rect 45836 7200 45888 7206
rect 45836 7142 45888 7148
rect 45848 6730 45876 7142
rect 46124 7002 46152 7822
rect 46112 6996 46164 7002
rect 46112 6938 46164 6944
rect 46216 6882 46244 8486
rect 46388 8434 46440 8440
rect 46296 8288 46348 8294
rect 46296 8230 46348 8236
rect 46308 7410 46336 8230
rect 46400 8090 46428 8434
rect 46388 8084 46440 8090
rect 46388 8026 46440 8032
rect 46492 7954 46520 8588
rect 46480 7948 46532 7954
rect 46480 7890 46532 7896
rect 46296 7404 46348 7410
rect 46296 7346 46348 7352
rect 46308 7002 46336 7346
rect 46492 7342 46520 7890
rect 46572 7812 46624 7818
rect 46572 7754 46624 7760
rect 46480 7336 46532 7342
rect 46480 7278 46532 7284
rect 46296 6996 46348 7002
rect 46296 6938 46348 6944
rect 46216 6854 46428 6882
rect 45836 6724 45888 6730
rect 45836 6666 45888 6672
rect 46400 6322 46428 6854
rect 46388 6316 46440 6322
rect 46388 6258 46440 6264
rect 45926 5400 45982 5409
rect 45926 5335 45982 5344
rect 45940 4146 45968 5335
rect 46020 4548 46072 4554
rect 46020 4490 46072 4496
rect 45928 4140 45980 4146
rect 45928 4082 45980 4088
rect 46032 3670 46060 4490
rect 46400 4078 46428 6258
rect 46584 6254 46612 7754
rect 46572 6248 46624 6254
rect 46572 6190 46624 6196
rect 46584 5166 46612 6190
rect 46572 5160 46624 5166
rect 46572 5102 46624 5108
rect 46768 4146 46796 9007
rect 46860 6866 46888 11750
rect 46952 11694 46980 11886
rect 46940 11688 46992 11694
rect 46940 11630 46992 11636
rect 46940 11144 46992 11150
rect 46940 11086 46992 11092
rect 46952 9926 46980 11086
rect 46940 9920 46992 9926
rect 46940 9862 46992 9868
rect 46848 6860 46900 6866
rect 46848 6802 46900 6808
rect 46860 6390 46888 6802
rect 46952 6798 46980 9862
rect 46940 6792 46992 6798
rect 46940 6734 46992 6740
rect 46848 6384 46900 6390
rect 46848 6326 46900 6332
rect 46952 5234 46980 6734
rect 46940 5228 46992 5234
rect 46940 5170 46992 5176
rect 46756 4140 46808 4146
rect 46756 4082 46808 4088
rect 46388 4072 46440 4078
rect 46388 4014 46440 4020
rect 47044 3738 47072 25638
rect 47124 18284 47176 18290
rect 47124 18226 47176 18232
rect 47136 18193 47164 18226
rect 47122 18184 47178 18193
rect 47122 18119 47178 18128
rect 47124 9376 47176 9382
rect 47124 9318 47176 9324
rect 47032 3732 47084 3738
rect 47032 3674 47084 3680
rect 46020 3664 46072 3670
rect 46020 3606 46072 3612
rect 46112 3528 46164 3534
rect 46112 3470 46164 3476
rect 45756 2746 45876 2774
rect 45848 2650 45876 2746
rect 45836 2644 45888 2650
rect 45836 2586 45888 2592
rect 45928 2372 45980 2378
rect 45928 2314 45980 2320
rect 45940 800 45968 2314
rect 46124 1154 46152 3470
rect 46756 3460 46808 3466
rect 46756 3402 46808 3408
rect 46204 3052 46256 3058
rect 46204 2994 46256 3000
rect 46112 1148 46164 1154
rect 46112 1090 46164 1096
rect 46216 800 46244 2994
rect 46296 2372 46348 2378
rect 46296 2314 46348 2320
rect 46308 950 46336 2314
rect 46296 944 46348 950
rect 46296 886 46348 892
rect 46480 944 46532 950
rect 46480 886 46532 892
rect 46492 800 46520 886
rect 46768 800 46796 3402
rect 47136 3126 47164 9318
rect 47124 3120 47176 3126
rect 47124 3062 47176 3068
rect 47032 3052 47084 3058
rect 47032 2994 47084 3000
rect 47044 800 47072 2994
rect 47412 2650 47440 28358
rect 47504 3194 47532 31146
rect 47596 20058 47624 34478
rect 47688 24886 47716 35566
rect 48964 31816 49016 31822
rect 48964 31758 49016 31764
rect 48872 29708 48924 29714
rect 48872 29650 48924 29656
rect 48780 26784 48832 26790
rect 48780 26726 48832 26732
rect 47676 24880 47728 24886
rect 47676 24822 47728 24828
rect 48412 24880 48464 24886
rect 48412 24822 48464 24828
rect 48424 22094 48452 24822
rect 48424 22066 48636 22094
rect 47860 20936 47912 20942
rect 47860 20878 47912 20884
rect 47676 20868 47728 20874
rect 47676 20810 47728 20816
rect 47688 20398 47716 20810
rect 47676 20392 47728 20398
rect 47676 20334 47728 20340
rect 47584 20052 47636 20058
rect 47584 19994 47636 20000
rect 47596 18698 47624 19994
rect 47872 19446 47900 20878
rect 48320 20800 48372 20806
rect 48320 20742 48372 20748
rect 48228 20392 48280 20398
rect 48228 20334 48280 20340
rect 48240 19922 48268 20334
rect 48228 19916 48280 19922
rect 48228 19858 48280 19864
rect 47860 19440 47912 19446
rect 47860 19382 47912 19388
rect 48136 19440 48188 19446
rect 48136 19382 48188 19388
rect 47676 19372 47728 19378
rect 47676 19314 47728 19320
rect 47584 18692 47636 18698
rect 47584 18634 47636 18640
rect 47688 18630 47716 19314
rect 47766 18728 47822 18737
rect 47766 18663 47768 18672
rect 47820 18663 47822 18672
rect 47768 18634 47820 18640
rect 47676 18624 47728 18630
rect 47676 18566 47728 18572
rect 47688 16522 47716 18566
rect 48148 18222 48176 19382
rect 48240 18442 48268 19858
rect 48332 19854 48360 20742
rect 48504 20460 48556 20466
rect 48504 20402 48556 20408
rect 48412 20256 48464 20262
rect 48412 20198 48464 20204
rect 48424 19990 48452 20198
rect 48516 20058 48544 20402
rect 48504 20052 48556 20058
rect 48504 19994 48556 20000
rect 48412 19984 48464 19990
rect 48412 19926 48464 19932
rect 48320 19848 48372 19854
rect 48320 19790 48372 19796
rect 48424 18766 48452 19926
rect 48504 18964 48556 18970
rect 48504 18906 48556 18912
rect 48412 18760 48464 18766
rect 48412 18702 48464 18708
rect 48240 18426 48360 18442
rect 48240 18420 48372 18426
rect 48240 18414 48320 18420
rect 48136 18216 48188 18222
rect 48136 18158 48188 18164
rect 48148 17746 48176 18158
rect 48136 17740 48188 17746
rect 48136 17682 48188 17688
rect 47952 17672 48004 17678
rect 47952 17614 48004 17620
rect 47964 17202 47992 17614
rect 47952 17196 48004 17202
rect 47952 17138 48004 17144
rect 47676 16516 47728 16522
rect 47676 16458 47728 16464
rect 47860 16108 47912 16114
rect 47860 16050 47912 16056
rect 47768 16040 47820 16046
rect 47768 15982 47820 15988
rect 47780 11150 47808 15982
rect 47872 15162 47900 16050
rect 48136 15904 48188 15910
rect 48136 15846 48188 15852
rect 48148 15348 48176 15846
rect 48240 15706 48268 18414
rect 48320 18362 48372 18368
rect 48516 18290 48544 18906
rect 48504 18284 48556 18290
rect 48504 18226 48556 18232
rect 48228 15700 48280 15706
rect 48228 15642 48280 15648
rect 48240 15502 48268 15642
rect 48228 15496 48280 15502
rect 48228 15438 48280 15444
rect 48148 15320 48268 15348
rect 47860 15156 47912 15162
rect 47860 15098 47912 15104
rect 48240 14958 48268 15320
rect 48412 15088 48464 15094
rect 48412 15030 48464 15036
rect 48228 14952 48280 14958
rect 48228 14894 48280 14900
rect 47768 11144 47820 11150
rect 47768 11086 47820 11092
rect 48240 8129 48268 14894
rect 48320 11756 48372 11762
rect 48320 11698 48372 11704
rect 48226 8120 48282 8129
rect 48226 8055 48282 8064
rect 48136 4140 48188 4146
rect 48136 4082 48188 4088
rect 47952 4004 48004 4010
rect 47952 3946 48004 3952
rect 47964 3738 47992 3946
rect 47952 3732 48004 3738
rect 47952 3674 48004 3680
rect 47584 3528 47636 3534
rect 47584 3470 47636 3476
rect 47492 3188 47544 3194
rect 47492 3130 47544 3136
rect 47400 2644 47452 2650
rect 47400 2586 47452 2592
rect 47400 2372 47452 2378
rect 47400 2314 47452 2320
rect 47216 2304 47268 2310
rect 47216 2246 47268 2252
rect 47228 2038 47256 2246
rect 47216 2032 47268 2038
rect 47216 1974 47268 1980
rect 47308 1012 47360 1018
rect 47308 954 47360 960
rect 47320 800 47348 954
rect 47412 950 47440 2314
rect 47400 944 47452 950
rect 47400 886 47452 892
rect 47596 800 47624 3470
rect 47872 882 47992 898
rect 47872 876 48004 882
rect 47872 870 47952 876
rect 47872 800 47900 870
rect 47952 818 48004 824
rect 48148 800 48176 4082
rect 48332 3670 48360 11698
rect 48424 4010 48452 15030
rect 48412 4004 48464 4010
rect 48412 3946 48464 3952
rect 48608 3738 48636 22066
rect 48688 18760 48740 18766
rect 48688 18702 48740 18708
rect 48700 17814 48728 18702
rect 48688 17808 48740 17814
rect 48688 17750 48740 17756
rect 48596 3732 48648 3738
rect 48596 3674 48648 3680
rect 48320 3664 48372 3670
rect 48320 3606 48372 3612
rect 48688 3528 48740 3534
rect 48688 3470 48740 3476
rect 48412 3052 48464 3058
rect 48412 2994 48464 3000
rect 48424 800 48452 2994
rect 48700 800 48728 3470
rect 48792 3194 48820 26726
rect 48780 3188 48832 3194
rect 48780 3130 48832 3136
rect 48884 2650 48912 29650
rect 48976 20874 49004 31758
rect 50080 28994 50108 41414
rect 49988 28966 50108 28994
rect 49792 28484 49844 28490
rect 49792 28426 49844 28432
rect 49056 21344 49108 21350
rect 49056 21286 49108 21292
rect 48964 20868 49016 20874
rect 48964 20810 49016 20816
rect 48964 18624 49016 18630
rect 48964 18566 49016 18572
rect 48976 18290 49004 18566
rect 48964 18284 49016 18290
rect 48964 18226 49016 18232
rect 49068 14414 49096 21286
rect 49608 20868 49660 20874
rect 49608 20810 49660 20816
rect 49620 20602 49648 20810
rect 49608 20596 49660 20602
rect 49608 20538 49660 20544
rect 49240 20392 49292 20398
rect 49240 20334 49292 20340
rect 49252 19990 49280 20334
rect 49240 19984 49292 19990
rect 49240 19926 49292 19932
rect 49700 19508 49752 19514
rect 49804 19496 49832 28426
rect 49804 19468 49924 19496
rect 49700 19450 49752 19456
rect 49712 19417 49740 19450
rect 49698 19408 49754 19417
rect 49698 19343 49754 19352
rect 49792 19372 49844 19378
rect 49792 19314 49844 19320
rect 49700 19236 49752 19242
rect 49700 19178 49752 19184
rect 49712 19145 49740 19178
rect 49698 19136 49754 19145
rect 49698 19071 49754 19080
rect 49804 18834 49832 19314
rect 49792 18828 49844 18834
rect 49792 18770 49844 18776
rect 49056 14408 49108 14414
rect 49056 14350 49108 14356
rect 49424 7744 49476 7750
rect 49424 7686 49476 7692
rect 49436 3738 49464 7686
rect 49608 6860 49660 6866
rect 49608 6802 49660 6808
rect 49620 4690 49648 6802
rect 49608 4684 49660 4690
rect 49608 4626 49660 4632
rect 49424 3732 49476 3738
rect 49424 3674 49476 3680
rect 49792 3460 49844 3466
rect 49792 3402 49844 3408
rect 49516 3120 49568 3126
rect 49516 3062 49568 3068
rect 48964 3052 49016 3058
rect 48964 2994 49016 3000
rect 48872 2644 48924 2650
rect 48872 2586 48924 2592
rect 48780 2372 48832 2378
rect 48780 2314 48832 2320
rect 48792 1018 48820 2314
rect 48780 1012 48832 1018
rect 48780 954 48832 960
rect 48976 800 49004 2994
rect 49240 944 49292 950
rect 49240 886 49292 892
rect 49252 800 49280 886
rect 49528 800 49556 3062
rect 49700 2848 49752 2854
rect 49700 2790 49752 2796
rect 49712 2650 49740 2790
rect 49700 2644 49752 2650
rect 49700 2586 49752 2592
rect 49700 2372 49752 2378
rect 49700 2314 49752 2320
rect 49712 882 49740 2314
rect 49700 876 49752 882
rect 49700 818 49752 824
rect 49804 800 49832 3402
rect 49896 3194 49924 19468
rect 49988 18426 50016 28966
rect 50172 24154 50200 51046
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 53484 39370 53512 61066
rect 54300 61056 54352 61062
rect 54300 60998 54352 61004
rect 53840 43784 53892 43790
rect 53840 43726 53892 43732
rect 53564 41608 53616 41614
rect 53564 41550 53616 41556
rect 53472 39364 53524 39370
rect 53472 39306 53524 39312
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 53472 37256 53524 37262
rect 53472 37198 53524 37204
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 53484 36650 53512 37198
rect 53472 36644 53524 36650
rect 53472 36586 53524 36592
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 53288 32496 53340 32502
rect 53288 32438 53340 32444
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 52552 25288 52604 25294
rect 52552 25230 52604 25236
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50080 24126 50200 24154
rect 51816 24132 51868 24138
rect 50080 18698 50108 24126
rect 51816 24074 51868 24080
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 51828 22094 51856 24074
rect 51736 22066 51856 22094
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50160 20460 50212 20466
rect 50160 20402 50212 20408
rect 51632 20460 51684 20466
rect 51632 20402 51684 20408
rect 50172 19174 50200 20402
rect 51448 20392 51500 20398
rect 51448 20334 51500 20340
rect 50528 20256 50580 20262
rect 50528 20198 50580 20204
rect 50540 19786 50568 20198
rect 50620 20052 50672 20058
rect 50620 19994 50672 20000
rect 50528 19780 50580 19786
rect 50528 19722 50580 19728
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50528 19440 50580 19446
rect 50528 19382 50580 19388
rect 50160 19168 50212 19174
rect 50436 19168 50488 19174
rect 50160 19110 50212 19116
rect 50434 19136 50436 19145
rect 50488 19136 50490 19145
rect 50434 19071 50490 19080
rect 50540 18970 50568 19382
rect 50632 19310 50660 19994
rect 51264 19440 51316 19446
rect 51262 19408 51264 19417
rect 51316 19408 51318 19417
rect 51262 19343 51318 19352
rect 50620 19304 50672 19310
rect 50620 19246 50672 19252
rect 50988 19304 51040 19310
rect 50988 19246 51040 19252
rect 50528 18964 50580 18970
rect 50528 18906 50580 18912
rect 50068 18692 50120 18698
rect 50068 18634 50120 18640
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 49976 18420 50028 18426
rect 49976 18362 50028 18368
rect 49988 17610 50016 18362
rect 51000 17678 51028 19246
rect 51460 19242 51488 20334
rect 51644 19514 51672 20402
rect 51632 19508 51684 19514
rect 51632 19450 51684 19456
rect 51448 19236 51500 19242
rect 51448 19178 51500 19184
rect 50988 17672 51040 17678
rect 50988 17614 51040 17620
rect 49976 17604 50028 17610
rect 49976 17546 50028 17552
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50712 16108 50764 16114
rect 50712 16050 50764 16056
rect 50724 15910 50752 16050
rect 51000 16046 51028 17614
rect 51080 17536 51132 17542
rect 51080 17478 51132 17484
rect 51092 16250 51120 17478
rect 51460 17202 51488 19178
rect 51632 17672 51684 17678
rect 51552 17632 51632 17660
rect 51448 17196 51500 17202
rect 51448 17138 51500 17144
rect 51552 16726 51580 17632
rect 51632 17614 51684 17620
rect 51632 17536 51684 17542
rect 51632 17478 51684 17484
rect 51644 17202 51672 17478
rect 51632 17196 51684 17202
rect 51632 17138 51684 17144
rect 51540 16720 51592 16726
rect 51540 16662 51592 16668
rect 51552 16266 51580 16662
rect 51632 16584 51684 16590
rect 51632 16526 51684 16532
rect 51080 16244 51132 16250
rect 51080 16186 51132 16192
rect 51460 16238 51580 16266
rect 51644 16250 51672 16526
rect 51632 16244 51684 16250
rect 51172 16176 51224 16182
rect 51172 16118 51224 16124
rect 50988 16040 51040 16046
rect 50988 15982 51040 15988
rect 50712 15904 50764 15910
rect 50712 15846 50764 15852
rect 50724 15366 50752 15846
rect 51184 15366 51212 16118
rect 51356 16108 51408 16114
rect 51356 16050 51408 16056
rect 51368 15706 51396 16050
rect 51356 15700 51408 15706
rect 51356 15642 51408 15648
rect 51460 15502 51488 16238
rect 51632 16186 51684 16192
rect 51540 16176 51592 16182
rect 51540 16118 51592 16124
rect 51552 15910 51580 16118
rect 51540 15904 51592 15910
rect 51540 15846 51592 15852
rect 51448 15496 51500 15502
rect 51448 15438 51500 15444
rect 50712 15360 50764 15366
rect 50712 15302 50764 15308
rect 51172 15360 51224 15366
rect 51172 15302 51224 15308
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50160 14816 50212 14822
rect 50160 14758 50212 14764
rect 50172 3738 50200 14758
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 51736 12434 51764 22066
rect 52368 20324 52420 20330
rect 52368 20266 52420 20272
rect 52380 19922 52408 20266
rect 52460 20256 52512 20262
rect 52460 20198 52512 20204
rect 52368 19916 52420 19922
rect 52368 19858 52420 19864
rect 52472 19854 52500 20198
rect 52460 19848 52512 19854
rect 52460 19790 52512 19796
rect 52368 19780 52420 19786
rect 52368 19722 52420 19728
rect 52380 19666 52408 19722
rect 52564 19666 52592 25230
rect 52920 20936 52972 20942
rect 52920 20878 52972 20884
rect 52644 20800 52696 20806
rect 52644 20742 52696 20748
rect 52380 19638 52592 19666
rect 52656 19281 52684 20742
rect 52642 19272 52698 19281
rect 52642 19207 52698 19216
rect 52368 18692 52420 18698
rect 52368 18634 52420 18640
rect 52092 18080 52144 18086
rect 52092 18022 52144 18028
rect 51908 17604 51960 17610
rect 51908 17546 51960 17552
rect 51920 17338 51948 17546
rect 51908 17332 51960 17338
rect 51908 17274 51960 17280
rect 51816 17128 51868 17134
rect 51816 17070 51868 17076
rect 51828 16658 51856 17070
rect 51816 16652 51868 16658
rect 51816 16594 51868 16600
rect 51816 16448 51868 16454
rect 51816 16390 51868 16396
rect 51828 15434 51856 16390
rect 51816 15428 51868 15434
rect 51816 15370 51868 15376
rect 52104 12434 52132 18022
rect 52380 14618 52408 18634
rect 52932 16794 52960 20878
rect 53012 17876 53064 17882
rect 53012 17818 53064 17824
rect 53024 17678 53052 17818
rect 53012 17672 53064 17678
rect 53012 17614 53064 17620
rect 52920 16788 52972 16794
rect 52920 16730 52972 16736
rect 52932 16454 52960 16730
rect 52920 16448 52972 16454
rect 52920 16390 52972 16396
rect 52932 16114 52960 16390
rect 52920 16108 52972 16114
rect 52920 16050 52972 16056
rect 53104 16108 53156 16114
rect 53104 16050 53156 16056
rect 53196 16108 53248 16114
rect 53196 16050 53248 16056
rect 53116 15706 53144 16050
rect 53104 15700 53156 15706
rect 53104 15642 53156 15648
rect 52368 14612 52420 14618
rect 52368 14554 52420 14560
rect 51736 12406 51856 12434
rect 52104 12406 52224 12434
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 51080 5024 51132 5030
rect 51080 4966 51132 4972
rect 51092 4622 51120 4966
rect 51356 4752 51408 4758
rect 51356 4694 51408 4700
rect 51080 4616 51132 4622
rect 51080 4558 51132 4564
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 51368 3738 51396 4694
rect 50160 3732 50212 3738
rect 50160 3674 50212 3680
rect 51356 3732 51408 3738
rect 51356 3674 51408 3680
rect 51264 3528 51316 3534
rect 51264 3470 51316 3476
rect 50620 3460 50672 3466
rect 50620 3402 50672 3408
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 49884 3188 49936 3194
rect 49884 3130 49936 3136
rect 50160 2848 50212 2854
rect 50160 2790 50212 2796
rect 50172 1442 50200 2790
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50172 1414 50384 1442
rect 50068 1012 50120 1018
rect 50068 954 50120 960
rect 50080 800 50108 954
rect 50356 800 50384 1414
rect 50632 800 50660 3402
rect 51080 3392 51132 3398
rect 51080 3334 51132 3340
rect 50896 3120 50948 3126
rect 50896 3062 50948 3068
rect 50908 800 50936 3062
rect 50988 3052 51040 3058
rect 50988 2994 51040 3000
rect 51000 2854 51028 2994
rect 50988 2848 51040 2854
rect 50988 2790 51040 2796
rect 51092 2582 51120 3334
rect 51080 2576 51132 2582
rect 51080 2518 51132 2524
rect 51080 2372 51132 2378
rect 51080 2314 51132 2320
rect 51092 950 51120 2314
rect 51276 1714 51304 3470
rect 51724 3460 51776 3466
rect 51724 3402 51776 3408
rect 51448 3052 51500 3058
rect 51448 2994 51500 3000
rect 51184 1686 51304 1714
rect 51080 944 51132 950
rect 51080 886 51132 892
rect 51184 800 51212 1686
rect 51460 800 51488 2994
rect 51736 800 51764 3402
rect 51828 2514 51856 12406
rect 52092 11552 52144 11558
rect 52092 11494 52144 11500
rect 52000 4208 52052 4214
rect 52000 4150 52052 4156
rect 51816 2508 51868 2514
rect 51816 2450 51868 2456
rect 51908 2372 51960 2378
rect 51908 2314 51960 2320
rect 51920 1018 51948 2314
rect 51908 1012 51960 1018
rect 51908 954 51960 960
rect 52012 800 52040 4150
rect 52104 2990 52132 11494
rect 52196 3194 52224 12406
rect 52368 10056 52420 10062
rect 52368 9998 52420 10004
rect 52380 9178 52408 9998
rect 52368 9172 52420 9178
rect 52368 9114 52420 9120
rect 52276 8900 52328 8906
rect 52276 8842 52328 8848
rect 52288 7818 52316 8842
rect 52368 8832 52420 8838
rect 52368 8774 52420 8780
rect 52380 8537 52408 8774
rect 52366 8528 52422 8537
rect 52366 8463 52422 8472
rect 53116 8430 53144 15642
rect 53208 15502 53236 16050
rect 53196 15496 53248 15502
rect 53196 15438 53248 15444
rect 53196 12436 53248 12442
rect 53196 12378 53248 12384
rect 53208 11150 53236 12378
rect 53196 11144 53248 11150
rect 53196 11086 53248 11092
rect 53104 8424 53156 8430
rect 53104 8366 53156 8372
rect 52276 7812 52328 7818
rect 52276 7754 52328 7760
rect 52276 7268 52328 7274
rect 52276 7210 52328 7216
rect 52288 4078 52316 7210
rect 52366 6216 52422 6225
rect 52366 6151 52422 6160
rect 52380 4146 52408 6151
rect 53104 5364 53156 5370
rect 53104 5306 53156 5312
rect 53116 4282 53144 5306
rect 53104 4276 53156 4282
rect 53104 4218 53156 4224
rect 52828 4208 52880 4214
rect 52828 4150 52880 4156
rect 52368 4140 52420 4146
rect 52368 4082 52420 4088
rect 52276 4072 52328 4078
rect 52276 4014 52328 4020
rect 52276 3936 52328 3942
rect 52276 3878 52328 3884
rect 52288 3602 52316 3878
rect 52276 3596 52328 3602
rect 52276 3538 52328 3544
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 52184 3188 52236 3194
rect 52184 3130 52236 3136
rect 52092 2984 52144 2990
rect 52092 2926 52144 2932
rect 52380 1714 52408 3334
rect 52458 2408 52514 2417
rect 52458 2343 52514 2352
rect 52552 2372 52604 2378
rect 52472 2310 52500 2343
rect 52552 2314 52604 2320
rect 52460 2304 52512 2310
rect 52460 2246 52512 2252
rect 52288 1686 52408 1714
rect 52288 800 52316 1686
rect 52564 800 52592 2314
rect 52840 800 52868 4150
rect 53104 3528 53156 3534
rect 53104 3470 53156 3476
rect 53116 800 53144 3470
rect 53300 3126 53328 32438
rect 53380 21072 53432 21078
rect 53378 21040 53380 21049
rect 53432 21040 53434 21049
rect 53378 20975 53434 20984
rect 53484 12374 53512 36586
rect 53576 20058 53604 41550
rect 53852 41478 53880 43726
rect 54312 42634 54340 60998
rect 54680 60722 54708 63294
rect 55310 63294 55536 63322
rect 55310 63200 55366 63294
rect 55508 61198 55536 63294
rect 56046 63200 56102 64000
rect 56782 63322 56838 64000
rect 56782 63294 56916 63322
rect 56782 63200 56838 63294
rect 56060 61198 56088 63200
rect 56692 61260 56744 61266
rect 56692 61202 56744 61208
rect 55496 61192 55548 61198
rect 55496 61134 55548 61140
rect 56048 61192 56100 61198
rect 56048 61134 56100 61140
rect 55772 61124 55824 61130
rect 55772 61066 55824 61072
rect 54668 60716 54720 60722
rect 54668 60658 54720 60664
rect 54852 60512 54904 60518
rect 54852 60454 54904 60460
rect 55588 60512 55640 60518
rect 55588 60454 55640 60460
rect 54864 43314 54892 60454
rect 55600 59770 55628 60454
rect 55588 59764 55640 59770
rect 55588 59706 55640 59712
rect 54852 43308 54904 43314
rect 54852 43250 54904 43256
rect 54300 42628 54352 42634
rect 54300 42570 54352 42576
rect 53840 41472 53892 41478
rect 53840 41414 53892 41420
rect 54668 40520 54720 40526
rect 54668 40462 54720 40468
rect 53748 37256 53800 37262
rect 53748 37198 53800 37204
rect 54484 37256 54536 37262
rect 54484 37198 54536 37204
rect 53656 36780 53708 36786
rect 53656 36722 53708 36728
rect 53564 20052 53616 20058
rect 53564 19994 53616 20000
rect 53576 19446 53604 19994
rect 53564 19440 53616 19446
rect 53564 19382 53616 19388
rect 53472 12368 53524 12374
rect 53472 12310 53524 12316
rect 53484 11150 53512 12310
rect 53564 12300 53616 12306
rect 53564 12242 53616 12248
rect 53576 11286 53604 12242
rect 53564 11280 53616 11286
rect 53564 11222 53616 11228
rect 53472 11144 53524 11150
rect 53472 11086 53524 11092
rect 53380 4208 53432 4214
rect 53380 4150 53432 4156
rect 53288 3120 53340 3126
rect 53288 3062 53340 3068
rect 53392 800 53420 4150
rect 53668 4010 53696 36722
rect 53760 4570 53788 37198
rect 53840 37188 53892 37194
rect 53840 37130 53892 37136
rect 53852 36786 53880 37130
rect 53840 36780 53892 36786
rect 53840 36722 53892 36728
rect 53852 35894 53880 36722
rect 54208 36576 54260 36582
rect 54208 36518 54260 36524
rect 54220 36378 54248 36518
rect 54208 36372 54260 36378
rect 54208 36314 54260 36320
rect 53852 35866 54432 35894
rect 54024 32564 54076 32570
rect 54024 32506 54076 32512
rect 53838 21040 53894 21049
rect 53838 20975 53840 20984
rect 53892 20975 53894 20984
rect 53840 20946 53892 20952
rect 53932 20936 53984 20942
rect 53932 20878 53984 20884
rect 53840 20800 53892 20806
rect 53840 20742 53892 20748
rect 53852 20058 53880 20742
rect 53840 20052 53892 20058
rect 53840 19994 53892 20000
rect 53840 17672 53892 17678
rect 53840 17614 53892 17620
rect 53852 16250 53880 17614
rect 53944 17338 53972 20878
rect 53932 17332 53984 17338
rect 53932 17274 53984 17280
rect 53944 17134 53972 17274
rect 53932 17128 53984 17134
rect 53932 17070 53984 17076
rect 53840 16244 53892 16250
rect 53840 16186 53892 16192
rect 53840 16108 53892 16114
rect 53840 16050 53892 16056
rect 53852 15910 53880 16050
rect 53840 15904 53892 15910
rect 53840 15846 53892 15852
rect 53760 4542 53880 4570
rect 53748 4480 53800 4486
rect 53748 4422 53800 4428
rect 53656 4004 53708 4010
rect 53656 3946 53708 3952
rect 53760 3466 53788 4422
rect 53852 3670 53880 4542
rect 53840 3664 53892 3670
rect 53840 3606 53892 3612
rect 53748 3460 53800 3466
rect 53748 3402 53800 3408
rect 53472 3392 53524 3398
rect 53472 3334 53524 3340
rect 53484 2582 53512 3334
rect 54036 3194 54064 32506
rect 54208 20800 54260 20806
rect 54208 20742 54260 20748
rect 54220 20466 54248 20742
rect 54208 20460 54260 20466
rect 54208 20402 54260 20408
rect 54300 19848 54352 19854
rect 54300 19790 54352 19796
rect 54312 18902 54340 19790
rect 54300 18896 54352 18902
rect 54300 18838 54352 18844
rect 54116 17196 54168 17202
rect 54116 17138 54168 17144
rect 54128 16250 54156 17138
rect 54300 16992 54352 16998
rect 54300 16934 54352 16940
rect 54312 16590 54340 16934
rect 54300 16584 54352 16590
rect 54300 16526 54352 16532
rect 54116 16244 54168 16250
rect 54116 16186 54168 16192
rect 54404 12442 54432 35866
rect 54496 20874 54524 37198
rect 54680 34542 54708 40462
rect 55680 35216 55732 35222
rect 55680 35158 55732 35164
rect 54944 35080 54996 35086
rect 54944 35022 54996 35028
rect 54668 34536 54720 34542
rect 54668 34478 54720 34484
rect 54760 32768 54812 32774
rect 54760 32710 54812 32716
rect 54668 28552 54720 28558
rect 54668 28494 54720 28500
rect 54680 22094 54708 28494
rect 54772 24274 54800 32710
rect 54760 24268 54812 24274
rect 54760 24210 54812 24216
rect 54588 22066 54708 22094
rect 54484 20868 54536 20874
rect 54484 20810 54536 20816
rect 54496 20330 54524 20810
rect 54484 20324 54536 20330
rect 54484 20266 54536 20272
rect 54588 18442 54616 22066
rect 54956 19990 54984 35022
rect 55220 26920 55272 26926
rect 55220 26862 55272 26868
rect 55036 20460 55088 20466
rect 55036 20402 55088 20408
rect 54944 19984 54996 19990
rect 54944 19926 54996 19932
rect 54668 19712 54720 19718
rect 54668 19654 54720 19660
rect 54760 19712 54812 19718
rect 54760 19654 54812 19660
rect 54680 19417 54708 19654
rect 54666 19408 54722 19417
rect 54772 19378 54800 19654
rect 55048 19514 55076 20402
rect 55128 20052 55180 20058
rect 55128 19994 55180 20000
rect 55140 19718 55168 19994
rect 55128 19712 55180 19718
rect 55128 19654 55180 19660
rect 55036 19508 55088 19514
rect 55036 19450 55088 19456
rect 54666 19343 54722 19352
rect 54760 19372 54812 19378
rect 54680 19258 54708 19343
rect 54760 19314 54812 19320
rect 54680 19230 54800 19258
rect 54496 18414 54616 18442
rect 54496 17882 54524 18414
rect 54772 18290 54800 19230
rect 54576 18284 54628 18290
rect 54576 18226 54628 18232
rect 54760 18284 54812 18290
rect 54760 18226 54812 18232
rect 54944 18284 54996 18290
rect 54944 18226 54996 18232
rect 54484 17876 54536 17882
rect 54484 17818 54536 17824
rect 54588 17270 54616 18226
rect 54772 17746 54800 18226
rect 54760 17740 54812 17746
rect 54760 17682 54812 17688
rect 54576 17264 54628 17270
rect 54576 17206 54628 17212
rect 54956 16114 54984 18226
rect 55140 17202 55168 19654
rect 55128 17196 55180 17202
rect 55128 17138 55180 17144
rect 54944 16108 54996 16114
rect 54944 16050 54996 16056
rect 55140 15910 55168 17138
rect 55128 15904 55180 15910
rect 55128 15846 55180 15852
rect 54392 12436 54444 12442
rect 54392 12378 54444 12384
rect 54208 11212 54260 11218
rect 54208 11154 54260 11160
rect 54220 3738 54248 11154
rect 54852 8288 54904 8294
rect 54852 8230 54904 8236
rect 54864 7478 54892 8230
rect 54852 7472 54904 7478
rect 54852 7414 54904 7420
rect 54484 4140 54536 4146
rect 54484 4082 54536 4088
rect 54208 3732 54260 3738
rect 54208 3674 54260 3680
rect 54024 3188 54076 3194
rect 54024 3130 54076 3136
rect 53932 3052 53984 3058
rect 53932 2994 53984 3000
rect 54208 3052 54260 3058
rect 54208 2994 54260 3000
rect 53472 2576 53524 2582
rect 53472 2518 53524 2524
rect 53840 2440 53892 2446
rect 53840 2382 53892 2388
rect 53852 898 53880 2382
rect 53668 870 53880 898
rect 53668 800 53696 870
rect 53944 800 53972 2994
rect 54220 800 54248 2994
rect 54496 800 54524 4082
rect 54760 3528 54812 3534
rect 54760 3470 54812 3476
rect 54772 800 54800 3470
rect 55232 3194 55260 26862
rect 55692 22094 55720 35158
rect 55600 22066 55720 22094
rect 55494 20904 55550 20913
rect 55494 20839 55550 20848
rect 55508 19854 55536 20839
rect 55312 19848 55364 19854
rect 55312 19790 55364 19796
rect 55496 19848 55548 19854
rect 55496 19790 55548 19796
rect 55324 17202 55352 19790
rect 55496 19236 55548 19242
rect 55496 19178 55548 19184
rect 55508 18834 55536 19178
rect 55496 18828 55548 18834
rect 55496 18770 55548 18776
rect 55312 17196 55364 17202
rect 55312 17138 55364 17144
rect 55324 16794 55352 17138
rect 55312 16788 55364 16794
rect 55312 16730 55364 16736
rect 55312 16448 55364 16454
rect 55312 16390 55364 16396
rect 55324 16182 55352 16390
rect 55312 16176 55364 16182
rect 55312 16118 55364 16124
rect 55600 12434 55628 22066
rect 55680 20936 55732 20942
rect 55680 20878 55732 20884
rect 55692 19242 55720 20878
rect 55680 19236 55732 19242
rect 55680 19178 55732 19184
rect 55680 18760 55732 18766
rect 55680 18702 55732 18708
rect 55692 18426 55720 18702
rect 55680 18420 55732 18426
rect 55680 18362 55732 18368
rect 55600 12406 55720 12434
rect 55312 9988 55364 9994
rect 55312 9930 55364 9936
rect 55324 3913 55352 9930
rect 55310 3904 55366 3913
rect 55310 3839 55366 3848
rect 55220 3188 55272 3194
rect 55220 3130 55272 3136
rect 55312 3052 55364 3058
rect 55312 2994 55364 3000
rect 55220 2440 55272 2446
rect 55220 2382 55272 2388
rect 55232 898 55260 2382
rect 55048 870 55260 898
rect 55048 800 55076 870
rect 55324 800 55352 2994
rect 55692 2514 55720 12406
rect 55784 10742 55812 61066
rect 56600 61056 56652 61062
rect 56600 60998 56652 61004
rect 56324 60512 56376 60518
rect 56324 60454 56376 60460
rect 56232 60172 56284 60178
rect 56232 60114 56284 60120
rect 56244 59770 56272 60114
rect 56232 59764 56284 59770
rect 56232 59706 56284 59712
rect 56336 59566 56364 60454
rect 56324 59560 56376 59566
rect 56324 59502 56376 59508
rect 56508 56976 56560 56982
rect 56508 56918 56560 56924
rect 55864 56772 55916 56778
rect 55864 56714 55916 56720
rect 55876 24206 55904 56714
rect 56520 56506 56548 56918
rect 56508 56500 56560 56506
rect 56508 56442 56560 56448
rect 56612 50386 56640 60998
rect 56704 60654 56732 61202
rect 56784 60784 56836 60790
rect 56784 60726 56836 60732
rect 56692 60648 56744 60654
rect 56692 60590 56744 60596
rect 56796 60110 56824 60726
rect 56888 60722 56916 63294
rect 57518 63200 57574 64000
rect 58254 63322 58310 64000
rect 58990 63322 59046 64000
rect 57992 63294 58310 63322
rect 57532 61198 57560 63200
rect 57520 61192 57572 61198
rect 57520 61134 57572 61140
rect 56876 60716 56928 60722
rect 56876 60658 56928 60664
rect 57060 60512 57112 60518
rect 57060 60454 57112 60460
rect 56784 60104 56836 60110
rect 56784 60046 56836 60052
rect 56692 60036 56744 60042
rect 56692 59978 56744 59984
rect 56600 50380 56652 50386
rect 56600 50322 56652 50328
rect 55956 48272 56008 48278
rect 55956 48214 56008 48220
rect 55864 24200 55916 24206
rect 55864 24142 55916 24148
rect 55864 20256 55916 20262
rect 55864 20198 55916 20204
rect 55876 19802 55904 20198
rect 55968 19938 55996 48214
rect 56048 40384 56100 40390
rect 56048 40326 56100 40332
rect 56060 29646 56088 40326
rect 56704 37194 56732 59978
rect 57072 45558 57100 60454
rect 57992 60110 58020 63294
rect 58254 63200 58310 63294
rect 58728 63294 59046 63322
rect 58348 61124 58400 61130
rect 58348 61066 58400 61072
rect 58072 60716 58124 60722
rect 58072 60658 58124 60664
rect 57980 60104 58032 60110
rect 57980 60046 58032 60052
rect 57336 59968 57388 59974
rect 58084 59945 58112 60658
rect 58164 60580 58216 60586
rect 58164 60522 58216 60528
rect 57336 59910 57388 59916
rect 58070 59936 58126 59945
rect 57152 59492 57204 59498
rect 57152 59434 57204 59440
rect 57164 59022 57192 59434
rect 57152 59016 57204 59022
rect 57152 58958 57204 58964
rect 57060 45552 57112 45558
rect 57060 45494 57112 45500
rect 56968 44872 57020 44878
rect 56968 44814 57020 44820
rect 56692 37188 56744 37194
rect 56692 37130 56744 37136
rect 56048 29640 56100 29646
rect 56048 29582 56100 29588
rect 56324 26376 56376 26382
rect 56324 26318 56376 26324
rect 56048 20936 56100 20942
rect 56048 20878 56100 20884
rect 56060 20058 56088 20878
rect 56336 20602 56364 26318
rect 56980 26234 57008 44814
rect 57348 36854 57376 59910
rect 58070 59871 58126 59880
rect 58176 59770 58204 60522
rect 58256 60512 58308 60518
rect 58256 60454 58308 60460
rect 58268 60314 58296 60454
rect 58256 60308 58308 60314
rect 58256 60250 58308 60256
rect 58164 59764 58216 59770
rect 58164 59706 58216 59712
rect 58072 59628 58124 59634
rect 58072 59570 58124 59576
rect 58084 59401 58112 59570
rect 58070 59392 58126 59401
rect 58070 59327 58126 59336
rect 58360 59158 58388 61066
rect 58728 59498 58756 63294
rect 58990 63200 59046 63294
rect 58806 62656 58862 62665
rect 58806 62591 58862 62600
rect 58820 59702 58848 62591
rect 58898 62112 58954 62121
rect 58898 62047 58954 62056
rect 58912 60858 58940 62047
rect 58990 61568 59046 61577
rect 58990 61503 59046 61512
rect 59004 61266 59032 61503
rect 58992 61260 59044 61266
rect 58992 61202 59044 61208
rect 58990 61024 59046 61033
rect 58990 60959 59046 60968
rect 58900 60852 58952 60858
rect 58900 60794 58952 60800
rect 59004 60790 59032 60959
rect 58992 60784 59044 60790
rect 58992 60726 59044 60732
rect 58990 60480 59046 60489
rect 58990 60415 59046 60424
rect 59004 60178 59032 60415
rect 58992 60172 59044 60178
rect 58992 60114 59044 60120
rect 59544 60036 59596 60042
rect 59544 59978 59596 59984
rect 58808 59696 58860 59702
rect 58808 59638 58860 59644
rect 58716 59492 58768 59498
rect 58716 59434 58768 59440
rect 58348 59152 58400 59158
rect 58348 59094 58400 59100
rect 58992 59016 59044 59022
rect 58992 58958 59044 58964
rect 58900 58948 58952 58954
rect 58900 58890 58952 58896
rect 58162 58848 58218 58857
rect 58162 58783 58218 58792
rect 58176 58614 58204 58783
rect 58164 58608 58216 58614
rect 58164 58550 58216 58556
rect 58256 58336 58308 58342
rect 58256 58278 58308 58284
rect 58268 57934 58296 58278
rect 58256 57928 58308 57934
rect 58256 57870 58308 57876
rect 57980 57860 58032 57866
rect 57980 57802 58032 57808
rect 57992 57769 58020 57802
rect 58072 57792 58124 57798
rect 57978 57760 58034 57769
rect 58072 57734 58124 57740
rect 57978 57695 58034 57704
rect 57520 50312 57572 50318
rect 57520 50254 57572 50260
rect 57336 36848 57388 36854
rect 57336 36790 57388 36796
rect 57428 32904 57480 32910
rect 57428 32846 57480 32852
rect 57244 29640 57296 29646
rect 57244 29582 57296 29588
rect 56888 26206 57008 26234
rect 56324 20596 56376 20602
rect 56324 20538 56376 20544
rect 56048 20052 56100 20058
rect 56048 19994 56100 20000
rect 55968 19910 56088 19938
rect 56336 19922 56364 20538
rect 55956 19848 56008 19854
rect 55876 19796 55956 19802
rect 55876 19790 56008 19796
rect 55876 19774 55996 19790
rect 55876 18222 55904 19774
rect 55864 18216 55916 18222
rect 55864 18158 55916 18164
rect 55876 17746 55904 18158
rect 55864 17740 55916 17746
rect 55864 17682 55916 17688
rect 55956 17332 56008 17338
rect 55956 17274 56008 17280
rect 55968 17134 55996 17274
rect 55956 17128 56008 17134
rect 55956 17070 56008 17076
rect 56060 11082 56088 19910
rect 56324 19916 56376 19922
rect 56324 19858 56376 19864
rect 56140 18624 56192 18630
rect 56140 18566 56192 18572
rect 56152 18358 56180 18566
rect 56140 18352 56192 18358
rect 56140 18294 56192 18300
rect 56324 17604 56376 17610
rect 56324 17546 56376 17552
rect 56336 17338 56364 17546
rect 56324 17332 56376 17338
rect 56324 17274 56376 17280
rect 56232 17196 56284 17202
rect 56232 17138 56284 17144
rect 56244 16454 56272 17138
rect 56600 16788 56652 16794
rect 56600 16730 56652 16736
rect 56232 16448 56284 16454
rect 56232 16390 56284 16396
rect 56612 12889 56640 16730
rect 56784 16516 56836 16522
rect 56784 16458 56836 16464
rect 56692 14068 56744 14074
rect 56692 14010 56744 14016
rect 56598 12880 56654 12889
rect 56140 12844 56192 12850
rect 56598 12815 56654 12824
rect 56140 12786 56192 12792
rect 56152 11150 56180 12786
rect 56416 11892 56468 11898
rect 56416 11834 56468 11840
rect 56428 11150 56456 11834
rect 56140 11144 56192 11150
rect 56140 11086 56192 11092
rect 56416 11144 56468 11150
rect 56416 11086 56468 11092
rect 56048 11076 56100 11082
rect 56048 11018 56100 11024
rect 55772 10736 55824 10742
rect 55772 10678 55824 10684
rect 56152 8974 56180 11086
rect 56324 9376 56376 9382
rect 56324 9318 56376 9324
rect 56336 8974 56364 9318
rect 56140 8968 56192 8974
rect 56140 8910 56192 8916
rect 56324 8968 56376 8974
rect 56324 8910 56376 8916
rect 56152 7818 56180 8910
rect 56416 8356 56468 8362
rect 56416 8298 56468 8304
rect 55772 7812 55824 7818
rect 55772 7754 55824 7760
rect 56140 7812 56192 7818
rect 56140 7754 56192 7760
rect 55784 7478 55812 7754
rect 56152 7478 56180 7754
rect 55772 7472 55824 7478
rect 55772 7414 55824 7420
rect 56140 7472 56192 7478
rect 56140 7414 56192 7420
rect 56428 6186 56456 8298
rect 56704 7410 56732 14010
rect 56796 10674 56824 16458
rect 56888 14278 56916 26206
rect 57060 22092 57112 22098
rect 57060 22034 57112 22040
rect 56968 20800 57020 20806
rect 56968 20742 57020 20748
rect 56980 19854 57008 20742
rect 56968 19848 57020 19854
rect 56968 19790 57020 19796
rect 57072 19718 57100 22034
rect 57152 22024 57204 22030
rect 57152 21966 57204 21972
rect 57060 19712 57112 19718
rect 57060 19654 57112 19660
rect 57164 17882 57192 21966
rect 57256 18426 57284 29582
rect 57440 22098 57468 32846
rect 57428 22092 57480 22098
rect 57428 22034 57480 22040
rect 57532 21978 57560 50254
rect 57980 49156 58032 49162
rect 57980 49098 58032 49104
rect 57992 49065 58020 49098
rect 57978 49056 58034 49065
rect 57978 48991 58034 49000
rect 58084 48278 58112 57734
rect 58346 56128 58402 56137
rect 58346 56063 58402 56072
rect 58360 55962 58388 56063
rect 58348 55956 58400 55962
rect 58348 55898 58400 55904
rect 58348 54664 58400 54670
rect 58348 54606 58400 54612
rect 58360 54505 58388 54606
rect 58346 54496 58402 54505
rect 58346 54431 58402 54440
rect 58348 52896 58400 52902
rect 58346 52864 58348 52873
rect 58400 52864 58402 52873
rect 58346 52799 58402 52808
rect 58348 51400 58400 51406
rect 58348 51342 58400 51348
rect 58360 51241 58388 51342
rect 58346 51232 58402 51241
rect 58346 51167 58402 51176
rect 58072 48272 58124 48278
rect 58072 48214 58124 48220
rect 57796 48136 57848 48142
rect 57796 48078 57848 48084
rect 57704 45960 57756 45966
rect 57704 45902 57756 45908
rect 57716 22094 57744 45902
rect 57348 21950 57560 21978
rect 57624 22066 57744 22094
rect 57244 18420 57296 18426
rect 57244 18362 57296 18368
rect 57152 17876 57204 17882
rect 57152 17818 57204 17824
rect 57164 16998 57192 17818
rect 57152 16992 57204 16998
rect 57152 16934 57204 16940
rect 56876 14272 56928 14278
rect 56876 14214 56928 14220
rect 57348 13462 57376 21950
rect 57624 21706 57652 22066
rect 57532 21678 57652 21706
rect 57532 13870 57560 21678
rect 57704 21480 57756 21486
rect 57704 21422 57756 21428
rect 57716 20534 57744 21422
rect 57704 20528 57756 20534
rect 57704 20470 57756 20476
rect 57808 14006 57836 48078
rect 58164 48068 58216 48074
rect 58164 48010 58216 48016
rect 58176 47977 58204 48010
rect 58162 47968 58218 47977
rect 58162 47903 58218 47912
rect 58072 47660 58124 47666
rect 58072 47602 58124 47608
rect 58084 47433 58112 47602
rect 58808 47456 58860 47462
rect 58070 47424 58126 47433
rect 58808 47398 58860 47404
rect 58070 47359 58126 47368
rect 58162 46336 58218 46345
rect 58162 46271 58218 46280
rect 58176 46034 58204 46271
rect 58164 46028 58216 46034
rect 58164 45970 58216 45976
rect 58440 45280 58492 45286
rect 58440 45222 58492 45228
rect 58348 44736 58400 44742
rect 58348 44678 58400 44684
rect 58164 43716 58216 43722
rect 58164 43658 58216 43664
rect 58176 43081 58204 43658
rect 58162 43072 58218 43081
rect 58162 43007 58218 43016
rect 57980 42628 58032 42634
rect 57980 42570 58032 42576
rect 57992 41993 58020 42570
rect 57978 41984 58034 41993
rect 57978 41919 58034 41928
rect 58360 40186 58388 44678
rect 58348 40180 58400 40186
rect 58348 40122 58400 40128
rect 57980 39364 58032 39370
rect 57980 39306 58032 39312
rect 58348 39364 58400 39370
rect 58348 39306 58400 39312
rect 57992 38729 58020 39306
rect 57978 38720 58034 38729
rect 57978 38655 58034 38664
rect 58164 38276 58216 38282
rect 58164 38218 58216 38224
rect 58176 38185 58204 38218
rect 58162 38176 58218 38185
rect 58162 38111 58218 38120
rect 58072 37868 58124 37874
rect 58072 37810 58124 37816
rect 58084 37641 58112 37810
rect 58070 37632 58126 37641
rect 58070 37567 58126 37576
rect 58164 37188 58216 37194
rect 58164 37130 58216 37136
rect 58176 36553 58204 37130
rect 58162 36544 58218 36553
rect 58162 36479 58218 36488
rect 57980 36100 58032 36106
rect 57980 36042 58032 36048
rect 57992 36009 58020 36042
rect 57978 36000 58034 36009
rect 57978 35935 58034 35944
rect 58164 35012 58216 35018
rect 58164 34954 58216 34960
rect 58176 34921 58204 34954
rect 58162 34912 58218 34921
rect 58162 34847 58218 34856
rect 58072 31340 58124 31346
rect 58072 31282 58124 31288
rect 58084 31113 58112 31282
rect 58070 31104 58126 31113
rect 58070 31039 58126 31048
rect 58162 30016 58218 30025
rect 58162 29951 58218 29960
rect 58176 29714 58204 29951
rect 58164 29708 58216 29714
rect 58164 29650 58216 29656
rect 58164 28484 58216 28490
rect 58164 28426 58216 28432
rect 58176 28393 58204 28426
rect 58162 28384 58218 28393
rect 58162 28319 58218 28328
rect 58162 26752 58218 26761
rect 58162 26687 58218 26696
rect 58176 26450 58204 26687
rect 58164 26444 58216 26450
rect 58164 26386 58216 26392
rect 58070 26208 58126 26217
rect 58070 26143 58126 26152
rect 58084 25906 58112 26143
rect 58072 25900 58124 25906
rect 58072 25842 58124 25848
rect 57980 25696 58032 25702
rect 57980 25638 58032 25644
rect 57888 23112 57940 23118
rect 57888 23054 57940 23060
rect 57900 21486 57928 23054
rect 57888 21480 57940 21486
rect 57888 21422 57940 21428
rect 57888 21344 57940 21350
rect 57888 21286 57940 21292
rect 57900 20942 57928 21286
rect 57992 21146 58020 25638
rect 58164 25220 58216 25226
rect 58164 25162 58216 25168
rect 58176 25129 58204 25162
rect 58162 25120 58218 25129
rect 58162 25055 58218 25064
rect 58072 24812 58124 24818
rect 58072 24754 58124 24760
rect 58084 24585 58112 24754
rect 58070 24576 58126 24585
rect 58070 24511 58126 24520
rect 58162 22944 58218 22953
rect 58162 22879 58218 22888
rect 58176 22710 58204 22879
rect 58164 22704 58216 22710
rect 58164 22646 58216 22652
rect 58164 21956 58216 21962
rect 58164 21898 58216 21904
rect 58176 21865 58204 21898
rect 58162 21856 58218 21865
rect 58162 21791 58218 21800
rect 58072 21548 58124 21554
rect 58072 21490 58124 21496
rect 58084 21321 58112 21490
rect 58256 21344 58308 21350
rect 58070 21312 58126 21321
rect 58256 21286 58308 21292
rect 58070 21247 58126 21256
rect 57980 21140 58032 21146
rect 57980 21082 58032 21088
rect 57888 20936 57940 20942
rect 57888 20878 57940 20884
rect 58072 18624 58124 18630
rect 58072 18566 58124 18572
rect 58084 17270 58112 18566
rect 58268 17678 58296 21286
rect 58256 17672 58308 17678
rect 58256 17614 58308 17620
rect 58072 17264 58124 17270
rect 58072 17206 58124 17212
rect 58072 16448 58124 16454
rect 58072 16390 58124 16396
rect 58084 15609 58112 16390
rect 58070 15600 58126 15609
rect 58070 15535 58126 15544
rect 58164 15428 58216 15434
rect 58164 15370 58216 15376
rect 58176 15337 58204 15370
rect 58162 15328 58218 15337
rect 58162 15263 58218 15272
rect 58070 15056 58126 15065
rect 58070 14991 58126 15000
rect 57978 14784 58034 14793
rect 57978 14719 58034 14728
rect 57992 14414 58020 14719
rect 58084 14618 58112 14991
rect 58072 14612 58124 14618
rect 58072 14554 58124 14560
rect 57980 14408 58032 14414
rect 57980 14350 58032 14356
rect 57796 14000 57848 14006
rect 57796 13942 57848 13948
rect 57520 13864 57572 13870
rect 57520 13806 57572 13812
rect 58162 13696 58218 13705
rect 58162 13631 58218 13640
rect 57336 13456 57388 13462
rect 57336 13398 57388 13404
rect 58176 13394 58204 13631
rect 58164 13388 58216 13394
rect 58164 13330 58216 13336
rect 57152 13184 57204 13190
rect 57152 13126 57204 13132
rect 56876 11144 56928 11150
rect 56876 11086 56928 11092
rect 56784 10668 56836 10674
rect 56784 10610 56836 10616
rect 56796 9586 56824 10610
rect 56888 9926 56916 11086
rect 56968 11076 57020 11082
rect 56968 11018 57020 11024
rect 56980 10810 57008 11018
rect 56968 10804 57020 10810
rect 56968 10746 57020 10752
rect 56876 9920 56928 9926
rect 56876 9862 56928 9868
rect 56784 9580 56836 9586
rect 56784 9522 56836 9528
rect 56796 8090 56824 9522
rect 56888 9042 56916 9862
rect 56876 9036 56928 9042
rect 56876 8978 56928 8984
rect 56784 8084 56836 8090
rect 56784 8026 56836 8032
rect 56796 7410 56824 8026
rect 56888 7954 56916 8978
rect 56876 7948 56928 7954
rect 56876 7890 56928 7896
rect 56692 7404 56744 7410
rect 56692 7346 56744 7352
rect 56784 7404 56836 7410
rect 56784 7346 56836 7352
rect 56416 6180 56468 6186
rect 56416 6122 56468 6128
rect 56704 4826 56732 7346
rect 56888 6866 56916 7890
rect 56968 7200 57020 7206
rect 56968 7142 57020 7148
rect 56876 6860 56928 6866
rect 56876 6802 56928 6808
rect 56692 4820 56744 4826
rect 56692 4762 56744 4768
rect 56888 3602 56916 6802
rect 56980 6798 57008 7142
rect 56968 6792 57020 6798
rect 56968 6734 57020 6740
rect 57164 5574 57192 13126
rect 57888 12232 57940 12238
rect 57888 12174 57940 12180
rect 57244 11552 57296 11558
rect 57244 11494 57296 11500
rect 57256 11354 57284 11494
rect 57244 11348 57296 11354
rect 57244 11290 57296 11296
rect 57900 11286 57928 12174
rect 58164 12164 58216 12170
rect 58164 12106 58216 12112
rect 58176 12073 58204 12106
rect 58162 12064 58218 12073
rect 58162 11999 58218 12008
rect 57888 11280 57940 11286
rect 57888 11222 57940 11228
rect 57900 10674 57928 11222
rect 57888 10668 57940 10674
rect 57888 10610 57940 10616
rect 58162 10432 58218 10441
rect 58162 10367 58218 10376
rect 58176 10130 58204 10367
rect 58164 10124 58216 10130
rect 58164 10066 58216 10072
rect 57244 9580 57296 9586
rect 57244 9522 57296 9528
rect 57256 8838 57284 9522
rect 58360 9178 58388 39306
rect 58452 15026 58480 45222
rect 58716 44804 58768 44810
rect 58716 44746 58768 44752
rect 58728 44169 58756 44746
rect 58714 44160 58770 44169
rect 58714 44095 58770 44104
rect 58532 42628 58584 42634
rect 58532 42570 58584 42576
rect 58544 15706 58572 42570
rect 58716 41540 58768 41546
rect 58716 41482 58768 41488
rect 58624 41472 58676 41478
rect 58624 41414 58676 41420
rect 58636 19174 58664 41414
rect 58728 40905 58756 41482
rect 58714 40896 58770 40905
rect 58714 40831 58770 40840
rect 58716 40384 58768 40390
rect 58714 40352 58716 40361
rect 58768 40352 58770 40361
rect 58714 40287 58770 40296
rect 58716 40180 58768 40186
rect 58716 40122 58768 40128
rect 58624 19168 58676 19174
rect 58624 19110 58676 19116
rect 58728 18426 58756 40122
rect 58716 18420 58768 18426
rect 58716 18362 58768 18368
rect 58820 18306 58848 47398
rect 58636 18278 58848 18306
rect 58532 15700 58584 15706
rect 58532 15642 58584 15648
rect 58636 15366 58664 18278
rect 58716 18148 58768 18154
rect 58716 18090 58768 18096
rect 58624 15360 58676 15366
rect 58624 15302 58676 15308
rect 58440 15020 58492 15026
rect 58440 14962 58492 14968
rect 58348 9172 58400 9178
rect 58348 9114 58400 9120
rect 57244 8832 57296 8838
rect 57244 8774 57296 8780
rect 57256 8498 57284 8774
rect 57244 8492 57296 8498
rect 57244 8434 57296 8440
rect 58728 8294 58756 18090
rect 58806 18048 58862 18057
rect 58806 17983 58862 17992
rect 58820 16590 58848 17983
rect 58808 16584 58860 16590
rect 58808 16526 58860 16532
rect 58912 8634 58940 58890
rect 59004 58313 59032 58958
rect 58990 58304 59046 58313
rect 58990 58239 59046 58248
rect 58990 57216 59046 57225
rect 58990 57151 59046 57160
rect 59004 56846 59032 57151
rect 58992 56840 59044 56846
rect 58992 56782 59044 56788
rect 58990 56672 59046 56681
rect 58990 56607 59046 56616
rect 59004 56438 59032 56607
rect 58992 56432 59044 56438
rect 58992 56374 59044 56380
rect 58992 50244 59044 50250
rect 58992 50186 59044 50192
rect 59004 49609 59032 50186
rect 58990 49600 59046 49609
rect 58990 49535 59046 49544
rect 59452 49156 59504 49162
rect 59452 49098 59504 49104
rect 58990 45792 59046 45801
rect 58990 45727 59046 45736
rect 59004 45490 59032 45727
rect 58992 45484 59044 45490
rect 58992 45426 59044 45432
rect 58992 44872 59044 44878
rect 58992 44814 59044 44820
rect 59004 44713 59032 44814
rect 58990 44704 59046 44713
rect 58990 44639 59046 44648
rect 58992 42696 59044 42702
rect 58992 42638 59044 42644
rect 59004 42537 59032 42638
rect 58990 42528 59046 42537
rect 58990 42463 59046 42472
rect 58992 41608 59044 41614
rect 58992 41550 59044 41556
rect 59004 41449 59032 41550
rect 58990 41440 59046 41449
rect 58990 41375 59046 41384
rect 58992 40452 59044 40458
rect 58992 40394 59044 40400
rect 59004 39817 59032 40394
rect 58990 39808 59046 39817
rect 58990 39743 59046 39752
rect 58992 39432 59044 39438
rect 58992 39374 59044 39380
rect 59004 39273 59032 39374
rect 58990 39264 59046 39273
rect 58990 39199 59046 39208
rect 59176 37664 59228 37670
rect 59176 37606 59228 37612
rect 59188 35894 59216 37606
rect 59268 36100 59320 36106
rect 59268 36042 59320 36048
rect 59096 35866 59216 35894
rect 58992 34604 59044 34610
rect 58992 34546 59044 34552
rect 59004 34377 59032 34546
rect 58990 34368 59046 34377
rect 58990 34303 59046 34312
rect 58990 33280 59046 33289
rect 58990 33215 59046 33224
rect 59004 32978 59032 33215
rect 58992 32972 59044 32978
rect 58992 32914 59044 32920
rect 58992 32836 59044 32842
rect 58992 32778 59044 32784
rect 59004 32745 59032 32778
rect 58990 32736 59046 32745
rect 58990 32671 59046 32680
rect 58992 31816 59044 31822
rect 58992 31758 59044 31764
rect 59004 31657 59032 31758
rect 58990 31648 59046 31657
rect 58990 31583 59046 31592
rect 58992 29572 59044 29578
rect 58992 29514 59044 29520
rect 59004 29481 59032 29514
rect 58990 29472 59046 29481
rect 58990 29407 59046 29416
rect 58990 27840 59046 27849
rect 58990 27775 59046 27784
rect 59004 27470 59032 27775
rect 58992 27464 59044 27470
rect 58992 27406 59044 27412
rect 58990 23488 59046 23497
rect 58990 23423 59046 23432
rect 59004 23186 59032 23423
rect 58992 23180 59044 23186
rect 58992 23122 59044 23128
rect 58992 20868 59044 20874
rect 58992 20810 59044 20816
rect 59004 20233 59032 20810
rect 58990 20224 59046 20233
rect 58990 20159 59046 20168
rect 58990 19680 59046 19689
rect 58990 19615 59046 19624
rect 59004 18766 59032 19615
rect 58992 18760 59044 18766
rect 58992 18702 59044 18708
rect 58992 18624 59044 18630
rect 58990 18592 58992 18601
rect 59044 18592 59046 18601
rect 58990 18527 59046 18536
rect 59096 17649 59124 35866
rect 59280 31090 59308 36042
rect 59360 34740 59412 34746
rect 59360 34682 59412 34688
rect 59188 31062 59308 31090
rect 59188 22778 59216 31062
rect 59372 26234 59400 34682
rect 59280 26206 59400 26234
rect 59176 22772 59228 22778
rect 59176 22714 59228 22720
rect 59280 21078 59308 26206
rect 59268 21072 59320 21078
rect 59268 21014 59320 21020
rect 59082 17640 59138 17649
rect 59082 17575 59138 17584
rect 58992 17128 59044 17134
rect 58992 17070 59044 17076
rect 59004 16969 59032 17070
rect 58990 16960 59046 16969
rect 58990 16895 59046 16904
rect 58992 16516 59044 16522
rect 58992 16458 59044 16464
rect 59004 16425 59032 16458
rect 58990 16416 59046 16425
rect 58990 16351 59046 16360
rect 58992 13252 59044 13258
rect 58992 13194 59044 13200
rect 59004 13161 59032 13194
rect 58990 13152 59046 13161
rect 58990 13087 59046 13096
rect 59464 11830 59492 49098
rect 59556 31958 59584 59978
rect 59544 31952 59596 31958
rect 59544 31894 59596 31900
rect 59452 11824 59504 11830
rect 59452 11766 59504 11772
rect 58992 11756 59044 11762
rect 58992 11698 59044 11704
rect 59004 11529 59032 11698
rect 58990 11520 59046 11529
rect 58990 11455 59046 11464
rect 58992 9988 59044 9994
rect 58992 9930 59044 9936
rect 59004 9897 59032 9930
rect 58990 9888 59046 9897
rect 58990 9823 59046 9832
rect 58990 8800 59046 8809
rect 58990 8735 59046 8744
rect 58900 8628 58952 8634
rect 58900 8570 58952 8576
rect 59004 8566 59032 8735
rect 58992 8560 59044 8566
rect 58992 8502 59044 8508
rect 58992 8424 59044 8430
rect 58992 8366 59044 8372
rect 58716 8288 58768 8294
rect 59004 8265 59032 8366
rect 58716 8230 58768 8236
rect 58990 8256 59046 8265
rect 58990 8191 59046 8200
rect 57888 7812 57940 7818
rect 57888 7754 57940 7760
rect 57900 5710 57928 7754
rect 58256 7404 58308 7410
rect 58256 7346 58308 7352
rect 58268 6662 58296 7346
rect 58898 7168 58954 7177
rect 58898 7103 58954 7112
rect 58256 6656 58308 6662
rect 58070 6624 58126 6633
rect 58256 6598 58308 6604
rect 58070 6559 58126 6568
rect 58084 6322 58112 6559
rect 58072 6316 58124 6322
rect 58072 6258 58124 6264
rect 58268 5846 58296 6598
rect 58256 5840 58308 5846
rect 58256 5782 58308 5788
rect 58912 5710 58940 7103
rect 58992 5772 59044 5778
rect 58992 5714 59044 5720
rect 57888 5704 57940 5710
rect 57888 5646 57940 5652
rect 58900 5704 58952 5710
rect 58900 5646 58952 5652
rect 57152 5568 57204 5574
rect 59004 5545 59032 5714
rect 57152 5510 57204 5516
rect 58990 5536 59046 5545
rect 58990 5471 59046 5480
rect 58072 5228 58124 5234
rect 58072 5170 58124 5176
rect 58084 5001 58112 5170
rect 58070 4992 58126 5001
rect 58070 4927 58126 4936
rect 58808 4616 58860 4622
rect 58808 4558 58860 4564
rect 57428 3936 57480 3942
rect 57428 3878 57480 3884
rect 56876 3596 56928 3602
rect 56876 3538 56928 3544
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 55680 2508 55732 2514
rect 55680 2450 55732 2456
rect 57256 2446 57284 3334
rect 57440 3194 57468 3878
rect 58162 3360 58218 3369
rect 58162 3295 58218 3304
rect 57428 3188 57480 3194
rect 57428 3130 57480 3136
rect 58176 3126 58204 3295
rect 58164 3120 58216 3126
rect 58164 3062 58216 3068
rect 58256 3052 58308 3058
rect 58256 2994 58308 3000
rect 58268 2650 58296 2994
rect 58256 2644 58308 2650
rect 58256 2586 58308 2592
rect 57244 2440 57296 2446
rect 57244 2382 57296 2388
rect 58820 1737 58848 4558
rect 58992 4208 59044 4214
rect 58992 4150 59044 4156
rect 59004 3913 59032 4150
rect 58990 3904 59046 3913
rect 58990 3839 59046 3848
rect 58990 2816 59046 2825
rect 58990 2751 59046 2760
rect 59004 2446 59032 2751
rect 58992 2440 59044 2446
rect 58992 2382 59044 2388
rect 58900 2372 58952 2378
rect 58900 2314 58952 2320
rect 58912 2281 58940 2314
rect 58898 2272 58954 2281
rect 58898 2207 58954 2216
rect 58806 1728 58862 1737
rect 58806 1663 58862 1672
rect 56508 1352 56560 1358
rect 56508 1294 56560 1300
rect 56520 1193 56548 1294
rect 56506 1184 56562 1193
rect 56506 1119 56562 1128
rect 38936 400 38988 406
rect 38936 342 38988 348
rect 38844 128 38896 134
rect 38844 70 38896 76
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 53930 0 53986 800
rect 54206 0 54262 800
rect 54482 0 54538 800
rect 54758 0 54814 800
rect 55034 0 55090 800
rect 55310 0 55366 800
<< via2 >>
rect 938 61784 994 61840
rect 1030 61124 1086 61160
rect 1030 61104 1032 61124
rect 1032 61104 1084 61124
rect 1084 61104 1086 61124
rect 938 60424 994 60480
rect 938 59744 994 59800
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 938 59064 994 59120
rect 938 58384 994 58440
rect 938 57704 994 57760
rect 938 57024 994 57080
rect 938 56344 994 56400
rect 938 55684 994 55720
rect 938 55664 940 55684
rect 940 55664 992 55684
rect 992 55664 994 55684
rect 938 54984 994 55040
rect 938 54304 994 54360
rect 938 53624 994 53680
rect 938 52944 994 53000
rect 2042 52536 2098 52592
rect 938 52264 994 52320
rect 938 51584 994 51640
rect 938 50904 994 50960
rect 938 50244 994 50280
rect 938 50224 940 50244
rect 940 50224 992 50244
rect 992 50224 994 50244
rect 938 49544 994 49600
rect 938 48864 994 48920
rect 938 48184 994 48240
rect 938 47504 994 47560
rect 938 46824 994 46880
rect 938 46144 994 46200
rect 938 45464 994 45520
rect 938 44820 940 44840
rect 940 44820 992 44840
rect 992 44820 994 44840
rect 938 44784 994 44820
rect 938 44104 994 44160
rect 938 43424 994 43480
rect 938 42744 994 42800
rect 938 42064 994 42120
rect 938 41384 994 41440
rect 938 40704 994 40760
rect 938 40024 994 40080
rect 1030 39344 1086 39400
rect 938 38664 994 38720
rect 1030 37984 1086 38040
rect 938 37304 994 37360
rect 938 36624 994 36680
rect 938 35944 994 36000
rect 1858 44820 1860 44840
rect 1860 44820 1912 44840
rect 1912 44820 1914 44840
rect 1858 44784 1914 44820
rect 938 35264 994 35320
rect 938 34584 994 34640
rect 938 33940 940 33960
rect 940 33940 992 33960
rect 992 33940 994 33960
rect 938 33904 994 33940
rect 938 33224 994 33280
rect 938 32544 994 32600
rect 938 31864 994 31920
rect 938 31184 994 31240
rect 938 30504 994 30560
rect 938 29824 994 29880
rect 938 29144 994 29200
rect 938 28464 994 28520
rect 938 27784 994 27840
rect 938 27104 994 27160
rect 938 26424 994 26480
rect 938 25780 940 25800
rect 940 25780 992 25800
rect 992 25780 994 25800
rect 938 25744 994 25780
rect 938 25064 994 25120
rect 938 24384 994 24440
rect 938 23704 994 23760
rect 938 23024 994 23080
rect 938 22344 994 22400
rect 938 21664 994 21720
rect 938 20984 994 21040
rect 938 20340 940 20360
rect 940 20340 992 20360
rect 992 20340 994 20360
rect 938 20304 994 20340
rect 938 19624 994 19680
rect 938 18944 994 19000
rect 938 18264 994 18320
rect 938 17584 994 17640
rect 938 16904 994 16960
rect 938 16224 994 16280
rect 938 15544 994 15600
rect 938 14900 940 14920
rect 940 14900 992 14920
rect 992 14900 994 14920
rect 938 14864 994 14900
rect 1582 14456 1638 14512
rect 938 14184 994 14240
rect 938 13504 994 13560
rect 1582 13368 1638 13424
rect 938 12824 994 12880
rect 938 12144 994 12200
rect 938 11464 994 11520
rect 938 10784 994 10840
rect 938 10124 994 10160
rect 938 10104 940 10124
rect 940 10104 992 10124
rect 992 10104 994 10124
rect 938 9460 940 9480
rect 940 9460 992 9480
rect 992 9460 994 9480
rect 938 9424 994 9460
rect 938 8744 994 8800
rect 938 8064 994 8120
rect 938 7384 994 7440
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 2410 9424 2466 9480
rect 2502 8880 2558 8936
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 6182 35128 6238 35184
rect 7746 44240 7802 44296
rect 5538 17720 5594 17776
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 7010 13232 7066 13288
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4066 12144 4122 12200
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 938 6704 994 6760
rect 1858 6704 1914 6760
rect 938 6024 994 6080
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 938 5344 994 5400
rect 5262 4936 5318 4992
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 938 4664 994 4720
rect 938 4020 940 4040
rect 940 4020 992 4040
rect 992 4020 994 4040
rect 938 3984 994 4020
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 5722 3984 5778 4040
rect 938 3304 994 3360
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 938 2624 994 2680
rect 938 1944 994 2000
rect 5814 3032 5870 3088
rect 9678 20440 9734 20496
rect 11886 18944 11942 19000
rect 12622 18808 12678 18864
rect 11242 17176 11298 17232
rect 5998 2896 6054 2952
rect 6918 3168 6974 3224
rect 7930 7928 7986 7984
rect 7654 2760 7710 2816
rect 9586 10668 9642 10704
rect 9586 10648 9588 10668
rect 9588 10648 9640 10668
rect 9640 10648 9642 10668
rect 9770 4684 9826 4720
rect 10874 10376 10930 10432
rect 9770 4664 9772 4684
rect 9772 4664 9824 4684
rect 9824 4664 9826 4684
rect 8942 4020 8944 4040
rect 8944 4020 8996 4040
rect 8996 4020 8998 4040
rect 8942 3984 8998 4020
rect 9310 3032 9366 3088
rect 9494 3052 9550 3088
rect 9494 3032 9496 3052
rect 9496 3032 9548 3052
rect 9548 3032 9550 3052
rect 13450 16652 13506 16688
rect 13450 16632 13452 16652
rect 13452 16632 13504 16652
rect 13504 16632 13506 16652
rect 13358 16532 13360 16552
rect 13360 16532 13412 16552
rect 13412 16532 13414 16552
rect 13358 16496 13414 16532
rect 10322 2760 10378 2816
rect 12898 4020 12900 4040
rect 12900 4020 12952 4040
rect 12952 4020 12954 4040
rect 12898 3984 12954 4020
rect 12622 3576 12678 3632
rect 13266 9968 13322 10024
rect 15198 47504 15254 47560
rect 17590 50224 17646 50280
rect 14462 18128 14518 18184
rect 13818 16108 13874 16144
rect 13818 16088 13820 16108
rect 13820 16088 13872 16108
rect 13872 16088 13874 16108
rect 13634 9152 13690 9208
rect 12990 3576 13046 3632
rect 15106 12688 15162 12744
rect 15198 9868 15200 9888
rect 15200 9868 15252 9888
rect 15252 9868 15254 9888
rect 15198 9832 15254 9868
rect 16486 15952 16542 16008
rect 14830 8064 14886 8120
rect 15198 7420 15200 7440
rect 15200 7420 15252 7440
rect 15252 7420 15254 7440
rect 15198 7384 15254 7420
rect 15658 11192 15714 11248
rect 15382 6316 15438 6352
rect 15382 6296 15384 6316
rect 15384 6296 15436 6316
rect 15436 6296 15438 6316
rect 14922 5208 14978 5264
rect 14830 4664 14886 4720
rect 14738 4528 14794 4584
rect 15290 4800 15346 4856
rect 15198 3712 15254 3768
rect 14830 2896 14886 2952
rect 15842 9580 15898 9616
rect 15842 9560 15844 9580
rect 15844 9560 15896 9580
rect 15896 9560 15898 9580
rect 15750 6860 15806 6896
rect 15750 6840 15752 6860
rect 15752 6840 15804 6860
rect 15804 6840 15806 6860
rect 15934 6160 15990 6216
rect 17314 19896 17370 19952
rect 17222 19352 17278 19408
rect 17222 18944 17278 19000
rect 16762 13776 16818 13832
rect 16670 12280 16726 12336
rect 16394 9832 16450 9888
rect 15842 3440 15898 3496
rect 19580 60954 19636 60956
rect 19660 60954 19716 60956
rect 19740 60954 19796 60956
rect 19820 60954 19876 60956
rect 19580 60902 19626 60954
rect 19626 60902 19636 60954
rect 19660 60902 19690 60954
rect 19690 60902 19702 60954
rect 19702 60902 19716 60954
rect 19740 60902 19754 60954
rect 19754 60902 19766 60954
rect 19766 60902 19796 60954
rect 19820 60902 19830 60954
rect 19830 60902 19876 60954
rect 19580 60900 19636 60902
rect 19660 60900 19716 60902
rect 19740 60900 19796 60902
rect 19820 60900 19876 60902
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 21822 59336 21878 59392
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 20626 37848 20682 37904
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 18142 20304 18198 20360
rect 17958 20052 18014 20088
rect 17958 20032 17960 20052
rect 17960 20032 18012 20052
rect 18012 20032 18014 20052
rect 18142 18128 18198 18184
rect 18326 16904 18382 16960
rect 17682 12688 17738 12744
rect 18142 12688 18198 12744
rect 17866 11328 17922 11384
rect 17590 11056 17646 11112
rect 17130 10512 17186 10568
rect 17222 10240 17278 10296
rect 17130 8472 17186 8528
rect 17682 10104 17738 10160
rect 17590 6840 17646 6896
rect 17774 9016 17830 9072
rect 17958 8064 18014 8120
rect 17958 4664 18014 4720
rect 18326 12688 18382 12744
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 18786 16632 18842 16688
rect 18694 13776 18750 13832
rect 18234 9288 18290 9344
rect 18510 5072 18566 5128
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19706 21292 19708 21312
rect 19708 21292 19760 21312
rect 19760 21292 19762 21312
rect 19706 21256 19762 21292
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19890 19216 19946 19272
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 20074 20984 20130 21040
rect 20810 34584 20866 34640
rect 21546 37848 21602 37904
rect 22190 60732 22192 60752
rect 22192 60732 22244 60752
rect 22244 60732 22246 60752
rect 22190 60696 22246 60732
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19522 13640 19578 13696
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19522 11600 19578 11656
rect 19430 11464 19486 11520
rect 21178 19216 21234 19272
rect 20626 14728 20682 14784
rect 20166 14048 20222 14104
rect 20350 11464 20406 11520
rect 22466 38664 22522 38720
rect 23110 38820 23166 38856
rect 23110 38800 23112 38820
rect 23112 38800 23164 38820
rect 23164 38800 23166 38820
rect 23018 37712 23074 37768
rect 22282 33360 22338 33416
rect 21454 18944 21510 19000
rect 19982 10920 20038 10976
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 20166 9832 20222 9888
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19982 9696 20038 9752
rect 19338 8200 19394 8256
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 20074 9016 20130 9072
rect 20074 8744 20130 8800
rect 19338 6024 19394 6080
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 20350 10784 20406 10840
rect 20534 10784 20590 10840
rect 21178 12724 21180 12744
rect 21180 12724 21232 12744
rect 21232 12724 21234 12744
rect 21178 12688 21234 12724
rect 20994 11464 21050 11520
rect 20442 4428 20444 4448
rect 20444 4428 20496 4448
rect 20496 4428 20498 4448
rect 20442 4392 20498 4428
rect 19706 3596 19762 3632
rect 19706 3576 19708 3596
rect 19708 3576 19760 3596
rect 19760 3576 19762 3596
rect 19338 3168 19394 3224
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21362 11600 21418 11656
rect 21454 9696 21510 9752
rect 20534 3304 20590 3360
rect 20718 2896 20774 2952
rect 21638 13640 21694 13696
rect 21638 12844 21694 12880
rect 21638 12824 21640 12844
rect 21640 12824 21692 12844
rect 21692 12824 21694 12844
rect 21638 11092 21640 11112
rect 21640 11092 21692 11112
rect 21692 11092 21694 11112
rect 21638 11056 21694 11092
rect 21822 12436 21878 12472
rect 21822 12416 21824 12436
rect 21824 12416 21876 12436
rect 21876 12416 21878 12436
rect 21730 9832 21786 9888
rect 21638 4800 21694 4856
rect 22190 19760 22246 19816
rect 22006 9152 22062 9208
rect 22006 7248 22062 7304
rect 22190 12844 22246 12880
rect 22190 12824 22192 12844
rect 22192 12824 22244 12844
rect 22244 12824 22246 12844
rect 22650 29824 22706 29880
rect 22834 18672 22890 18728
rect 22834 16632 22890 16688
rect 22742 16360 22798 16416
rect 23938 55276 23994 55312
rect 23938 55256 23940 55276
rect 23940 55256 23992 55276
rect 23992 55256 23994 55276
rect 23754 27648 23810 27704
rect 23202 19760 23258 19816
rect 23202 18944 23258 19000
rect 22466 14320 22522 14376
rect 22374 14068 22430 14104
rect 22374 14048 22376 14068
rect 22376 14048 22428 14068
rect 22428 14048 22430 14068
rect 22558 11464 22614 11520
rect 22374 6976 22430 7032
rect 22190 6296 22246 6352
rect 22374 5480 22430 5536
rect 23294 13912 23350 13968
rect 23386 13640 23442 13696
rect 23018 12688 23074 12744
rect 22742 4800 22798 4856
rect 22558 4120 22614 4176
rect 22650 3984 22706 4040
rect 22650 3576 22706 3632
rect 22926 8336 22982 8392
rect 23202 11600 23258 11656
rect 23294 10376 23350 10432
rect 24122 34584 24178 34640
rect 25134 37868 25190 37904
rect 25134 37848 25136 37868
rect 25136 37848 25188 37868
rect 25188 37848 25190 37868
rect 25226 27648 25282 27704
rect 24030 20848 24086 20904
rect 23478 8900 23534 8936
rect 23478 8880 23480 8900
rect 23480 8880 23532 8900
rect 23532 8880 23534 8900
rect 23386 8628 23442 8664
rect 23386 8608 23388 8628
rect 23388 8608 23440 8628
rect 23440 8608 23442 8628
rect 23386 4936 23442 4992
rect 23662 4664 23718 4720
rect 24306 12280 24362 12336
rect 24674 19216 24730 19272
rect 24766 17856 24822 17912
rect 24766 13776 24822 13832
rect 24950 14456 25006 14512
rect 25778 20984 25834 21040
rect 25318 16904 25374 16960
rect 25410 16360 25466 16416
rect 25226 15136 25282 15192
rect 25042 13932 25098 13968
rect 25042 13912 25044 13932
rect 25044 13912 25096 13932
rect 25096 13912 25098 13932
rect 25318 14492 25320 14512
rect 25320 14492 25372 14512
rect 25372 14492 25374 14512
rect 25318 14456 25374 14492
rect 25318 14220 25320 14240
rect 25320 14220 25372 14240
rect 25372 14220 25374 14240
rect 25318 14184 25374 14220
rect 24214 8064 24270 8120
rect 23662 3440 23718 3496
rect 23662 3188 23718 3224
rect 23662 3168 23664 3188
rect 23664 3168 23716 3188
rect 23716 3168 23718 3188
rect 24858 12008 24914 12064
rect 25594 19372 25650 19408
rect 25594 19352 25596 19372
rect 25596 19352 25648 19372
rect 25648 19352 25650 19372
rect 25042 10376 25098 10432
rect 24766 7792 24822 7848
rect 25778 15020 25834 15056
rect 25778 15000 25780 15020
rect 25780 15000 25832 15020
rect 25832 15000 25834 15020
rect 26146 21256 26202 21312
rect 26790 20984 26846 21040
rect 25962 20440 26018 20496
rect 26146 20052 26202 20088
rect 26146 20032 26148 20052
rect 26148 20032 26200 20052
rect 26200 20032 26202 20052
rect 26054 16904 26110 16960
rect 25962 14492 25964 14512
rect 25964 14492 26016 14512
rect 26016 14492 26018 14512
rect 25962 14456 26018 14492
rect 25686 11600 25742 11656
rect 25594 8064 25650 8120
rect 26146 14068 26202 14104
rect 26146 14048 26148 14068
rect 26148 14048 26200 14068
rect 26200 14048 26202 14068
rect 26238 12824 26294 12880
rect 26054 10376 26110 10432
rect 26054 9696 26110 9752
rect 25870 9152 25926 9208
rect 25778 8916 25780 8936
rect 25780 8916 25832 8936
rect 25832 8916 25834 8936
rect 25778 8880 25834 8916
rect 26146 9288 26202 9344
rect 26514 12416 26570 12472
rect 26514 12044 26516 12064
rect 26516 12044 26568 12064
rect 26568 12044 26570 12064
rect 26514 12008 26570 12044
rect 26514 9696 26570 9752
rect 26330 9288 26386 9344
rect 26698 14728 26754 14784
rect 27066 17620 27068 17640
rect 27068 17620 27120 17640
rect 27120 17620 27122 17640
rect 27066 17584 27122 17620
rect 29090 59916 29092 59936
rect 29092 59916 29144 59936
rect 29144 59916 29146 59936
rect 29090 59880 29146 59916
rect 29734 59472 29790 59528
rect 27526 19780 27582 19816
rect 27526 19760 27528 19780
rect 27528 19760 27580 19780
rect 27580 19760 27582 19780
rect 26790 9288 26846 9344
rect 27158 10376 27214 10432
rect 26790 8744 26846 8800
rect 26330 8608 26386 8664
rect 25226 5208 25282 5264
rect 24122 2760 24178 2816
rect 26514 8336 26570 8392
rect 26698 8064 26754 8120
rect 25778 3984 25834 4040
rect 26698 7384 26754 7440
rect 26882 8336 26938 8392
rect 26974 6840 27030 6896
rect 27710 14592 27766 14648
rect 28998 20576 29054 20632
rect 28906 19896 28962 19952
rect 28538 18692 28594 18728
rect 28538 18672 28540 18692
rect 28540 18672 28592 18692
rect 28592 18672 28594 18692
rect 27986 17856 28042 17912
rect 27986 15544 28042 15600
rect 27986 14320 28042 14376
rect 27342 11092 27344 11112
rect 27344 11092 27396 11112
rect 27396 11092 27398 11112
rect 27342 11056 27398 11092
rect 27434 10512 27490 10568
rect 27342 9288 27398 9344
rect 27710 10240 27766 10296
rect 27618 9016 27674 9072
rect 27250 7112 27306 7168
rect 27342 6840 27398 6896
rect 27342 6024 27398 6080
rect 28354 17040 28410 17096
rect 27802 6568 27858 6624
rect 28262 10512 28318 10568
rect 28446 9444 28502 9480
rect 28446 9424 28448 9444
rect 28448 9424 28500 9444
rect 28500 9424 28502 9444
rect 28262 7792 28318 7848
rect 28262 7268 28318 7304
rect 28262 7248 28264 7268
rect 28264 7248 28316 7268
rect 28316 7248 28318 7268
rect 28814 10512 28870 10568
rect 27710 5788 27712 5808
rect 27712 5788 27764 5808
rect 27764 5788 27766 5808
rect 27710 5752 27766 5788
rect 27526 3052 27582 3088
rect 27526 3032 27528 3052
rect 27528 3032 27580 3052
rect 27580 3032 27582 3052
rect 28722 6604 28724 6624
rect 28724 6604 28776 6624
rect 28776 6604 28778 6624
rect 28722 6568 28778 6604
rect 29550 15952 29606 16008
rect 28262 4120 28318 4176
rect 28722 4428 28724 4448
rect 28724 4428 28776 4448
rect 28776 4428 28778 4448
rect 28722 4392 28778 4428
rect 29274 9424 29330 9480
rect 29182 8744 29238 8800
rect 31114 60052 31116 60072
rect 31116 60052 31168 60072
rect 31168 60052 31170 60072
rect 31114 60016 31170 60052
rect 30654 59472 30710 59528
rect 32218 59916 32220 59936
rect 32220 59916 32272 59936
rect 32272 59916 32274 59936
rect 32218 59880 32274 59916
rect 29918 18400 29974 18456
rect 29826 18128 29882 18184
rect 29826 17756 29828 17776
rect 29828 17756 29880 17776
rect 29880 17756 29882 17776
rect 29826 17720 29882 17756
rect 29734 16224 29790 16280
rect 30010 15272 30066 15328
rect 29826 13096 29882 13152
rect 29734 12144 29790 12200
rect 29458 11192 29514 11248
rect 28998 5344 29054 5400
rect 28998 4664 29054 4720
rect 29550 8200 29606 8256
rect 30470 17176 30526 17232
rect 30286 11328 30342 11384
rect 30102 9016 30158 9072
rect 30010 8880 30066 8936
rect 29918 8608 29974 8664
rect 29642 5652 29644 5672
rect 29644 5652 29696 5672
rect 29696 5652 29698 5672
rect 29642 5616 29698 5652
rect 30286 10104 30342 10160
rect 30378 9424 30434 9480
rect 31390 20304 31446 20360
rect 31390 18672 31446 18728
rect 31206 16496 31262 16552
rect 30286 7656 30342 7712
rect 30654 8880 30710 8936
rect 30654 6976 30710 7032
rect 30930 13368 30986 13424
rect 31022 12688 31078 12744
rect 31666 20440 31722 20496
rect 31942 14864 31998 14920
rect 31850 14320 31906 14376
rect 30746 4800 30802 4856
rect 31850 13096 31906 13152
rect 31942 11736 31998 11792
rect 31574 9016 31630 9072
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 32678 42780 32680 42800
rect 32680 42780 32732 42800
rect 32732 42780 32734 42800
rect 32678 42744 32734 42780
rect 32586 24112 32642 24168
rect 32402 18808 32458 18864
rect 32586 18164 32588 18184
rect 32588 18164 32640 18184
rect 32640 18164 32642 18184
rect 32586 18128 32642 18164
rect 32034 10376 32090 10432
rect 32126 9152 32182 9208
rect 31390 8200 31446 8256
rect 31206 7112 31262 7168
rect 31206 6724 31262 6760
rect 31206 6704 31208 6724
rect 31208 6704 31260 6724
rect 31260 6704 31262 6724
rect 31022 3168 31078 3224
rect 31482 4528 31538 4584
rect 31666 8200 31722 8256
rect 31482 3848 31538 3904
rect 31758 3712 31814 3768
rect 32586 13524 32642 13560
rect 32586 13504 32588 13524
rect 32588 13504 32640 13524
rect 32640 13504 32642 13524
rect 32402 8744 32458 8800
rect 33782 20576 33838 20632
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34334 19760 34390 19816
rect 33414 10376 33470 10432
rect 32862 8744 32918 8800
rect 33046 8492 33102 8528
rect 33046 8472 33048 8492
rect 33048 8472 33100 8492
rect 33100 8472 33102 8492
rect 33506 9016 33562 9072
rect 32954 4936 33010 4992
rect 33598 7656 33654 7712
rect 34426 17040 34482 17096
rect 34058 16224 34114 16280
rect 33966 8744 34022 8800
rect 33322 5616 33378 5672
rect 34518 11192 34574 11248
rect 34334 10376 34390 10432
rect 34150 9560 34206 9616
rect 34150 8916 34152 8936
rect 34152 8916 34204 8936
rect 34204 8916 34206 8936
rect 34150 8880 34206 8916
rect 34150 8336 34206 8392
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35254 12688 35310 12744
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34794 11056 34850 11112
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35254 9832 35310 9888
rect 33046 4120 33102 4176
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 37278 15272 37334 15328
rect 37002 13912 37058 13968
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35898 9696 35954 9752
rect 35990 9152 36046 9208
rect 36082 8880 36138 8936
rect 35714 8472 35770 8528
rect 36174 7928 36230 7984
rect 35162 5208 35218 5264
rect 34702 4120 34758 4176
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35898 3984 35954 4040
rect 36174 5208 36230 5264
rect 37830 18672 37886 18728
rect 36542 7928 36598 7984
rect 36358 4664 36414 4720
rect 36450 4120 36506 4176
rect 37186 6160 37242 6216
rect 37094 3984 37150 4040
rect 37738 10104 37794 10160
rect 37554 9424 37610 9480
rect 37462 9288 37518 9344
rect 39210 17604 39266 17640
rect 39210 17584 39212 17604
rect 39212 17584 39264 17604
rect 39264 17584 39266 17604
rect 38198 11600 38254 11656
rect 38014 10104 38070 10160
rect 38382 10512 38438 10568
rect 38658 10920 38714 10976
rect 38014 9560 38070 9616
rect 37922 9424 37978 9480
rect 38290 10104 38346 10160
rect 38566 10104 38622 10160
rect 38382 9868 38384 9888
rect 38384 9868 38436 9888
rect 38436 9868 38438 9888
rect 38382 9832 38438 9868
rect 38566 9832 38622 9888
rect 38290 9152 38346 9208
rect 38566 8744 38622 8800
rect 37830 3712 37886 3768
rect 38382 5772 38438 5808
rect 38382 5752 38384 5772
rect 38384 5752 38436 5772
rect 38436 5752 38438 5772
rect 37738 3304 37794 3360
rect 38198 4156 38200 4176
rect 38200 4156 38252 4176
rect 38252 4156 38254 4176
rect 38198 4120 38254 4156
rect 38198 4004 38254 4040
rect 38198 3984 38200 4004
rect 38200 3984 38252 4004
rect 38252 3984 38254 4004
rect 38290 3712 38346 3768
rect 39118 8608 39174 8664
rect 39302 8608 39358 8664
rect 40038 19080 40094 19136
rect 40222 16632 40278 16688
rect 40038 12280 40094 12336
rect 39946 8064 40002 8120
rect 40130 6840 40186 6896
rect 40774 14864 40830 14920
rect 40774 14184 40830 14240
rect 40406 8880 40462 8936
rect 40406 3612 40408 3632
rect 40408 3612 40460 3632
rect 40460 3612 40462 3632
rect 40406 3576 40462 3612
rect 42062 59336 42118 59392
rect 41510 16632 41566 16688
rect 41142 12180 41144 12200
rect 41144 12180 41196 12200
rect 41196 12180 41198 12200
rect 41142 12144 41198 12180
rect 41050 11872 41106 11928
rect 40958 11736 41014 11792
rect 41510 14864 41566 14920
rect 41786 13932 41842 13968
rect 41786 13912 41788 13932
rect 41788 13912 41840 13932
rect 41840 13912 41842 13932
rect 41510 12280 41566 12336
rect 41326 11736 41382 11792
rect 41510 11736 41566 11792
rect 41326 3848 41382 3904
rect 41694 5344 41750 5400
rect 41786 3984 41842 4040
rect 42430 18400 42486 18456
rect 42430 18128 42486 18184
rect 42246 11892 42302 11928
rect 42246 11872 42248 11892
rect 42248 11872 42300 11892
rect 42300 11872 42302 11892
rect 42338 8608 42394 8664
rect 42706 56616 42762 56672
rect 42706 19080 42762 19136
rect 42890 18692 42946 18728
rect 42890 18672 42892 18692
rect 42892 18672 42944 18692
rect 42944 18672 42946 18692
rect 42890 18536 42946 18592
rect 50300 60954 50356 60956
rect 50380 60954 50436 60956
rect 50460 60954 50516 60956
rect 50540 60954 50596 60956
rect 50300 60902 50346 60954
rect 50346 60902 50356 60954
rect 50380 60902 50410 60954
rect 50410 60902 50422 60954
rect 50422 60902 50436 60954
rect 50460 60902 50474 60954
rect 50474 60902 50486 60954
rect 50486 60902 50516 60954
rect 50540 60902 50550 60954
rect 50550 60902 50596 60954
rect 50300 60900 50356 60902
rect 50380 60900 50436 60902
rect 50460 60900 50516 60902
rect 50540 60900 50596 60902
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 43442 18400 43498 18456
rect 42706 5480 42762 5536
rect 42522 5072 42578 5128
rect 42614 3168 42670 3224
rect 42614 3068 42616 3088
rect 42616 3068 42668 3088
rect 42668 3068 42670 3088
rect 42614 3032 42670 3068
rect 43534 13912 43590 13968
rect 43994 10648 44050 10704
rect 43718 3576 43774 3632
rect 44178 2488 44234 2544
rect 45926 16632 45982 16688
rect 46570 16088 46626 16144
rect 46754 9016 46810 9072
rect 45926 5344 45982 5400
rect 47122 18128 47178 18184
rect 47766 18692 47822 18728
rect 47766 18672 47768 18692
rect 47768 18672 47820 18692
rect 47820 18672 47822 18692
rect 48226 8064 48282 8120
rect 49698 19352 49754 19408
rect 49698 19080 49754 19136
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50434 19116 50436 19136
rect 50436 19116 50488 19136
rect 50488 19116 50490 19136
rect 50434 19080 50490 19116
rect 51262 19388 51264 19408
rect 51264 19388 51316 19408
rect 51316 19388 51318 19408
rect 51262 19352 51318 19388
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 52642 19216 52698 19272
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 52366 8472 52422 8528
rect 52366 6160 52422 6216
rect 52458 2352 52514 2408
rect 53378 21020 53380 21040
rect 53380 21020 53432 21040
rect 53432 21020 53434 21040
rect 53378 20984 53434 21020
rect 53838 21004 53894 21040
rect 53838 20984 53840 21004
rect 53840 20984 53892 21004
rect 53892 20984 53894 21004
rect 54666 19352 54722 19408
rect 55494 20848 55550 20904
rect 55310 3848 55366 3904
rect 58070 59880 58126 59936
rect 58070 59336 58126 59392
rect 58806 62600 58862 62656
rect 58898 62056 58954 62112
rect 58990 61512 59046 61568
rect 58990 60968 59046 61024
rect 58990 60424 59046 60480
rect 58162 58792 58218 58848
rect 57978 57704 58034 57760
rect 56598 12824 56654 12880
rect 57978 49000 58034 49056
rect 58346 56072 58402 56128
rect 58346 54440 58402 54496
rect 58346 52844 58348 52864
rect 58348 52844 58400 52864
rect 58400 52844 58402 52864
rect 58346 52808 58402 52844
rect 58346 51176 58402 51232
rect 58162 47912 58218 47968
rect 58070 47368 58126 47424
rect 58162 46280 58218 46336
rect 58162 43016 58218 43072
rect 57978 41928 58034 41984
rect 57978 38664 58034 38720
rect 58162 38120 58218 38176
rect 58070 37576 58126 37632
rect 58162 36488 58218 36544
rect 57978 35944 58034 36000
rect 58162 34856 58218 34912
rect 58070 31048 58126 31104
rect 58162 29960 58218 30016
rect 58162 28328 58218 28384
rect 58162 26696 58218 26752
rect 58070 26152 58126 26208
rect 58162 25064 58218 25120
rect 58070 24520 58126 24576
rect 58162 22888 58218 22944
rect 58162 21800 58218 21856
rect 58070 21256 58126 21312
rect 58070 15544 58126 15600
rect 58162 15272 58218 15328
rect 58070 15000 58126 15056
rect 57978 14728 58034 14784
rect 58162 13640 58218 13696
rect 58162 12008 58218 12064
rect 58162 10376 58218 10432
rect 58714 44104 58770 44160
rect 58714 40840 58770 40896
rect 58714 40332 58716 40352
rect 58716 40332 58768 40352
rect 58768 40332 58770 40352
rect 58714 40296 58770 40332
rect 58806 17992 58862 18048
rect 58990 58248 59046 58304
rect 58990 57160 59046 57216
rect 58990 56616 59046 56672
rect 58990 49544 59046 49600
rect 58990 45736 59046 45792
rect 58990 44648 59046 44704
rect 58990 42472 59046 42528
rect 58990 41384 59046 41440
rect 58990 39752 59046 39808
rect 58990 39208 59046 39264
rect 58990 34312 59046 34368
rect 58990 33224 59046 33280
rect 58990 32680 59046 32736
rect 58990 31592 59046 31648
rect 58990 29416 59046 29472
rect 58990 27784 59046 27840
rect 58990 23432 59046 23488
rect 58990 20168 59046 20224
rect 58990 19624 59046 19680
rect 58990 18572 58992 18592
rect 58992 18572 59044 18592
rect 59044 18572 59046 18592
rect 58990 18536 59046 18572
rect 59082 17584 59138 17640
rect 58990 16904 59046 16960
rect 58990 16360 59046 16416
rect 58990 13096 59046 13152
rect 58990 11464 59046 11520
rect 58990 9832 59046 9888
rect 58990 8744 59046 8800
rect 58990 8200 59046 8256
rect 58898 7112 58954 7168
rect 58070 6568 58126 6624
rect 58990 5480 59046 5536
rect 58070 4936 58126 4992
rect 58162 3304 58218 3360
rect 58990 3848 59046 3904
rect 58990 2760 59046 2816
rect 58898 2216 58954 2272
rect 58806 1672 58862 1728
rect 56506 1128 56562 1184
<< metal3 >>
rect 58801 62658 58867 62661
rect 59200 62658 60000 62688
rect 58801 62656 60000 62658
rect 58801 62600 58806 62656
rect 58862 62600 60000 62656
rect 58801 62598 60000 62600
rect 58801 62595 58867 62598
rect 59200 62568 60000 62598
rect 58893 62114 58959 62117
rect 59200 62114 60000 62144
rect 58893 62112 60000 62114
rect 58893 62056 58898 62112
rect 58954 62056 60000 62112
rect 58893 62054 60000 62056
rect 58893 62051 58959 62054
rect 59200 62024 60000 62054
rect 0 61842 800 61872
rect 933 61842 999 61845
rect 0 61840 999 61842
rect 0 61784 938 61840
rect 994 61784 999 61840
rect 0 61782 999 61784
rect 0 61752 800 61782
rect 933 61779 999 61782
rect 58985 61570 59051 61573
rect 59200 61570 60000 61600
rect 58985 61568 60000 61570
rect 58985 61512 58990 61568
rect 59046 61512 60000 61568
rect 58985 61510 60000 61512
rect 58985 61507 59051 61510
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 34930 61504 35246 61505
rect 34930 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35246 61504
rect 59200 61480 60000 61510
rect 34930 61439 35246 61440
rect 0 61162 800 61192
rect 1025 61162 1091 61165
rect 0 61160 1091 61162
rect 0 61104 1030 61160
rect 1086 61104 1091 61160
rect 0 61102 1091 61104
rect 0 61072 800 61102
rect 1025 61099 1091 61102
rect 58985 61026 59051 61029
rect 59200 61026 60000 61056
rect 58985 61024 60000 61026
rect 58985 60968 58990 61024
rect 59046 60968 60000 61024
rect 58985 60966 60000 60968
rect 58985 60963 59051 60966
rect 19570 60960 19886 60961
rect 19570 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19886 60960
rect 19570 60895 19886 60896
rect 50290 60960 50606 60961
rect 50290 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50606 60960
rect 59200 60936 60000 60966
rect 50290 60895 50606 60896
rect 20478 60692 20484 60756
rect 20548 60754 20554 60756
rect 22185 60754 22251 60757
rect 20548 60752 22251 60754
rect 20548 60696 22190 60752
rect 22246 60696 22251 60752
rect 20548 60694 22251 60696
rect 20548 60692 20554 60694
rect 22185 60691 22251 60694
rect 0 60482 800 60512
rect 933 60482 999 60485
rect 0 60480 999 60482
rect 0 60424 938 60480
rect 994 60424 999 60480
rect 0 60422 999 60424
rect 0 60392 800 60422
rect 933 60419 999 60422
rect 58985 60482 59051 60485
rect 59200 60482 60000 60512
rect 58985 60480 60000 60482
rect 58985 60424 58990 60480
rect 59046 60424 60000 60480
rect 58985 60422 60000 60424
rect 58985 60419 59051 60422
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 34930 60416 35246 60417
rect 34930 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35246 60416
rect 59200 60392 60000 60422
rect 34930 60351 35246 60352
rect 31109 60076 31175 60077
rect 31109 60074 31156 60076
rect 31064 60072 31156 60074
rect 31064 60016 31114 60072
rect 31064 60014 31156 60016
rect 31109 60012 31156 60014
rect 31220 60012 31226 60076
rect 31109 60011 31175 60012
rect 29085 59940 29151 59941
rect 29085 59938 29132 59940
rect 29040 59936 29132 59938
rect 29040 59880 29090 59936
rect 29040 59878 29132 59880
rect 29085 59876 29132 59878
rect 29196 59876 29202 59940
rect 32213 59938 32279 59941
rect 32438 59938 32444 59940
rect 32213 59936 32444 59938
rect 32213 59880 32218 59936
rect 32274 59880 32444 59936
rect 32213 59878 32444 59880
rect 29085 59875 29151 59876
rect 32213 59875 32279 59878
rect 32438 59876 32444 59878
rect 32508 59876 32514 59940
rect 58065 59938 58131 59941
rect 59200 59938 60000 59968
rect 58065 59936 60000 59938
rect 58065 59880 58070 59936
rect 58126 59880 60000 59936
rect 58065 59878 60000 59880
rect 58065 59875 58131 59878
rect 19570 59872 19886 59873
rect 0 59802 800 59832
rect 19570 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19886 59872
rect 19570 59807 19886 59808
rect 50290 59872 50606 59873
rect 50290 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50606 59872
rect 59200 59848 60000 59878
rect 50290 59807 50606 59808
rect 933 59802 999 59805
rect 0 59800 999 59802
rect 0 59744 938 59800
rect 994 59744 999 59800
rect 0 59742 999 59744
rect 0 59712 800 59742
rect 933 59739 999 59742
rect 29729 59530 29795 59533
rect 30649 59530 30715 59533
rect 29729 59528 30715 59530
rect 29729 59472 29734 59528
rect 29790 59472 30654 59528
rect 30710 59472 30715 59528
rect 29729 59470 30715 59472
rect 29729 59467 29795 59470
rect 30649 59467 30715 59470
rect 21817 59394 21883 59397
rect 21950 59394 21956 59396
rect 21817 59392 21956 59394
rect 21817 59336 21822 59392
rect 21878 59336 21956 59392
rect 21817 59334 21956 59336
rect 21817 59331 21883 59334
rect 21950 59332 21956 59334
rect 22020 59332 22026 59396
rect 42057 59394 42123 59397
rect 42558 59394 42564 59396
rect 42057 59392 42564 59394
rect 42057 59336 42062 59392
rect 42118 59336 42564 59392
rect 42057 59334 42564 59336
rect 42057 59331 42123 59334
rect 42558 59332 42564 59334
rect 42628 59332 42634 59396
rect 58065 59394 58131 59397
rect 59200 59394 60000 59424
rect 58065 59392 60000 59394
rect 58065 59336 58070 59392
rect 58126 59336 60000 59392
rect 58065 59334 60000 59336
rect 58065 59331 58131 59334
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 34930 59328 35246 59329
rect 34930 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35246 59328
rect 59200 59304 60000 59334
rect 34930 59263 35246 59264
rect 0 59122 800 59152
rect 933 59122 999 59125
rect 0 59120 999 59122
rect 0 59064 938 59120
rect 994 59064 999 59120
rect 0 59062 999 59064
rect 0 59032 800 59062
rect 933 59059 999 59062
rect 58157 58850 58223 58853
rect 59200 58850 60000 58880
rect 58157 58848 60000 58850
rect 58157 58792 58162 58848
rect 58218 58792 60000 58848
rect 58157 58790 60000 58792
rect 58157 58787 58223 58790
rect 19570 58784 19886 58785
rect 19570 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19886 58784
rect 19570 58719 19886 58720
rect 50290 58784 50606 58785
rect 50290 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50606 58784
rect 59200 58760 60000 58790
rect 50290 58719 50606 58720
rect 0 58442 800 58472
rect 933 58442 999 58445
rect 0 58440 999 58442
rect 0 58384 938 58440
rect 994 58384 999 58440
rect 0 58382 999 58384
rect 0 58352 800 58382
rect 933 58379 999 58382
rect 58985 58306 59051 58309
rect 59200 58306 60000 58336
rect 58985 58304 60000 58306
rect 58985 58248 58990 58304
rect 59046 58248 60000 58304
rect 58985 58246 60000 58248
rect 58985 58243 59051 58246
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 34930 58240 35246 58241
rect 34930 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35246 58240
rect 59200 58216 60000 58246
rect 34930 58175 35246 58176
rect 0 57762 800 57792
rect 933 57762 999 57765
rect 0 57760 999 57762
rect 0 57704 938 57760
rect 994 57704 999 57760
rect 0 57702 999 57704
rect 0 57672 800 57702
rect 933 57699 999 57702
rect 57973 57762 58039 57765
rect 59200 57762 60000 57792
rect 57973 57760 60000 57762
rect 57973 57704 57978 57760
rect 58034 57704 60000 57760
rect 57973 57702 60000 57704
rect 57973 57699 58039 57702
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 59200 57672 60000 57702
rect 50290 57631 50606 57632
rect 58985 57218 59051 57221
rect 59200 57218 60000 57248
rect 58985 57216 60000 57218
rect 58985 57160 58990 57216
rect 59046 57160 60000 57216
rect 58985 57158 60000 57160
rect 58985 57155 59051 57158
rect 4210 57152 4526 57153
rect 0 57082 800 57112
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 59200 57128 60000 57158
rect 34930 57087 35246 57088
rect 933 57082 999 57085
rect 0 57080 999 57082
rect 0 57024 938 57080
rect 994 57024 999 57080
rect 0 57022 999 57024
rect 0 56992 800 57022
rect 933 57019 999 57022
rect 42701 56674 42767 56677
rect 43846 56674 43852 56676
rect 42701 56672 43852 56674
rect 42701 56616 42706 56672
rect 42762 56616 43852 56672
rect 42701 56614 43852 56616
rect 42701 56611 42767 56614
rect 43846 56612 43852 56614
rect 43916 56612 43922 56676
rect 58985 56674 59051 56677
rect 59200 56674 60000 56704
rect 58985 56672 60000 56674
rect 58985 56616 58990 56672
rect 59046 56616 60000 56672
rect 58985 56614 60000 56616
rect 58985 56611 59051 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 59200 56584 60000 56614
rect 50290 56543 50606 56544
rect 0 56402 800 56432
rect 933 56402 999 56405
rect 0 56400 999 56402
rect 0 56344 938 56400
rect 994 56344 999 56400
rect 0 56342 999 56344
rect 0 56312 800 56342
rect 933 56339 999 56342
rect 58341 56130 58407 56133
rect 59200 56130 60000 56160
rect 58341 56128 60000 56130
rect 58341 56072 58346 56128
rect 58402 56072 60000 56128
rect 58341 56070 60000 56072
rect 58341 56067 58407 56070
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 59200 56040 60000 56070
rect 34930 55999 35246 56000
rect 0 55722 800 55752
rect 933 55722 999 55725
rect 0 55720 999 55722
rect 0 55664 938 55720
rect 994 55664 999 55720
rect 0 55662 999 55664
rect 0 55632 800 55662
rect 933 55659 999 55662
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 59200 55496 60000 55616
rect 50290 55455 50606 55456
rect 23933 55314 23999 55317
rect 25262 55314 25268 55316
rect 23933 55312 25268 55314
rect 23933 55256 23938 55312
rect 23994 55256 25268 55312
rect 23933 55254 25268 55256
rect 23933 55251 23999 55254
rect 25262 55252 25268 55254
rect 25332 55252 25338 55316
rect 0 55042 800 55072
rect 933 55042 999 55045
rect 0 55040 999 55042
rect 0 54984 938 55040
rect 994 54984 999 55040
rect 0 54982 999 54984
rect 0 54952 800 54982
rect 933 54979 999 54982
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 59200 54952 60000 55072
rect 34930 54911 35246 54912
rect 58341 54498 58407 54501
rect 59200 54498 60000 54528
rect 58341 54496 60000 54498
rect 58341 54440 58346 54496
rect 58402 54440 60000 54496
rect 58341 54438 60000 54440
rect 58341 54435 58407 54438
rect 19570 54432 19886 54433
rect 0 54362 800 54392
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 59200 54408 60000 54438
rect 50290 54367 50606 54368
rect 933 54362 999 54365
rect 0 54360 999 54362
rect 0 54304 938 54360
rect 994 54304 999 54360
rect 0 54302 999 54304
rect 0 54272 800 54302
rect 933 54299 999 54302
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 59200 53864 60000 53984
rect 34930 53823 35246 53824
rect 0 53682 800 53712
rect 933 53682 999 53685
rect 0 53680 999 53682
rect 0 53624 938 53680
rect 994 53624 999 53680
rect 0 53622 999 53624
rect 0 53592 800 53622
rect 933 53619 999 53622
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 59200 53320 60000 53440
rect 50290 53279 50606 53280
rect 0 53002 800 53032
rect 933 53002 999 53005
rect 0 53000 999 53002
rect 0 52944 938 53000
rect 994 52944 999 53000
rect 0 52942 999 52944
rect 0 52912 800 52942
rect 933 52939 999 52942
rect 58341 52866 58407 52869
rect 59200 52866 60000 52896
rect 58341 52864 60000 52866
rect 58341 52808 58346 52864
rect 58402 52808 60000 52864
rect 58341 52806 60000 52808
rect 58341 52803 58407 52806
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 59200 52776 60000 52806
rect 34930 52735 35246 52736
rect 2037 52594 2103 52597
rect 25078 52594 25084 52596
rect 2037 52592 25084 52594
rect 2037 52536 2042 52592
rect 2098 52536 25084 52592
rect 2037 52534 25084 52536
rect 2037 52531 2103 52534
rect 25078 52532 25084 52534
rect 25148 52532 25154 52596
rect 0 52322 800 52352
rect 933 52322 999 52325
rect 0 52320 999 52322
rect 0 52264 938 52320
rect 994 52264 999 52320
rect 0 52262 999 52264
rect 0 52232 800 52262
rect 933 52259 999 52262
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 59200 52232 60000 52352
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 0 51642 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 59200 51688 60000 51808
rect 34930 51647 35246 51648
rect 933 51642 999 51645
rect 0 51640 999 51642
rect 0 51584 938 51640
rect 994 51584 999 51640
rect 0 51582 999 51584
rect 0 51552 800 51582
rect 933 51579 999 51582
rect 58341 51234 58407 51237
rect 59200 51234 60000 51264
rect 58341 51232 60000 51234
rect 58341 51176 58346 51232
rect 58402 51176 60000 51232
rect 58341 51174 60000 51176
rect 58341 51171 58407 51174
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 59200 51144 60000 51174
rect 50290 51103 50606 51104
rect 0 50962 800 50992
rect 933 50962 999 50965
rect 0 50960 999 50962
rect 0 50904 938 50960
rect 994 50904 999 50960
rect 0 50902 999 50904
rect 0 50872 800 50902
rect 933 50899 999 50902
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 59200 50600 60000 50720
rect 34930 50559 35246 50560
rect 0 50282 800 50312
rect 933 50282 999 50285
rect 0 50280 999 50282
rect 0 50224 938 50280
rect 994 50224 999 50280
rect 0 50222 999 50224
rect 0 50192 800 50222
rect 933 50219 999 50222
rect 17585 50282 17651 50285
rect 35934 50282 35940 50284
rect 17585 50280 35940 50282
rect 17585 50224 17590 50280
rect 17646 50224 35940 50280
rect 17585 50222 35940 50224
rect 17585 50219 17651 50222
rect 35934 50220 35940 50222
rect 36004 50220 36010 50284
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 59200 50056 60000 50176
rect 50290 50015 50606 50016
rect 0 49602 800 49632
rect 933 49602 999 49605
rect 0 49600 999 49602
rect 0 49544 938 49600
rect 994 49544 999 49600
rect 0 49542 999 49544
rect 0 49512 800 49542
rect 933 49539 999 49542
rect 58985 49602 59051 49605
rect 59200 49602 60000 49632
rect 58985 49600 60000 49602
rect 58985 49544 58990 49600
rect 59046 49544 60000 49600
rect 58985 49542 60000 49544
rect 58985 49539 59051 49542
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 59200 49512 60000 49542
rect 34930 49471 35246 49472
rect 57973 49058 58039 49061
rect 59200 49058 60000 49088
rect 57973 49056 60000 49058
rect 57973 49000 57978 49056
rect 58034 49000 60000 49056
rect 57973 48998 60000 49000
rect 57973 48995 58039 48998
rect 19570 48992 19886 48993
rect 0 48922 800 48952
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 59200 48968 60000 48998
rect 50290 48927 50606 48928
rect 933 48922 999 48925
rect 0 48920 999 48922
rect 0 48864 938 48920
rect 994 48864 999 48920
rect 0 48862 999 48864
rect 0 48832 800 48862
rect 933 48859 999 48862
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 59200 48424 60000 48544
rect 34930 48383 35246 48384
rect 0 48242 800 48272
rect 933 48242 999 48245
rect 0 48240 999 48242
rect 0 48184 938 48240
rect 994 48184 999 48240
rect 0 48182 999 48184
rect 0 48152 800 48182
rect 933 48179 999 48182
rect 58157 47970 58223 47973
rect 59200 47970 60000 48000
rect 58157 47968 60000 47970
rect 58157 47912 58162 47968
rect 58218 47912 60000 47968
rect 58157 47910 60000 47912
rect 58157 47907 58223 47910
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 59200 47880 60000 47910
rect 50290 47839 50606 47840
rect 0 47562 800 47592
rect 933 47562 999 47565
rect 0 47560 999 47562
rect 0 47504 938 47560
rect 994 47504 999 47560
rect 0 47502 999 47504
rect 0 47472 800 47502
rect 933 47499 999 47502
rect 15193 47562 15259 47565
rect 38694 47562 38700 47564
rect 15193 47560 38700 47562
rect 15193 47504 15198 47560
rect 15254 47504 38700 47560
rect 15193 47502 38700 47504
rect 15193 47499 15259 47502
rect 38694 47500 38700 47502
rect 38764 47500 38770 47564
rect 58065 47426 58131 47429
rect 59200 47426 60000 47456
rect 58065 47424 60000 47426
rect 58065 47368 58070 47424
rect 58126 47368 60000 47424
rect 58065 47366 60000 47368
rect 58065 47363 58131 47366
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 59200 47336 60000 47366
rect 34930 47295 35246 47296
rect 0 46882 800 46912
rect 933 46882 999 46885
rect 0 46880 999 46882
rect 0 46824 938 46880
rect 994 46824 999 46880
rect 0 46822 999 46824
rect 0 46792 800 46822
rect 933 46819 999 46822
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 59200 46792 60000 46912
rect 50290 46751 50606 46752
rect 58157 46338 58223 46341
rect 59200 46338 60000 46368
rect 58157 46336 60000 46338
rect 58157 46280 58162 46336
rect 58218 46280 60000 46336
rect 58157 46278 60000 46280
rect 58157 46275 58223 46278
rect 4210 46272 4526 46273
rect 0 46202 800 46232
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 59200 46248 60000 46278
rect 34930 46207 35246 46208
rect 933 46202 999 46205
rect 0 46200 999 46202
rect 0 46144 938 46200
rect 994 46144 999 46200
rect 0 46142 999 46144
rect 0 46112 800 46142
rect 933 46139 999 46142
rect 58985 45794 59051 45797
rect 59200 45794 60000 45824
rect 58985 45792 60000 45794
rect 58985 45736 58990 45792
rect 59046 45736 60000 45792
rect 58985 45734 60000 45736
rect 58985 45731 59051 45734
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 59200 45704 60000 45734
rect 50290 45663 50606 45664
rect 0 45522 800 45552
rect 933 45522 999 45525
rect 0 45520 999 45522
rect 0 45464 938 45520
rect 994 45464 999 45520
rect 0 45462 999 45464
rect 0 45432 800 45462
rect 933 45459 999 45462
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 59200 45160 60000 45280
rect 34930 45119 35246 45120
rect 0 44842 800 44872
rect 933 44842 999 44845
rect 0 44840 999 44842
rect 0 44784 938 44840
rect 994 44784 999 44840
rect 0 44782 999 44784
rect 0 44752 800 44782
rect 933 44779 999 44782
rect 1853 44842 1919 44845
rect 37590 44842 37596 44844
rect 1853 44840 37596 44842
rect 1853 44784 1858 44840
rect 1914 44784 37596 44840
rect 1853 44782 37596 44784
rect 1853 44779 1919 44782
rect 37590 44780 37596 44782
rect 37660 44780 37666 44844
rect 58985 44706 59051 44709
rect 59200 44706 60000 44736
rect 58985 44704 60000 44706
rect 58985 44648 58990 44704
rect 59046 44648 60000 44704
rect 58985 44646 60000 44648
rect 58985 44643 59051 44646
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 59200 44616 60000 44646
rect 50290 44575 50606 44576
rect 7741 44298 7807 44301
rect 15878 44298 15884 44300
rect 7741 44296 15884 44298
rect 7741 44240 7746 44296
rect 7802 44240 15884 44296
rect 7741 44238 15884 44240
rect 7741 44235 7807 44238
rect 15878 44236 15884 44238
rect 15948 44236 15954 44300
rect 0 44162 800 44192
rect 933 44162 999 44165
rect 0 44160 999 44162
rect 0 44104 938 44160
rect 994 44104 999 44160
rect 0 44102 999 44104
rect 0 44072 800 44102
rect 933 44099 999 44102
rect 58709 44162 58775 44165
rect 59200 44162 60000 44192
rect 58709 44160 60000 44162
rect 58709 44104 58714 44160
rect 58770 44104 60000 44160
rect 58709 44102 60000 44104
rect 58709 44099 58775 44102
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 59200 44072 60000 44102
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 0 43482 800 43512
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 59200 43528 60000 43648
rect 50290 43487 50606 43488
rect 933 43482 999 43485
rect 0 43480 999 43482
rect 0 43424 938 43480
rect 994 43424 999 43480
rect 0 43422 999 43424
rect 0 43392 800 43422
rect 933 43419 999 43422
rect 58157 43074 58223 43077
rect 59200 43074 60000 43104
rect 58157 43072 60000 43074
rect 58157 43016 58162 43072
rect 58218 43016 60000 43072
rect 58157 43014 60000 43016
rect 58157 43011 58223 43014
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 59200 42984 60000 43014
rect 34930 42943 35246 42944
rect 0 42802 800 42832
rect 933 42802 999 42805
rect 0 42800 999 42802
rect 0 42744 938 42800
rect 994 42744 999 42800
rect 0 42742 999 42744
rect 0 42712 800 42742
rect 933 42739 999 42742
rect 26734 42740 26740 42804
rect 26804 42802 26810 42804
rect 32673 42802 32739 42805
rect 26804 42800 32739 42802
rect 26804 42744 32678 42800
rect 32734 42744 32739 42800
rect 26804 42742 32739 42744
rect 26804 42740 26810 42742
rect 32673 42739 32739 42742
rect 58985 42530 59051 42533
rect 59200 42530 60000 42560
rect 58985 42528 60000 42530
rect 58985 42472 58990 42528
rect 59046 42472 60000 42528
rect 58985 42470 60000 42472
rect 58985 42467 59051 42470
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 59200 42440 60000 42470
rect 50290 42399 50606 42400
rect 0 42122 800 42152
rect 933 42122 999 42125
rect 0 42120 999 42122
rect 0 42064 938 42120
rect 994 42064 999 42120
rect 0 42062 999 42064
rect 0 42032 800 42062
rect 933 42059 999 42062
rect 57973 41986 58039 41989
rect 59200 41986 60000 42016
rect 57973 41984 60000 41986
rect 57973 41928 57978 41984
rect 58034 41928 60000 41984
rect 57973 41926 60000 41928
rect 57973 41923 58039 41926
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 59200 41896 60000 41926
rect 34930 41855 35246 41856
rect 0 41442 800 41472
rect 933 41442 999 41445
rect 0 41440 999 41442
rect 0 41384 938 41440
rect 994 41384 999 41440
rect 0 41382 999 41384
rect 0 41352 800 41382
rect 933 41379 999 41382
rect 58985 41442 59051 41445
rect 59200 41442 60000 41472
rect 58985 41440 60000 41442
rect 58985 41384 58990 41440
rect 59046 41384 60000 41440
rect 58985 41382 60000 41384
rect 58985 41379 59051 41382
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 59200 41352 60000 41382
rect 50290 41311 50606 41312
rect 58709 40898 58775 40901
rect 59200 40898 60000 40928
rect 58709 40896 60000 40898
rect 58709 40840 58714 40896
rect 58770 40840 60000 40896
rect 58709 40838 60000 40840
rect 58709 40835 58775 40838
rect 4210 40832 4526 40833
rect 0 40762 800 40792
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 59200 40808 60000 40838
rect 34930 40767 35246 40768
rect 933 40762 999 40765
rect 0 40760 999 40762
rect 0 40704 938 40760
rect 994 40704 999 40760
rect 0 40702 999 40704
rect 0 40672 800 40702
rect 933 40699 999 40702
rect 58709 40354 58775 40357
rect 59200 40354 60000 40384
rect 58709 40352 60000 40354
rect 58709 40296 58714 40352
rect 58770 40296 60000 40352
rect 58709 40294 60000 40296
rect 58709 40291 58775 40294
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 59200 40264 60000 40294
rect 50290 40223 50606 40224
rect 0 40082 800 40112
rect 933 40082 999 40085
rect 0 40080 999 40082
rect 0 40024 938 40080
rect 994 40024 999 40080
rect 0 40022 999 40024
rect 0 39992 800 40022
rect 933 40019 999 40022
rect 58985 39810 59051 39813
rect 59200 39810 60000 39840
rect 58985 39808 60000 39810
rect 58985 39752 58990 39808
rect 59046 39752 60000 39808
rect 58985 39750 60000 39752
rect 58985 39747 59051 39750
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 59200 39720 60000 39750
rect 34930 39679 35246 39680
rect 0 39402 800 39432
rect 1025 39402 1091 39405
rect 0 39400 1091 39402
rect 0 39344 1030 39400
rect 1086 39344 1091 39400
rect 0 39342 1091 39344
rect 0 39312 800 39342
rect 1025 39339 1091 39342
rect 58985 39266 59051 39269
rect 59200 39266 60000 39296
rect 58985 39264 60000 39266
rect 58985 39208 58990 39264
rect 59046 39208 60000 39264
rect 58985 39206 60000 39208
rect 58985 39203 59051 39206
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 59200 39176 60000 39206
rect 50290 39135 50606 39136
rect 23105 38858 23171 38861
rect 39246 38858 39252 38860
rect 23105 38856 39252 38858
rect 23105 38800 23110 38856
rect 23166 38800 39252 38856
rect 23105 38798 39252 38800
rect 23105 38795 23171 38798
rect 39246 38796 39252 38798
rect 39316 38796 39322 38860
rect 0 38722 800 38752
rect 933 38722 999 38725
rect 0 38720 999 38722
rect 0 38664 938 38720
rect 994 38664 999 38720
rect 0 38662 999 38664
rect 0 38632 800 38662
rect 933 38659 999 38662
rect 22461 38724 22527 38725
rect 22461 38720 22508 38724
rect 22572 38722 22578 38724
rect 57973 38722 58039 38725
rect 59200 38722 60000 38752
rect 22461 38664 22466 38720
rect 22461 38660 22508 38664
rect 22572 38662 22618 38722
rect 57973 38720 60000 38722
rect 57973 38664 57978 38720
rect 58034 38664 60000 38720
rect 57973 38662 60000 38664
rect 22572 38660 22578 38662
rect 22461 38659 22527 38660
rect 57973 38659 58039 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 59200 38632 60000 38662
rect 34930 38591 35246 38592
rect 58157 38178 58223 38181
rect 59200 38178 60000 38208
rect 58157 38176 60000 38178
rect 58157 38120 58162 38176
rect 58218 38120 60000 38176
rect 58157 38118 60000 38120
rect 58157 38115 58223 38118
rect 19570 38112 19886 38113
rect 0 38042 800 38072
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 59200 38088 60000 38118
rect 50290 38047 50606 38048
rect 1025 38042 1091 38045
rect 0 38040 1091 38042
rect 0 37984 1030 38040
rect 1086 37984 1091 38040
rect 0 37982 1091 37984
rect 0 37952 800 37982
rect 1025 37979 1091 37982
rect 20621 37906 20687 37909
rect 21541 37906 21607 37909
rect 25129 37906 25195 37909
rect 20621 37904 25195 37906
rect 20621 37848 20626 37904
rect 20682 37848 21546 37904
rect 21602 37848 25134 37904
rect 25190 37848 25195 37904
rect 20621 37846 25195 37848
rect 20621 37843 20687 37846
rect 21541 37843 21607 37846
rect 25129 37843 25195 37846
rect 23013 37770 23079 37773
rect 23422 37770 23428 37772
rect 23013 37768 23428 37770
rect 23013 37712 23018 37768
rect 23074 37712 23428 37768
rect 23013 37710 23428 37712
rect 23013 37707 23079 37710
rect 23422 37708 23428 37710
rect 23492 37708 23498 37772
rect 58065 37634 58131 37637
rect 59200 37634 60000 37664
rect 58065 37632 60000 37634
rect 58065 37576 58070 37632
rect 58126 37576 60000 37632
rect 58065 37574 60000 37576
rect 58065 37571 58131 37574
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 59200 37544 60000 37574
rect 34930 37503 35246 37504
rect 0 37362 800 37392
rect 933 37362 999 37365
rect 0 37360 999 37362
rect 0 37304 938 37360
rect 994 37304 999 37360
rect 0 37302 999 37304
rect 0 37272 800 37302
rect 933 37299 999 37302
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 59200 37000 60000 37120
rect 50290 36959 50606 36960
rect 0 36682 800 36712
rect 933 36682 999 36685
rect 0 36680 999 36682
rect 0 36624 938 36680
rect 994 36624 999 36680
rect 0 36622 999 36624
rect 0 36592 800 36622
rect 933 36619 999 36622
rect 58157 36546 58223 36549
rect 59200 36546 60000 36576
rect 58157 36544 60000 36546
rect 58157 36488 58162 36544
rect 58218 36488 60000 36544
rect 58157 36486 60000 36488
rect 58157 36483 58223 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 59200 36456 60000 36486
rect 34930 36415 35246 36416
rect 0 36002 800 36032
rect 933 36002 999 36005
rect 0 36000 999 36002
rect 0 35944 938 36000
rect 994 35944 999 36000
rect 0 35942 999 35944
rect 0 35912 800 35942
rect 933 35939 999 35942
rect 57973 36002 58039 36005
rect 59200 36002 60000 36032
rect 57973 36000 60000 36002
rect 57973 35944 57978 36000
rect 58034 35944 60000 36000
rect 57973 35942 60000 35944
rect 57973 35939 58039 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 59200 35912 60000 35942
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 0 35322 800 35352
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 59200 35368 60000 35488
rect 34930 35327 35246 35328
rect 933 35322 999 35325
rect 0 35320 999 35322
rect 0 35264 938 35320
rect 994 35264 999 35320
rect 0 35262 999 35264
rect 0 35232 800 35262
rect 933 35259 999 35262
rect 6177 35186 6243 35189
rect 16798 35186 16804 35188
rect 6177 35184 16804 35186
rect 6177 35128 6182 35184
rect 6238 35128 16804 35184
rect 6177 35126 16804 35128
rect 6177 35123 6243 35126
rect 16798 35124 16804 35126
rect 16868 35124 16874 35188
rect 58157 34914 58223 34917
rect 59200 34914 60000 34944
rect 58157 34912 60000 34914
rect 58157 34856 58162 34912
rect 58218 34856 60000 34912
rect 58157 34854 60000 34856
rect 58157 34851 58223 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 59200 34824 60000 34854
rect 50290 34783 50606 34784
rect 0 34642 800 34672
rect 933 34642 999 34645
rect 0 34640 999 34642
rect 0 34584 938 34640
rect 994 34584 999 34640
rect 0 34582 999 34584
rect 0 34552 800 34582
rect 933 34579 999 34582
rect 17534 34580 17540 34644
rect 17604 34642 17610 34644
rect 20805 34642 20871 34645
rect 17604 34640 20871 34642
rect 17604 34584 20810 34640
rect 20866 34584 20871 34640
rect 17604 34582 20871 34584
rect 17604 34580 17610 34582
rect 20805 34579 20871 34582
rect 24117 34642 24183 34645
rect 24710 34642 24716 34644
rect 24117 34640 24716 34642
rect 24117 34584 24122 34640
rect 24178 34584 24716 34640
rect 24117 34582 24716 34584
rect 24117 34579 24183 34582
rect 24710 34580 24716 34582
rect 24780 34580 24786 34644
rect 58985 34370 59051 34373
rect 59200 34370 60000 34400
rect 58985 34368 60000 34370
rect 58985 34312 58990 34368
rect 59046 34312 60000 34368
rect 58985 34310 60000 34312
rect 58985 34307 59051 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 59200 34280 60000 34310
rect 34930 34239 35246 34240
rect 0 33962 800 33992
rect 933 33962 999 33965
rect 0 33960 999 33962
rect 0 33904 938 33960
rect 994 33904 999 33960
rect 0 33902 999 33904
rect 0 33872 800 33902
rect 933 33899 999 33902
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 59200 33736 60000 33856
rect 50290 33695 50606 33696
rect 21214 33356 21220 33420
rect 21284 33418 21290 33420
rect 22277 33418 22343 33421
rect 21284 33416 22343 33418
rect 21284 33360 22282 33416
rect 22338 33360 22343 33416
rect 21284 33358 22343 33360
rect 21284 33356 21290 33358
rect 22277 33355 22343 33358
rect 0 33282 800 33312
rect 933 33282 999 33285
rect 0 33280 999 33282
rect 0 33224 938 33280
rect 994 33224 999 33280
rect 0 33222 999 33224
rect 0 33192 800 33222
rect 933 33219 999 33222
rect 58985 33282 59051 33285
rect 59200 33282 60000 33312
rect 58985 33280 60000 33282
rect 58985 33224 58990 33280
rect 59046 33224 60000 33280
rect 58985 33222 60000 33224
rect 58985 33219 59051 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 59200 33192 60000 33222
rect 34930 33151 35246 33152
rect 58985 32738 59051 32741
rect 59200 32738 60000 32768
rect 58985 32736 60000 32738
rect 58985 32680 58990 32736
rect 59046 32680 60000 32736
rect 58985 32678 60000 32680
rect 58985 32675 59051 32678
rect 19570 32672 19886 32673
rect 0 32602 800 32632
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 59200 32648 60000 32678
rect 50290 32607 50606 32608
rect 933 32602 999 32605
rect 0 32600 999 32602
rect 0 32544 938 32600
rect 994 32544 999 32600
rect 0 32542 999 32544
rect 0 32512 800 32542
rect 933 32539 999 32542
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 59200 32104 60000 32224
rect 34930 32063 35246 32064
rect 0 31922 800 31952
rect 933 31922 999 31925
rect 0 31920 999 31922
rect 0 31864 938 31920
rect 994 31864 999 31920
rect 0 31862 999 31864
rect 0 31832 800 31862
rect 933 31859 999 31862
rect 58985 31650 59051 31653
rect 59200 31650 60000 31680
rect 58985 31648 60000 31650
rect 58985 31592 58990 31648
rect 59046 31592 60000 31648
rect 58985 31590 60000 31592
rect 58985 31587 59051 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 59200 31560 60000 31590
rect 50290 31519 50606 31520
rect 0 31242 800 31272
rect 933 31242 999 31245
rect 0 31240 999 31242
rect 0 31184 938 31240
rect 994 31184 999 31240
rect 0 31182 999 31184
rect 0 31152 800 31182
rect 933 31179 999 31182
rect 23422 31180 23428 31244
rect 23492 31242 23498 31244
rect 41822 31242 41828 31244
rect 23492 31182 41828 31242
rect 23492 31180 23498 31182
rect 41822 31180 41828 31182
rect 41892 31180 41898 31244
rect 58065 31106 58131 31109
rect 59200 31106 60000 31136
rect 58065 31104 60000 31106
rect 58065 31048 58070 31104
rect 58126 31048 60000 31104
rect 58065 31046 60000 31048
rect 58065 31043 58131 31046
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 59200 31016 60000 31046
rect 34930 30975 35246 30976
rect 0 30562 800 30592
rect 933 30562 999 30565
rect 0 30560 999 30562
rect 0 30504 938 30560
rect 994 30504 999 30560
rect 0 30502 999 30504
rect 0 30472 800 30502
rect 933 30499 999 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 59200 30472 60000 30592
rect 50290 30431 50606 30432
rect 58157 30018 58223 30021
rect 59200 30018 60000 30048
rect 58157 30016 60000 30018
rect 58157 29960 58162 30016
rect 58218 29960 60000 30016
rect 58157 29958 60000 29960
rect 58157 29955 58223 29958
rect 4210 29952 4526 29953
rect 0 29882 800 29912
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 59200 29928 60000 29958
rect 34930 29887 35246 29888
rect 933 29882 999 29885
rect 0 29880 999 29882
rect 0 29824 938 29880
rect 994 29824 999 29880
rect 0 29822 999 29824
rect 0 29792 800 29822
rect 933 29819 999 29822
rect 21950 29820 21956 29884
rect 22020 29882 22026 29884
rect 22645 29882 22711 29885
rect 22020 29880 22711 29882
rect 22020 29824 22650 29880
rect 22706 29824 22711 29880
rect 22020 29822 22711 29824
rect 22020 29820 22026 29822
rect 22645 29819 22711 29822
rect 58985 29474 59051 29477
rect 59200 29474 60000 29504
rect 58985 29472 60000 29474
rect 58985 29416 58990 29472
rect 59046 29416 60000 29472
rect 58985 29414 60000 29416
rect 58985 29411 59051 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 59200 29384 60000 29414
rect 50290 29343 50606 29344
rect 0 29202 800 29232
rect 933 29202 999 29205
rect 0 29200 999 29202
rect 0 29144 938 29200
rect 994 29144 999 29200
rect 0 29142 999 29144
rect 0 29112 800 29142
rect 933 29139 999 29142
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 59200 28840 60000 28960
rect 34930 28799 35246 28800
rect 0 28522 800 28552
rect 933 28522 999 28525
rect 0 28520 999 28522
rect 0 28464 938 28520
rect 994 28464 999 28520
rect 0 28462 999 28464
rect 0 28432 800 28462
rect 933 28459 999 28462
rect 58157 28386 58223 28389
rect 59200 28386 60000 28416
rect 58157 28384 60000 28386
rect 58157 28328 58162 28384
rect 58218 28328 60000 28384
rect 58157 28326 60000 28328
rect 58157 28323 58223 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 59200 28296 60000 28326
rect 50290 28255 50606 28256
rect 0 27842 800 27872
rect 933 27842 999 27845
rect 0 27840 999 27842
rect 0 27784 938 27840
rect 994 27784 999 27840
rect 0 27782 999 27784
rect 0 27752 800 27782
rect 933 27779 999 27782
rect 58985 27842 59051 27845
rect 59200 27842 60000 27872
rect 58985 27840 60000 27842
rect 58985 27784 58990 27840
rect 59046 27784 60000 27840
rect 58985 27782 60000 27784
rect 58985 27779 59051 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 59200 27752 60000 27782
rect 34930 27711 35246 27712
rect 23749 27706 23815 27709
rect 25221 27706 25287 27709
rect 23749 27704 25287 27706
rect 23749 27648 23754 27704
rect 23810 27648 25226 27704
rect 25282 27648 25287 27704
rect 23749 27646 25287 27648
rect 23749 27643 23815 27646
rect 25221 27643 25287 27646
rect 19570 27232 19886 27233
rect 0 27162 800 27192
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 59200 27208 60000 27328
rect 50290 27167 50606 27168
rect 933 27162 999 27165
rect 0 27160 999 27162
rect 0 27104 938 27160
rect 994 27104 999 27160
rect 0 27102 999 27104
rect 0 27072 800 27102
rect 933 27099 999 27102
rect 58157 26754 58223 26757
rect 59200 26754 60000 26784
rect 58157 26752 60000 26754
rect 58157 26696 58162 26752
rect 58218 26696 60000 26752
rect 58157 26694 60000 26696
rect 58157 26691 58223 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 59200 26664 60000 26694
rect 34930 26623 35246 26624
rect 0 26482 800 26512
rect 933 26482 999 26485
rect 0 26480 999 26482
rect 0 26424 938 26480
rect 994 26424 999 26480
rect 0 26422 999 26424
rect 0 26392 800 26422
rect 933 26419 999 26422
rect 58065 26210 58131 26213
rect 59200 26210 60000 26240
rect 58065 26208 60000 26210
rect 58065 26152 58070 26208
rect 58126 26152 60000 26208
rect 58065 26150 60000 26152
rect 58065 26147 58131 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 59200 26120 60000 26150
rect 50290 26079 50606 26080
rect 0 25802 800 25832
rect 933 25802 999 25805
rect 0 25800 999 25802
rect 0 25744 938 25800
rect 994 25744 999 25800
rect 0 25742 999 25744
rect 0 25712 800 25742
rect 933 25739 999 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 59200 25576 60000 25696
rect 34930 25535 35246 25536
rect 0 25122 800 25152
rect 933 25122 999 25125
rect 0 25120 999 25122
rect 0 25064 938 25120
rect 994 25064 999 25120
rect 0 25062 999 25064
rect 0 25032 800 25062
rect 933 25059 999 25062
rect 58157 25122 58223 25125
rect 59200 25122 60000 25152
rect 58157 25120 60000 25122
rect 58157 25064 58162 25120
rect 58218 25064 60000 25120
rect 58157 25062 60000 25064
rect 58157 25059 58223 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 59200 25032 60000 25062
rect 50290 24991 50606 24992
rect 58065 24578 58131 24581
rect 59200 24578 60000 24608
rect 58065 24576 60000 24578
rect 58065 24520 58070 24576
rect 58126 24520 60000 24576
rect 58065 24518 60000 24520
rect 58065 24515 58131 24518
rect 4210 24512 4526 24513
rect 0 24442 800 24472
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 59200 24488 60000 24518
rect 34930 24447 35246 24448
rect 933 24442 999 24445
rect 0 24440 999 24442
rect 0 24384 938 24440
rect 994 24384 999 24440
rect 0 24382 999 24384
rect 0 24352 800 24382
rect 933 24379 999 24382
rect 32581 24170 32647 24173
rect 40534 24170 40540 24172
rect 32581 24168 40540 24170
rect 32581 24112 32586 24168
rect 32642 24112 40540 24168
rect 32581 24110 40540 24112
rect 32581 24107 32647 24110
rect 40534 24108 40540 24110
rect 40604 24108 40610 24172
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 59200 23944 60000 24064
rect 50290 23903 50606 23904
rect 0 23762 800 23792
rect 933 23762 999 23765
rect 0 23760 999 23762
rect 0 23704 938 23760
rect 994 23704 999 23760
rect 0 23702 999 23704
rect 0 23672 800 23702
rect 933 23699 999 23702
rect 58985 23490 59051 23493
rect 59200 23490 60000 23520
rect 58985 23488 60000 23490
rect 58985 23432 58990 23488
rect 59046 23432 60000 23488
rect 58985 23430 60000 23432
rect 58985 23427 59051 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 59200 23400 60000 23430
rect 34930 23359 35246 23360
rect 0 23082 800 23112
rect 933 23082 999 23085
rect 0 23080 999 23082
rect 0 23024 938 23080
rect 994 23024 999 23080
rect 0 23022 999 23024
rect 0 22992 800 23022
rect 933 23019 999 23022
rect 58157 22946 58223 22949
rect 59200 22946 60000 22976
rect 58157 22944 60000 22946
rect 58157 22888 58162 22944
rect 58218 22888 60000 22944
rect 58157 22886 60000 22888
rect 58157 22883 58223 22886
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 59200 22856 60000 22886
rect 50290 22815 50606 22816
rect 0 22402 800 22432
rect 933 22402 999 22405
rect 0 22400 999 22402
rect 0 22344 938 22400
rect 994 22344 999 22400
rect 0 22342 999 22344
rect 0 22312 800 22342
rect 933 22339 999 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 59200 22312 60000 22432
rect 34930 22271 35246 22272
rect 58157 21858 58223 21861
rect 59200 21858 60000 21888
rect 58157 21856 60000 21858
rect 58157 21800 58162 21856
rect 58218 21800 60000 21856
rect 58157 21798 60000 21800
rect 58157 21795 58223 21798
rect 19570 21792 19886 21793
rect 0 21722 800 21752
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 59200 21768 60000 21798
rect 50290 21727 50606 21728
rect 933 21722 999 21725
rect 0 21720 999 21722
rect 0 21664 938 21720
rect 994 21664 999 21720
rect 0 21662 999 21664
rect 0 21632 800 21662
rect 933 21659 999 21662
rect 19701 21314 19767 21317
rect 26141 21314 26207 21317
rect 19701 21312 26207 21314
rect 19701 21256 19706 21312
rect 19762 21256 26146 21312
rect 26202 21256 26207 21312
rect 19701 21254 26207 21256
rect 19701 21251 19767 21254
rect 26141 21251 26207 21254
rect 58065 21314 58131 21317
rect 59200 21314 60000 21344
rect 58065 21312 60000 21314
rect 58065 21256 58070 21312
rect 58126 21256 60000 21312
rect 58065 21254 60000 21256
rect 58065 21251 58131 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 59200 21224 60000 21254
rect 34930 21183 35246 21184
rect 0 21042 800 21072
rect 933 21042 999 21045
rect 0 21040 999 21042
rect 0 20984 938 21040
rect 994 20984 999 21040
rect 0 20982 999 20984
rect 0 20952 800 20982
rect 933 20979 999 20982
rect 20069 21042 20135 21045
rect 25773 21042 25839 21045
rect 26785 21042 26851 21045
rect 20069 21040 26851 21042
rect 20069 20984 20074 21040
rect 20130 20984 25778 21040
rect 25834 20984 26790 21040
rect 26846 20984 26851 21040
rect 20069 20982 26851 20984
rect 20069 20979 20135 20982
rect 25773 20979 25839 20982
rect 26785 20979 26851 20982
rect 53373 21042 53439 21045
rect 53833 21042 53899 21045
rect 53373 21040 53899 21042
rect 53373 20984 53378 21040
rect 53434 20984 53838 21040
rect 53894 20984 53899 21040
rect 53373 20982 53899 20984
rect 53373 20979 53439 20982
rect 53833 20979 53899 20982
rect 24025 20906 24091 20909
rect 55489 20906 55555 20909
rect 24025 20904 55555 20906
rect 24025 20848 24030 20904
rect 24086 20848 55494 20904
rect 55550 20848 55555 20904
rect 24025 20846 55555 20848
rect 24025 20843 24091 20846
rect 55489 20843 55555 20846
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 59200 20680 60000 20800
rect 50290 20639 50606 20640
rect 28993 20634 29059 20637
rect 33777 20634 33843 20637
rect 28993 20632 33843 20634
rect 28993 20576 28998 20632
rect 29054 20576 33782 20632
rect 33838 20576 33843 20632
rect 28993 20574 33843 20576
rect 28993 20571 29059 20574
rect 33777 20571 33843 20574
rect 9673 20498 9739 20501
rect 25957 20498 26023 20501
rect 31661 20498 31727 20501
rect 9673 20496 31727 20498
rect 9673 20440 9678 20496
rect 9734 20440 25962 20496
rect 26018 20440 31666 20496
rect 31722 20440 31727 20496
rect 9673 20438 31727 20440
rect 9673 20435 9739 20438
rect 25957 20435 26023 20438
rect 31661 20435 31727 20438
rect 0 20362 800 20392
rect 933 20362 999 20365
rect 0 20360 999 20362
rect 0 20304 938 20360
rect 994 20304 999 20360
rect 0 20302 999 20304
rect 0 20272 800 20302
rect 933 20299 999 20302
rect 18137 20362 18203 20365
rect 31385 20362 31451 20365
rect 18137 20360 31451 20362
rect 18137 20304 18142 20360
rect 18198 20304 31390 20360
rect 31446 20304 31451 20360
rect 18137 20302 31451 20304
rect 18137 20299 18203 20302
rect 31385 20299 31451 20302
rect 58985 20226 59051 20229
rect 59200 20226 60000 20256
rect 58985 20224 60000 20226
rect 58985 20168 58990 20224
rect 59046 20168 60000 20224
rect 58985 20166 60000 20168
rect 58985 20163 59051 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 59200 20136 60000 20166
rect 34930 20095 35246 20096
rect 17953 20090 18019 20093
rect 26141 20090 26207 20093
rect 17953 20088 26207 20090
rect 17953 20032 17958 20088
rect 18014 20032 26146 20088
rect 26202 20032 26207 20088
rect 17953 20030 26207 20032
rect 17953 20027 18019 20030
rect 26141 20027 26207 20030
rect 17309 19954 17375 19957
rect 28901 19954 28967 19957
rect 17309 19952 28967 19954
rect 17309 19896 17314 19952
rect 17370 19896 28906 19952
rect 28962 19896 28967 19952
rect 17309 19894 28967 19896
rect 17309 19891 17375 19894
rect 28901 19891 28967 19894
rect 22185 19818 22251 19821
rect 22318 19818 22324 19820
rect 22185 19816 22324 19818
rect 22185 19760 22190 19816
rect 22246 19760 22324 19816
rect 22185 19758 22324 19760
rect 22185 19755 22251 19758
rect 22318 19756 22324 19758
rect 22388 19818 22394 19820
rect 23197 19818 23263 19821
rect 22388 19816 23263 19818
rect 22388 19760 23202 19816
rect 23258 19760 23263 19816
rect 22388 19758 23263 19760
rect 22388 19756 22394 19758
rect 23197 19755 23263 19758
rect 27521 19818 27587 19821
rect 34329 19818 34395 19821
rect 27521 19816 34395 19818
rect 27521 19760 27526 19816
rect 27582 19760 34334 19816
rect 34390 19760 34395 19816
rect 27521 19758 34395 19760
rect 27521 19755 27587 19758
rect 34329 19755 34395 19758
rect 0 19682 800 19712
rect 933 19682 999 19685
rect 0 19680 999 19682
rect 0 19624 938 19680
rect 994 19624 999 19680
rect 0 19622 999 19624
rect 0 19592 800 19622
rect 933 19619 999 19622
rect 58985 19682 59051 19685
rect 59200 19682 60000 19712
rect 58985 19680 60000 19682
rect 58985 19624 58990 19680
rect 59046 19624 60000 19680
rect 58985 19622 60000 19624
rect 58985 19619 59051 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 59200 19592 60000 19622
rect 50290 19551 50606 19552
rect 17217 19410 17283 19413
rect 25589 19410 25655 19413
rect 17217 19408 25655 19410
rect 17217 19352 17222 19408
rect 17278 19352 25594 19408
rect 25650 19352 25655 19408
rect 17217 19350 25655 19352
rect 17217 19347 17283 19350
rect 25589 19347 25655 19350
rect 49693 19410 49759 19413
rect 51257 19410 51323 19413
rect 54661 19410 54727 19413
rect 49693 19408 54727 19410
rect 49693 19352 49698 19408
rect 49754 19352 51262 19408
rect 51318 19352 54666 19408
rect 54722 19352 54727 19408
rect 49693 19350 54727 19352
rect 49693 19347 49759 19350
rect 51257 19347 51323 19350
rect 54661 19347 54727 19350
rect 19885 19274 19951 19277
rect 21173 19274 21239 19277
rect 19885 19272 21239 19274
rect 19885 19216 19890 19272
rect 19946 19216 21178 19272
rect 21234 19216 21239 19272
rect 19885 19214 21239 19216
rect 19885 19211 19951 19214
rect 21173 19211 21239 19214
rect 24669 19274 24735 19277
rect 52637 19274 52703 19277
rect 24669 19272 52703 19274
rect 24669 19216 24674 19272
rect 24730 19216 52642 19272
rect 52698 19216 52703 19272
rect 24669 19214 52703 19216
rect 24669 19211 24735 19214
rect 52637 19211 52703 19214
rect 40033 19138 40099 19141
rect 42701 19138 42767 19141
rect 40033 19136 42767 19138
rect 40033 19080 40038 19136
rect 40094 19080 42706 19136
rect 42762 19080 42767 19136
rect 40033 19078 42767 19080
rect 40033 19075 40099 19078
rect 42701 19075 42767 19078
rect 49693 19138 49759 19141
rect 50429 19138 50495 19141
rect 49693 19136 50495 19138
rect 49693 19080 49698 19136
rect 49754 19080 50434 19136
rect 50490 19080 50495 19136
rect 49693 19078 50495 19080
rect 49693 19075 49759 19078
rect 50429 19075 50495 19078
rect 4210 19072 4526 19073
rect 0 19002 800 19032
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 59200 19048 60000 19168
rect 34930 19007 35246 19008
rect 933 19002 999 19005
rect 0 19000 999 19002
rect 0 18944 938 19000
rect 994 18944 999 19000
rect 0 18942 999 18944
rect 0 18912 800 18942
rect 933 18939 999 18942
rect 11881 19002 11947 19005
rect 17217 19002 17283 19005
rect 11881 19000 17283 19002
rect 11881 18944 11886 19000
rect 11942 18944 17222 19000
rect 17278 18944 17283 19000
rect 11881 18942 17283 18944
rect 11881 18939 11947 18942
rect 17217 18939 17283 18942
rect 21449 19002 21515 19005
rect 23197 19002 23263 19005
rect 21449 19000 23263 19002
rect 21449 18944 21454 19000
rect 21510 18944 23202 19000
rect 23258 18944 23263 19000
rect 21449 18942 23263 18944
rect 21449 18939 21515 18942
rect 23197 18939 23263 18942
rect 12617 18866 12683 18869
rect 32397 18866 32463 18869
rect 12617 18864 32463 18866
rect 12617 18808 12622 18864
rect 12678 18808 32402 18864
rect 32458 18808 32463 18864
rect 12617 18806 32463 18808
rect 12617 18803 12683 18806
rect 32397 18803 32463 18806
rect 22829 18730 22895 18733
rect 28533 18730 28599 18733
rect 22829 18728 28599 18730
rect 22829 18672 22834 18728
rect 22890 18672 28538 18728
rect 28594 18672 28599 18728
rect 22829 18670 28599 18672
rect 22829 18667 22895 18670
rect 28533 18667 28599 18670
rect 31385 18730 31451 18733
rect 37825 18730 37891 18733
rect 31385 18728 37891 18730
rect 31385 18672 31390 18728
rect 31446 18672 37830 18728
rect 37886 18672 37891 18728
rect 31385 18670 37891 18672
rect 31385 18667 31451 18670
rect 37825 18667 37891 18670
rect 42885 18730 42951 18733
rect 47761 18730 47827 18733
rect 42885 18728 47827 18730
rect 42885 18672 42890 18728
rect 42946 18672 47766 18728
rect 47822 18672 47827 18728
rect 42885 18670 47827 18672
rect 42885 18667 42951 18670
rect 47761 18667 47827 18670
rect 42885 18594 42951 18597
rect 38610 18592 42951 18594
rect 38610 18536 42890 18592
rect 42946 18536 42951 18592
rect 38610 18534 42951 18536
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 29913 18458 29979 18461
rect 38610 18458 38670 18534
rect 42885 18531 42951 18534
rect 58985 18594 59051 18597
rect 59200 18594 60000 18624
rect 58985 18592 60000 18594
rect 58985 18536 58990 18592
rect 59046 18536 60000 18592
rect 58985 18534 60000 18536
rect 58985 18531 59051 18534
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 59200 18504 60000 18534
rect 50290 18463 50606 18464
rect 29913 18456 38670 18458
rect 29913 18400 29918 18456
rect 29974 18400 38670 18456
rect 29913 18398 38670 18400
rect 42425 18458 42491 18461
rect 43437 18458 43503 18461
rect 42425 18456 43503 18458
rect 42425 18400 42430 18456
rect 42486 18400 43442 18456
rect 43498 18400 43503 18456
rect 42425 18398 43503 18400
rect 29913 18395 29979 18398
rect 42425 18395 42491 18398
rect 43437 18395 43503 18398
rect 0 18322 800 18352
rect 933 18322 999 18325
rect 0 18320 999 18322
rect 0 18264 938 18320
rect 994 18264 999 18320
rect 0 18262 999 18264
rect 0 18232 800 18262
rect 933 18259 999 18262
rect 14457 18186 14523 18189
rect 18137 18186 18203 18189
rect 14457 18184 18203 18186
rect 14457 18128 14462 18184
rect 14518 18128 18142 18184
rect 18198 18128 18203 18184
rect 14457 18126 18203 18128
rect 14457 18123 14523 18126
rect 18137 18123 18203 18126
rect 27286 18124 27292 18188
rect 27356 18186 27362 18188
rect 29821 18186 29887 18189
rect 32581 18186 32647 18189
rect 27356 18184 32647 18186
rect 27356 18128 29826 18184
rect 29882 18128 32586 18184
rect 32642 18128 32647 18184
rect 27356 18126 32647 18128
rect 27356 18124 27362 18126
rect 29821 18123 29887 18126
rect 32581 18123 32647 18126
rect 42425 18186 42491 18189
rect 47117 18186 47183 18189
rect 42425 18184 47183 18186
rect 42425 18128 42430 18184
rect 42486 18128 47122 18184
rect 47178 18128 47183 18184
rect 42425 18126 47183 18128
rect 42425 18123 42491 18126
rect 47117 18123 47183 18126
rect 58801 18050 58867 18053
rect 59200 18050 60000 18080
rect 58801 18048 60000 18050
rect 58801 17992 58806 18048
rect 58862 17992 60000 18048
rect 58801 17990 60000 17992
rect 58801 17987 58867 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 59200 17960 60000 17990
rect 34930 17919 35246 17920
rect 22686 17852 22692 17916
rect 22756 17914 22762 17916
rect 24761 17914 24827 17917
rect 22756 17912 24827 17914
rect 22756 17856 24766 17912
rect 24822 17856 24827 17912
rect 22756 17854 24827 17856
rect 22756 17852 22762 17854
rect 24761 17851 24827 17854
rect 26182 17852 26188 17916
rect 26252 17914 26258 17916
rect 27981 17914 28047 17917
rect 26252 17912 28047 17914
rect 26252 17856 27986 17912
rect 28042 17856 28047 17912
rect 26252 17854 28047 17856
rect 26252 17852 26258 17854
rect 27981 17851 28047 17854
rect 5533 17778 5599 17781
rect 29821 17778 29887 17781
rect 5533 17776 29887 17778
rect 5533 17720 5538 17776
rect 5594 17720 29826 17776
rect 29882 17720 29887 17776
rect 5533 17718 29887 17720
rect 5533 17715 5599 17718
rect 29821 17715 29887 17718
rect 0 17642 800 17672
rect 933 17642 999 17645
rect 27061 17644 27127 17645
rect 27061 17642 27108 17644
rect 0 17640 999 17642
rect 0 17584 938 17640
rect 994 17584 999 17640
rect 0 17582 999 17584
rect 27016 17640 27108 17642
rect 27016 17584 27066 17640
rect 27016 17582 27108 17584
rect 0 17552 800 17582
rect 933 17579 999 17582
rect 27061 17580 27108 17582
rect 27172 17580 27178 17644
rect 39205 17642 39271 17645
rect 59077 17642 59143 17645
rect 39205 17640 59143 17642
rect 39205 17584 39210 17640
rect 39266 17584 59082 17640
rect 59138 17584 59143 17640
rect 39205 17582 59143 17584
rect 27061 17579 27127 17580
rect 39205 17579 39271 17582
rect 59077 17579 59143 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 59200 17416 60000 17536
rect 50290 17375 50606 17376
rect 11237 17234 11303 17237
rect 30465 17234 30531 17237
rect 11237 17232 30531 17234
rect 11237 17176 11242 17232
rect 11298 17176 30470 17232
rect 30526 17176 30531 17232
rect 11237 17174 30531 17176
rect 11237 17171 11303 17174
rect 30465 17171 30531 17174
rect 28349 17098 28415 17101
rect 34421 17098 34487 17101
rect 28349 17096 34487 17098
rect 28349 17040 28354 17096
rect 28410 17040 34426 17096
rect 34482 17040 34487 17096
rect 28349 17038 34487 17040
rect 28349 17035 28415 17038
rect 34421 17035 34487 17038
rect 0 16962 800 16992
rect 933 16962 999 16965
rect 0 16960 999 16962
rect 0 16904 938 16960
rect 994 16904 999 16960
rect 0 16902 999 16904
rect 0 16872 800 16902
rect 933 16899 999 16902
rect 18321 16962 18387 16965
rect 25313 16962 25379 16965
rect 26049 16962 26115 16965
rect 18321 16960 26115 16962
rect 18321 16904 18326 16960
rect 18382 16904 25318 16960
rect 25374 16904 26054 16960
rect 26110 16904 26115 16960
rect 18321 16902 26115 16904
rect 18321 16899 18387 16902
rect 25313 16899 25379 16902
rect 26049 16899 26115 16902
rect 58985 16962 59051 16965
rect 59200 16962 60000 16992
rect 58985 16960 60000 16962
rect 58985 16904 58990 16960
rect 59046 16904 60000 16960
rect 58985 16902 60000 16904
rect 58985 16899 59051 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 59200 16872 60000 16902
rect 34930 16831 35246 16832
rect 13445 16690 13511 16693
rect 18781 16690 18847 16693
rect 22829 16692 22895 16693
rect 22829 16690 22876 16692
rect 13445 16688 18847 16690
rect 13445 16632 13450 16688
rect 13506 16632 18786 16688
rect 18842 16632 18847 16688
rect 13445 16630 18847 16632
rect 22784 16688 22876 16690
rect 22784 16632 22834 16688
rect 22784 16630 22876 16632
rect 13445 16627 13511 16630
rect 18781 16627 18847 16630
rect 22829 16628 22876 16630
rect 22940 16628 22946 16692
rect 40217 16690 40283 16693
rect 41505 16690 41571 16693
rect 45921 16690 45987 16693
rect 40217 16688 45987 16690
rect 40217 16632 40222 16688
rect 40278 16632 41510 16688
rect 41566 16632 45926 16688
rect 45982 16632 45987 16688
rect 40217 16630 45987 16632
rect 22829 16627 22895 16628
rect 40217 16627 40283 16630
rect 41505 16627 41571 16630
rect 45921 16627 45987 16630
rect 13353 16554 13419 16557
rect 31201 16554 31267 16557
rect 13353 16552 31267 16554
rect 13353 16496 13358 16552
rect 13414 16496 31206 16552
rect 31262 16496 31267 16552
rect 13353 16494 31267 16496
rect 13353 16491 13419 16494
rect 31201 16491 31267 16494
rect 22737 16418 22803 16421
rect 25405 16418 25471 16421
rect 22737 16416 25471 16418
rect 22737 16360 22742 16416
rect 22798 16360 25410 16416
rect 25466 16360 25471 16416
rect 22737 16358 25471 16360
rect 22737 16355 22803 16358
rect 25405 16355 25471 16358
rect 58985 16418 59051 16421
rect 59200 16418 60000 16448
rect 58985 16416 60000 16418
rect 58985 16360 58990 16416
rect 59046 16360 60000 16416
rect 58985 16358 60000 16360
rect 58985 16355 59051 16358
rect 19570 16352 19886 16353
rect 0 16282 800 16312
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 59200 16328 60000 16358
rect 50290 16287 50606 16288
rect 933 16282 999 16285
rect 0 16280 999 16282
rect 0 16224 938 16280
rect 994 16224 999 16280
rect 0 16222 999 16224
rect 0 16192 800 16222
rect 933 16219 999 16222
rect 29729 16282 29795 16285
rect 34053 16282 34119 16285
rect 29729 16280 34119 16282
rect 29729 16224 29734 16280
rect 29790 16224 34058 16280
rect 34114 16224 34119 16280
rect 29729 16222 34119 16224
rect 29729 16219 29795 16222
rect 34053 16219 34119 16222
rect 13813 16146 13879 16149
rect 46565 16146 46631 16149
rect 13813 16144 46631 16146
rect 13813 16088 13818 16144
rect 13874 16088 46570 16144
rect 46626 16088 46631 16144
rect 13813 16086 46631 16088
rect 13813 16083 13879 16086
rect 46565 16083 46631 16086
rect 16481 16010 16547 16013
rect 29545 16010 29611 16013
rect 16481 16008 29611 16010
rect 16481 15952 16486 16008
rect 16542 15952 29550 16008
rect 29606 15952 29611 16008
rect 16481 15950 29611 15952
rect 16481 15947 16547 15950
rect 29545 15947 29611 15950
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 59200 15784 60000 15904
rect 34930 15743 35246 15744
rect 0 15602 800 15632
rect 933 15602 999 15605
rect 0 15600 999 15602
rect 0 15544 938 15600
rect 994 15544 999 15600
rect 0 15542 999 15544
rect 0 15512 800 15542
rect 933 15539 999 15542
rect 27981 15602 28047 15605
rect 58065 15602 58131 15605
rect 27981 15600 58131 15602
rect 27981 15544 27986 15600
rect 28042 15544 58070 15600
rect 58126 15544 58131 15600
rect 27981 15542 58131 15544
rect 27981 15539 28047 15542
rect 58065 15539 58131 15542
rect 30005 15330 30071 15333
rect 37273 15330 37339 15333
rect 30005 15328 37339 15330
rect 30005 15272 30010 15328
rect 30066 15272 37278 15328
rect 37334 15272 37339 15328
rect 30005 15270 37339 15272
rect 30005 15267 30071 15270
rect 37273 15267 37339 15270
rect 58157 15330 58223 15333
rect 59200 15330 60000 15360
rect 58157 15328 60000 15330
rect 58157 15272 58162 15328
rect 58218 15272 60000 15328
rect 58157 15270 60000 15272
rect 58157 15267 58223 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 59200 15240 60000 15270
rect 50290 15199 50606 15200
rect 25221 15196 25287 15197
rect 25221 15192 25268 15196
rect 25332 15194 25338 15196
rect 25221 15136 25226 15192
rect 25221 15132 25268 15136
rect 25332 15134 25378 15194
rect 25332 15132 25338 15134
rect 25221 15131 25287 15132
rect 25773 15060 25839 15061
rect 25773 15058 25820 15060
rect 25732 15056 25820 15058
rect 25884 15058 25890 15060
rect 58065 15058 58131 15061
rect 25884 15056 58131 15058
rect 25732 15000 25778 15056
rect 25884 15000 58070 15056
rect 58126 15000 58131 15056
rect 25732 14998 25820 15000
rect 25773 14996 25820 14998
rect 25884 14998 58131 15000
rect 25884 14996 25890 14998
rect 25773 14995 25839 14996
rect 58065 14995 58131 14998
rect 0 14922 800 14952
rect 933 14922 999 14925
rect 31937 14922 32003 14925
rect 0 14920 999 14922
rect 0 14864 938 14920
rect 994 14864 999 14920
rect 0 14862 999 14864
rect 0 14832 800 14862
rect 933 14859 999 14862
rect 31894 14920 32003 14922
rect 31894 14864 31942 14920
rect 31998 14864 32003 14920
rect 31894 14859 32003 14864
rect 40769 14922 40835 14925
rect 41505 14922 41571 14925
rect 40769 14920 41571 14922
rect 40769 14864 40774 14920
rect 40830 14864 41510 14920
rect 41566 14864 41571 14920
rect 40769 14862 41571 14864
rect 40769 14859 40835 14862
rect 41505 14859 41571 14862
rect 20621 14786 20687 14789
rect 26693 14786 26759 14789
rect 20621 14784 26759 14786
rect 20621 14728 20626 14784
rect 20682 14728 26698 14784
rect 26754 14728 26759 14784
rect 20621 14726 26759 14728
rect 20621 14723 20687 14726
rect 26693 14723 26759 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 27705 14650 27771 14653
rect 12390 14648 27771 14650
rect 12390 14592 27710 14648
rect 27766 14592 27771 14648
rect 12390 14590 27771 14592
rect 1577 14514 1643 14517
rect 12390 14514 12450 14590
rect 27705 14587 27771 14590
rect 1577 14512 12450 14514
rect 1577 14456 1582 14512
rect 1638 14456 12450 14512
rect 1577 14454 12450 14456
rect 24945 14514 25011 14517
rect 25078 14514 25084 14516
rect 24945 14512 25084 14514
rect 24945 14456 24950 14512
rect 25006 14456 25084 14512
rect 24945 14454 25084 14456
rect 1577 14451 1643 14454
rect 24945 14451 25011 14454
rect 25078 14452 25084 14454
rect 25148 14452 25154 14516
rect 25313 14514 25379 14517
rect 25957 14514 26023 14517
rect 25313 14512 26023 14514
rect 25313 14456 25318 14512
rect 25374 14456 25962 14512
rect 26018 14456 26023 14512
rect 25313 14454 26023 14456
rect 25313 14451 25379 14454
rect 25957 14451 26023 14454
rect 31894 14381 31954 14859
rect 57973 14786 58039 14789
rect 59200 14786 60000 14816
rect 57973 14784 60000 14786
rect 57973 14728 57978 14784
rect 58034 14728 60000 14784
rect 57973 14726 60000 14728
rect 57973 14723 58039 14726
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 59200 14696 60000 14726
rect 34930 14655 35246 14656
rect 22461 14378 22527 14381
rect 27981 14378 28047 14381
rect 22461 14376 28047 14378
rect 22461 14320 22466 14376
rect 22522 14320 27986 14376
rect 28042 14320 28047 14376
rect 22461 14318 28047 14320
rect 22461 14315 22527 14318
rect 27981 14315 28047 14318
rect 31845 14376 31954 14381
rect 31845 14320 31850 14376
rect 31906 14320 31954 14376
rect 31845 14318 31954 14320
rect 31845 14315 31911 14318
rect 0 14242 800 14272
rect 933 14242 999 14245
rect 0 14240 999 14242
rect 0 14184 938 14240
rect 994 14184 999 14240
rect 0 14182 999 14184
rect 0 14152 800 14182
rect 933 14179 999 14182
rect 25313 14242 25379 14245
rect 40769 14242 40835 14245
rect 25313 14240 40835 14242
rect 25313 14184 25318 14240
rect 25374 14184 40774 14240
rect 40830 14184 40835 14240
rect 25313 14182 40835 14184
rect 25313 14179 25379 14182
rect 40769 14179 40835 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 59200 14152 60000 14272
rect 50290 14111 50606 14112
rect 20161 14106 20227 14109
rect 22369 14106 22435 14109
rect 20161 14104 22435 14106
rect 20161 14048 20166 14104
rect 20222 14048 22374 14104
rect 22430 14048 22435 14104
rect 20161 14046 22435 14048
rect 20161 14043 20227 14046
rect 22369 14043 22435 14046
rect 26141 14108 26207 14109
rect 26141 14104 26188 14108
rect 26252 14106 26258 14108
rect 26141 14048 26146 14104
rect 26141 14044 26188 14048
rect 26252 14046 26298 14106
rect 26252 14044 26258 14046
rect 26141 14043 26207 14044
rect 23289 13970 23355 13973
rect 16806 13968 23355 13970
rect 16806 13912 23294 13968
rect 23350 13912 23355 13968
rect 16806 13910 23355 13912
rect 16806 13837 16866 13910
rect 23289 13907 23355 13910
rect 25037 13970 25103 13973
rect 36997 13970 37063 13973
rect 25037 13968 37063 13970
rect 25037 13912 25042 13968
rect 25098 13912 37002 13968
rect 37058 13912 37063 13968
rect 25037 13910 37063 13912
rect 25037 13907 25103 13910
rect 36997 13907 37063 13910
rect 41781 13970 41847 13973
rect 43529 13970 43595 13973
rect 41781 13968 43595 13970
rect 41781 13912 41786 13968
rect 41842 13912 43534 13968
rect 43590 13912 43595 13968
rect 41781 13910 43595 13912
rect 41781 13907 41847 13910
rect 43529 13907 43595 13910
rect 16757 13832 16866 13837
rect 16757 13776 16762 13832
rect 16818 13776 16866 13832
rect 16757 13774 16866 13776
rect 18689 13834 18755 13837
rect 24761 13834 24827 13837
rect 18689 13832 24827 13834
rect 18689 13776 18694 13832
rect 18750 13776 24766 13832
rect 24822 13776 24827 13832
rect 18689 13774 24827 13776
rect 16757 13771 16823 13774
rect 18689 13771 18755 13774
rect 24761 13771 24827 13774
rect 19517 13698 19583 13701
rect 21633 13698 21699 13701
rect 19517 13696 21699 13698
rect 19517 13640 19522 13696
rect 19578 13640 21638 13696
rect 21694 13640 21699 13696
rect 19517 13638 21699 13640
rect 19517 13635 19583 13638
rect 21633 13635 21699 13638
rect 22502 13636 22508 13700
rect 22572 13698 22578 13700
rect 23381 13698 23447 13701
rect 22572 13696 23447 13698
rect 22572 13640 23386 13696
rect 23442 13640 23447 13696
rect 22572 13638 23447 13640
rect 22572 13636 22578 13638
rect 23381 13635 23447 13638
rect 58157 13698 58223 13701
rect 59200 13698 60000 13728
rect 58157 13696 60000 13698
rect 58157 13640 58162 13696
rect 58218 13640 60000 13696
rect 58157 13638 60000 13640
rect 58157 13635 58223 13638
rect 4210 13632 4526 13633
rect 0 13562 800 13592
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 59200 13608 60000 13638
rect 34930 13567 35246 13568
rect 933 13562 999 13565
rect 0 13560 999 13562
rect 0 13504 938 13560
rect 994 13504 999 13560
rect 0 13502 999 13504
rect 0 13472 800 13502
rect 933 13499 999 13502
rect 32438 13500 32444 13564
rect 32508 13562 32514 13564
rect 32581 13562 32647 13565
rect 32508 13560 32647 13562
rect 32508 13504 32586 13560
rect 32642 13504 32647 13560
rect 32508 13502 32647 13504
rect 32508 13500 32514 13502
rect 32581 13499 32647 13502
rect 1577 13426 1643 13429
rect 30925 13426 30991 13429
rect 1577 13424 30991 13426
rect 1577 13368 1582 13424
rect 1638 13368 30930 13424
rect 30986 13368 30991 13424
rect 1577 13366 30991 13368
rect 1577 13363 1643 13366
rect 30925 13363 30991 13366
rect 7005 13290 7071 13293
rect 7005 13288 31770 13290
rect 7005 13232 7010 13288
rect 7066 13232 31770 13288
rect 7005 13230 31770 13232
rect 7005 13227 7071 13230
rect 29494 13092 29500 13156
rect 29564 13154 29570 13156
rect 29821 13154 29887 13157
rect 29564 13152 29887 13154
rect 29564 13096 29826 13152
rect 29882 13096 29887 13152
rect 29564 13094 29887 13096
rect 31710 13154 31770 13230
rect 31845 13154 31911 13157
rect 31710 13152 31911 13154
rect 31710 13096 31850 13152
rect 31906 13096 31911 13152
rect 31710 13094 31911 13096
rect 29564 13092 29570 13094
rect 29821 13091 29887 13094
rect 31845 13091 31911 13094
rect 58985 13154 59051 13157
rect 59200 13154 60000 13184
rect 58985 13152 60000 13154
rect 58985 13096 58990 13152
rect 59046 13096 60000 13152
rect 58985 13094 60000 13096
rect 58985 13091 59051 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 59200 13064 60000 13094
rect 50290 13023 50606 13024
rect 0 12882 800 12912
rect 933 12882 999 12885
rect 0 12880 999 12882
rect 0 12824 938 12880
rect 994 12824 999 12880
rect 0 12822 999 12824
rect 0 12792 800 12822
rect 933 12819 999 12822
rect 21633 12882 21699 12885
rect 22185 12882 22251 12885
rect 26233 12882 26299 12885
rect 56593 12882 56659 12885
rect 21633 12880 22251 12882
rect 21633 12824 21638 12880
rect 21694 12824 22190 12880
rect 22246 12824 22251 12880
rect 21633 12822 22251 12824
rect 21633 12819 21699 12822
rect 22185 12819 22251 12822
rect 22326 12880 56659 12882
rect 22326 12824 26238 12880
rect 26294 12824 56598 12880
rect 56654 12824 56659 12880
rect 22326 12822 56659 12824
rect 15101 12746 15167 12749
rect 17677 12746 17743 12749
rect 15101 12744 17743 12746
rect 15101 12688 15106 12744
rect 15162 12688 17682 12744
rect 17738 12688 17743 12744
rect 15101 12686 17743 12688
rect 15101 12683 15167 12686
rect 17677 12683 17743 12686
rect 18137 12746 18203 12749
rect 18321 12746 18387 12749
rect 18137 12744 18387 12746
rect 18137 12688 18142 12744
rect 18198 12688 18326 12744
rect 18382 12688 18387 12744
rect 18137 12686 18387 12688
rect 18137 12683 18203 12686
rect 18321 12683 18387 12686
rect 21173 12746 21239 12749
rect 22326 12746 22386 12822
rect 26233 12819 26299 12822
rect 56593 12819 56659 12822
rect 21173 12744 22386 12746
rect 21173 12688 21178 12744
rect 21234 12688 22386 12744
rect 21173 12686 22386 12688
rect 21173 12683 21239 12686
rect 22870 12684 22876 12748
rect 22940 12746 22946 12748
rect 23013 12746 23079 12749
rect 22940 12744 23079 12746
rect 22940 12688 23018 12744
rect 23074 12688 23079 12744
rect 22940 12686 23079 12688
rect 22940 12684 22946 12686
rect 23013 12683 23079 12686
rect 31017 12746 31083 12749
rect 35249 12746 35315 12749
rect 31017 12744 35315 12746
rect 31017 12688 31022 12744
rect 31078 12688 35254 12744
rect 35310 12688 35315 12744
rect 31017 12686 35315 12688
rect 31017 12683 31083 12686
rect 35249 12683 35315 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 59200 12520 60000 12640
rect 34930 12479 35246 12480
rect 21817 12474 21883 12477
rect 26509 12474 26575 12477
rect 21817 12472 26575 12474
rect 21817 12416 21822 12472
rect 21878 12416 26514 12472
rect 26570 12416 26575 12472
rect 21817 12414 26575 12416
rect 21817 12411 21883 12414
rect 26509 12411 26575 12414
rect 16665 12338 16731 12341
rect 16798 12338 16804 12340
rect 16665 12336 16804 12338
rect 16665 12280 16670 12336
rect 16726 12280 16804 12336
rect 16665 12278 16804 12280
rect 16665 12275 16731 12278
rect 16798 12276 16804 12278
rect 16868 12276 16874 12340
rect 24301 12338 24367 12341
rect 24710 12338 24716 12340
rect 24301 12336 24716 12338
rect 24301 12280 24306 12336
rect 24362 12280 24716 12336
rect 24301 12278 24716 12280
rect 24301 12275 24367 12278
rect 24710 12276 24716 12278
rect 24780 12338 24786 12340
rect 40033 12338 40099 12341
rect 24780 12336 40418 12338
rect 24780 12280 40038 12336
rect 40094 12280 40418 12336
rect 24780 12278 40418 12280
rect 24780 12276 24786 12278
rect 40033 12275 40099 12278
rect 0 12202 800 12232
rect 933 12202 999 12205
rect 0 12200 999 12202
rect 0 12144 938 12200
rect 994 12144 999 12200
rect 0 12142 999 12144
rect 0 12112 800 12142
rect 933 12139 999 12142
rect 4061 12202 4127 12205
rect 29729 12202 29795 12205
rect 4061 12200 29795 12202
rect 4061 12144 4066 12200
rect 4122 12144 29734 12200
rect 29790 12144 29795 12200
rect 4061 12142 29795 12144
rect 40358 12202 40418 12278
rect 40534 12276 40540 12340
rect 40604 12338 40610 12340
rect 41505 12338 41571 12341
rect 40604 12336 41571 12338
rect 40604 12280 41510 12336
rect 41566 12280 41571 12336
rect 40604 12278 41571 12280
rect 40604 12276 40610 12278
rect 41505 12275 41571 12278
rect 41137 12202 41203 12205
rect 40358 12200 41203 12202
rect 40358 12144 41142 12200
rect 41198 12144 41203 12200
rect 40358 12142 41203 12144
rect 4061 12139 4127 12142
rect 29729 12139 29795 12142
rect 41137 12139 41203 12142
rect 24853 12066 24919 12069
rect 26509 12066 26575 12069
rect 24853 12064 26575 12066
rect 24853 12008 24858 12064
rect 24914 12008 26514 12064
rect 26570 12008 26575 12064
rect 24853 12006 26575 12008
rect 24853 12003 24919 12006
rect 26509 12003 26575 12006
rect 58157 12066 58223 12069
rect 59200 12066 60000 12096
rect 58157 12064 60000 12066
rect 58157 12008 58162 12064
rect 58218 12008 60000 12064
rect 58157 12006 60000 12008
rect 58157 12003 58223 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 59200 11976 60000 12006
rect 50290 11935 50606 11936
rect 41045 11930 41111 11933
rect 42241 11930 42307 11933
rect 41045 11928 42307 11930
rect 41045 11872 41050 11928
rect 41106 11872 42246 11928
rect 42302 11872 42307 11928
rect 41045 11870 42307 11872
rect 41045 11867 41111 11870
rect 42241 11867 42307 11870
rect 31937 11794 32003 11797
rect 40953 11794 41019 11797
rect 31937 11792 41019 11794
rect 31937 11736 31942 11792
rect 31998 11736 40958 11792
rect 41014 11736 41019 11792
rect 31937 11734 41019 11736
rect 31937 11731 32003 11734
rect 40953 11731 41019 11734
rect 41321 11794 41387 11797
rect 41505 11794 41571 11797
rect 41321 11792 41571 11794
rect 41321 11736 41326 11792
rect 41382 11736 41510 11792
rect 41566 11736 41571 11792
rect 41321 11734 41571 11736
rect 41321 11731 41387 11734
rect 41505 11731 41571 11734
rect 19517 11658 19583 11661
rect 21357 11658 21423 11661
rect 19517 11656 21423 11658
rect 19517 11600 19522 11656
rect 19578 11600 21362 11656
rect 21418 11600 21423 11656
rect 19517 11598 21423 11600
rect 19517 11595 19583 11598
rect 21357 11595 21423 11598
rect 23197 11658 23263 11661
rect 25681 11658 25747 11661
rect 38193 11658 38259 11661
rect 23197 11656 25747 11658
rect 23197 11600 23202 11656
rect 23258 11600 25686 11656
rect 25742 11600 25747 11656
rect 23197 11598 25747 11600
rect 23197 11595 23263 11598
rect 25681 11595 25747 11598
rect 31710 11656 38259 11658
rect 31710 11600 38198 11656
rect 38254 11600 38259 11656
rect 31710 11598 38259 11600
rect 0 11522 800 11552
rect 933 11522 999 11525
rect 0 11520 999 11522
rect 0 11464 938 11520
rect 994 11464 999 11520
rect 0 11462 999 11464
rect 0 11432 800 11462
rect 933 11459 999 11462
rect 19425 11522 19491 11525
rect 20110 11522 20116 11524
rect 19425 11520 20116 11522
rect 19425 11464 19430 11520
rect 19486 11464 20116 11520
rect 19425 11462 20116 11464
rect 19425 11459 19491 11462
rect 20110 11460 20116 11462
rect 20180 11460 20186 11524
rect 20345 11522 20411 11525
rect 20989 11522 21055 11525
rect 20345 11520 21055 11522
rect 20345 11464 20350 11520
rect 20406 11464 20994 11520
rect 21050 11464 21055 11520
rect 20345 11462 21055 11464
rect 20345 11459 20411 11462
rect 20989 11459 21055 11462
rect 22553 11522 22619 11525
rect 31710 11522 31770 11598
rect 38193 11595 38259 11598
rect 22553 11520 31770 11522
rect 22553 11464 22558 11520
rect 22614 11464 31770 11520
rect 22553 11462 31770 11464
rect 58985 11522 59051 11525
rect 59200 11522 60000 11552
rect 58985 11520 60000 11522
rect 58985 11464 58990 11520
rect 59046 11464 60000 11520
rect 58985 11462 60000 11464
rect 22553 11459 22619 11462
rect 58985 11459 59051 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 59200 11432 60000 11462
rect 34930 11391 35246 11392
rect 17861 11386 17927 11389
rect 30281 11386 30347 11389
rect 17861 11384 30347 11386
rect 17861 11328 17866 11384
rect 17922 11328 30286 11384
rect 30342 11328 30347 11384
rect 17861 11326 30347 11328
rect 17861 11323 17927 11326
rect 30281 11323 30347 11326
rect 15653 11250 15719 11253
rect 29453 11250 29519 11253
rect 34513 11250 34579 11253
rect 15653 11248 27538 11250
rect 15653 11192 15658 11248
rect 15714 11192 27538 11248
rect 15653 11190 27538 11192
rect 15653 11187 15719 11190
rect 17585 11114 17651 11117
rect 21633 11114 21699 11117
rect 27337 11114 27403 11117
rect 17585 11112 21699 11114
rect 17585 11056 17590 11112
rect 17646 11056 21638 11112
rect 21694 11056 21699 11112
rect 17585 11054 21699 11056
rect 17585 11051 17651 11054
rect 21633 11051 21699 11054
rect 22050 11112 27403 11114
rect 22050 11056 27342 11112
rect 27398 11056 27403 11112
rect 22050 11054 27403 11056
rect 27478 11114 27538 11190
rect 29453 11248 34579 11250
rect 29453 11192 29458 11248
rect 29514 11192 34518 11248
rect 34574 11192 34579 11248
rect 29453 11190 34579 11192
rect 29453 11187 29519 11190
rect 34513 11187 34579 11190
rect 34789 11114 34855 11117
rect 27478 11112 34855 11114
rect 27478 11056 34794 11112
rect 34850 11056 34855 11112
rect 27478 11054 34855 11056
rect 19977 10978 20043 10981
rect 20478 10978 20484 10980
rect 19977 10976 20484 10978
rect 19977 10920 19982 10976
rect 20038 10920 20484 10976
rect 19977 10918 20484 10920
rect 19977 10915 20043 10918
rect 20478 10916 20484 10918
rect 20548 10978 20554 10980
rect 22050 10978 22110 11054
rect 27337 11051 27403 11054
rect 34789 11051 34855 11054
rect 20548 10918 22110 10978
rect 38653 10980 38719 10981
rect 38653 10976 38700 10980
rect 38764 10978 38770 10980
rect 38653 10920 38658 10976
rect 20548 10916 20554 10918
rect 38653 10916 38700 10920
rect 38764 10918 38810 10978
rect 38764 10916 38770 10918
rect 38653 10915 38719 10916
rect 19570 10912 19886 10913
rect 0 10842 800 10872
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 59200 10888 60000 11008
rect 50290 10847 50606 10848
rect 933 10842 999 10845
rect 0 10840 999 10842
rect 0 10784 938 10840
rect 994 10784 999 10840
rect 0 10782 999 10784
rect 0 10752 800 10782
rect 933 10779 999 10782
rect 20345 10842 20411 10845
rect 20529 10842 20595 10845
rect 20345 10840 20595 10842
rect 20345 10784 20350 10840
rect 20406 10784 20534 10840
rect 20590 10784 20595 10840
rect 20345 10782 20595 10784
rect 20345 10779 20411 10782
rect 20529 10779 20595 10782
rect 9581 10706 9647 10709
rect 43989 10706 44055 10709
rect 9581 10704 44055 10706
rect 9581 10648 9586 10704
rect 9642 10648 43994 10704
rect 44050 10648 44055 10704
rect 9581 10646 44055 10648
rect 9581 10643 9647 10646
rect 43989 10643 44055 10646
rect 17125 10570 17191 10573
rect 27429 10570 27495 10573
rect 17125 10568 27495 10570
rect 17125 10512 17130 10568
rect 17186 10512 27434 10568
rect 27490 10512 27495 10568
rect 17125 10510 27495 10512
rect 17125 10507 17191 10510
rect 27429 10507 27495 10510
rect 28257 10570 28323 10573
rect 28809 10570 28875 10573
rect 38377 10570 38443 10573
rect 28257 10568 28875 10570
rect 28257 10512 28262 10568
rect 28318 10512 28814 10568
rect 28870 10512 28875 10568
rect 28257 10510 28875 10512
rect 28257 10507 28323 10510
rect 28809 10507 28875 10510
rect 31710 10568 38443 10570
rect 31710 10512 38382 10568
rect 38438 10512 38443 10568
rect 31710 10510 38443 10512
rect 10869 10434 10935 10437
rect 23289 10434 23355 10437
rect 10869 10432 23355 10434
rect 10869 10376 10874 10432
rect 10930 10376 23294 10432
rect 23350 10376 23355 10432
rect 10869 10374 23355 10376
rect 10869 10371 10935 10374
rect 23289 10371 23355 10374
rect 25037 10434 25103 10437
rect 26049 10434 26115 10437
rect 27153 10434 27219 10437
rect 31710 10434 31770 10510
rect 38377 10507 38443 10510
rect 25037 10432 31770 10434
rect 25037 10376 25042 10432
rect 25098 10376 26054 10432
rect 26110 10376 27158 10432
rect 27214 10376 31770 10432
rect 25037 10374 31770 10376
rect 32029 10434 32095 10437
rect 33409 10434 33475 10437
rect 34329 10434 34395 10437
rect 58157 10434 58223 10437
rect 59200 10434 60000 10464
rect 32029 10432 34714 10434
rect 32029 10376 32034 10432
rect 32090 10376 33414 10432
rect 33470 10376 34334 10432
rect 34390 10376 34714 10432
rect 32029 10374 34714 10376
rect 25037 10371 25103 10374
rect 26049 10371 26115 10374
rect 27153 10371 27219 10374
rect 32029 10371 32095 10374
rect 33409 10371 33475 10374
rect 34329 10371 34395 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 17217 10298 17283 10301
rect 27705 10298 27771 10301
rect 17217 10296 27771 10298
rect 17217 10240 17222 10296
rect 17278 10240 27710 10296
rect 27766 10240 27771 10296
rect 17217 10238 27771 10240
rect 17217 10235 17283 10238
rect 27705 10235 27771 10238
rect 0 10162 800 10192
rect 933 10162 999 10165
rect 0 10160 999 10162
rect 0 10104 938 10160
rect 994 10104 999 10160
rect 0 10102 999 10104
rect 0 10072 800 10102
rect 933 10099 999 10102
rect 17534 10100 17540 10164
rect 17604 10162 17610 10164
rect 17677 10162 17743 10165
rect 30281 10162 30347 10165
rect 17604 10160 17743 10162
rect 17604 10104 17682 10160
rect 17738 10104 17743 10160
rect 17604 10102 17743 10104
rect 17604 10100 17610 10102
rect 17677 10099 17743 10102
rect 17910 10160 30347 10162
rect 17910 10104 30286 10160
rect 30342 10104 30347 10160
rect 17910 10102 30347 10104
rect 34654 10162 34714 10374
rect 58157 10432 60000 10434
rect 58157 10376 58162 10432
rect 58218 10376 60000 10432
rect 58157 10374 60000 10376
rect 58157 10371 58223 10374
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 59200 10344 60000 10374
rect 34930 10303 35246 10304
rect 37733 10162 37799 10165
rect 34654 10160 37799 10162
rect 34654 10104 37738 10160
rect 37794 10104 37799 10160
rect 34654 10102 37799 10104
rect 13261 10026 13327 10029
rect 17910 10026 17970 10102
rect 30281 10099 30347 10102
rect 37733 10099 37799 10102
rect 38009 10162 38075 10165
rect 38285 10162 38351 10165
rect 38561 10162 38627 10165
rect 38009 10160 38351 10162
rect 38009 10104 38014 10160
rect 38070 10104 38290 10160
rect 38346 10104 38351 10160
rect 38009 10102 38351 10104
rect 38009 10099 38075 10102
rect 38285 10099 38351 10102
rect 38518 10160 38627 10162
rect 38518 10104 38566 10160
rect 38622 10104 38627 10160
rect 38518 10099 38627 10104
rect 13261 10024 17970 10026
rect 13261 9968 13266 10024
rect 13322 9968 17970 10024
rect 13261 9966 17970 9968
rect 18094 9966 31770 10026
rect 13261 9963 13327 9966
rect 15193 9890 15259 9893
rect 16389 9890 16455 9893
rect 18094 9890 18154 9966
rect 15193 9888 18154 9890
rect 15193 9832 15198 9888
rect 15254 9832 16394 9888
rect 16450 9832 18154 9888
rect 15193 9830 18154 9832
rect 20161 9890 20227 9893
rect 21725 9890 21791 9893
rect 20161 9888 21791 9890
rect 20161 9832 20166 9888
rect 20222 9832 21730 9888
rect 21786 9832 21791 9888
rect 20161 9830 21791 9832
rect 15193 9827 15259 9830
rect 16389 9827 16455 9830
rect 20161 9827 20227 9830
rect 21725 9827 21791 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 19977 9754 20043 9757
rect 20110 9754 20116 9756
rect 19977 9752 20116 9754
rect 19977 9696 19982 9752
rect 20038 9696 20116 9752
rect 19977 9694 20116 9696
rect 19977 9691 20043 9694
rect 20110 9692 20116 9694
rect 20180 9692 20186 9756
rect 21449 9754 21515 9757
rect 26049 9754 26115 9757
rect 26509 9754 26575 9757
rect 26918 9754 26924 9756
rect 21449 9752 26115 9754
rect 21449 9696 21454 9752
rect 21510 9696 26054 9752
rect 26110 9696 26115 9752
rect 21449 9694 26115 9696
rect 21449 9691 21515 9694
rect 26049 9691 26115 9694
rect 26374 9752 26924 9754
rect 26374 9696 26514 9752
rect 26570 9696 26924 9752
rect 26374 9694 26924 9696
rect 15837 9620 15903 9621
rect 15837 9618 15884 9620
rect 15796 9616 15884 9618
rect 15948 9618 15954 9620
rect 26374 9618 26434 9694
rect 26509 9691 26575 9694
rect 26918 9692 26924 9694
rect 26988 9692 26994 9756
rect 31710 9754 31770 9966
rect 38518 9893 38578 10099
rect 35249 9890 35315 9893
rect 38377 9890 38443 9893
rect 35249 9888 38443 9890
rect 35249 9832 35254 9888
rect 35310 9832 38382 9888
rect 38438 9832 38443 9888
rect 35249 9830 38443 9832
rect 38518 9888 38627 9893
rect 38518 9832 38566 9888
rect 38622 9832 38627 9888
rect 38518 9830 38627 9832
rect 35249 9827 35315 9830
rect 38377 9827 38443 9830
rect 38561 9827 38627 9830
rect 58985 9890 59051 9893
rect 59200 9890 60000 9920
rect 58985 9888 60000 9890
rect 58985 9832 58990 9888
rect 59046 9832 60000 9888
rect 58985 9830 60000 9832
rect 58985 9827 59051 9830
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 59200 9800 60000 9830
rect 50290 9759 50606 9760
rect 35893 9754 35959 9757
rect 31710 9752 35959 9754
rect 31710 9696 35898 9752
rect 35954 9696 35959 9752
rect 31710 9694 35959 9696
rect 35893 9691 35959 9694
rect 15796 9560 15842 9616
rect 15796 9558 15884 9560
rect 15837 9556 15884 9558
rect 15948 9558 26434 9618
rect 34145 9618 34211 9621
rect 38009 9618 38075 9621
rect 34145 9616 38075 9618
rect 34145 9560 34150 9616
rect 34206 9560 38014 9616
rect 38070 9560 38075 9616
rect 34145 9558 38075 9560
rect 15948 9556 15954 9558
rect 15837 9555 15903 9556
rect 34145 9555 34211 9558
rect 38009 9555 38075 9558
rect 0 9482 800 9512
rect 933 9482 999 9485
rect 0 9480 999 9482
rect 0 9424 938 9480
rect 994 9424 999 9480
rect 0 9422 999 9424
rect 0 9392 800 9422
rect 933 9419 999 9422
rect 2405 9482 2471 9485
rect 28441 9482 28507 9485
rect 2405 9480 28507 9482
rect 2405 9424 2410 9480
rect 2466 9424 28446 9480
rect 28502 9424 28507 9480
rect 2405 9422 28507 9424
rect 2405 9419 2471 9422
rect 28441 9419 28507 9422
rect 29269 9482 29335 9485
rect 30373 9482 30439 9485
rect 29269 9480 30439 9482
rect 29269 9424 29274 9480
rect 29330 9424 30378 9480
rect 30434 9424 30439 9480
rect 29269 9422 30439 9424
rect 29269 9419 29335 9422
rect 30373 9419 30439 9422
rect 37549 9482 37615 9485
rect 37917 9482 37983 9485
rect 37549 9480 37983 9482
rect 37549 9424 37554 9480
rect 37610 9424 37922 9480
rect 37978 9424 37983 9480
rect 37549 9422 37983 9424
rect 37549 9419 37615 9422
rect 37917 9419 37983 9422
rect 18229 9346 18295 9349
rect 26141 9346 26207 9349
rect 18229 9344 26207 9346
rect 18229 9288 18234 9344
rect 18290 9288 26146 9344
rect 26202 9288 26207 9344
rect 18229 9286 26207 9288
rect 18229 9283 18295 9286
rect 26141 9283 26207 9286
rect 26325 9346 26391 9349
rect 26785 9346 26851 9349
rect 27337 9346 27403 9349
rect 26325 9344 27403 9346
rect 26325 9288 26330 9344
rect 26386 9288 26790 9344
rect 26846 9288 27342 9344
rect 27398 9288 27403 9344
rect 26325 9286 27403 9288
rect 26325 9283 26391 9286
rect 26785 9283 26851 9286
rect 27337 9283 27403 9286
rect 37457 9346 37523 9349
rect 37590 9346 37596 9348
rect 37457 9344 37596 9346
rect 37457 9288 37462 9344
rect 37518 9288 37596 9344
rect 37457 9286 37596 9288
rect 37457 9283 37523 9286
rect 37590 9284 37596 9286
rect 37660 9284 37666 9348
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 59200 9256 60000 9376
rect 34930 9215 35246 9216
rect 13629 9210 13695 9213
rect 22001 9210 22067 9213
rect 25865 9210 25931 9213
rect 32121 9210 32187 9213
rect 13629 9208 20362 9210
rect 13629 9152 13634 9208
rect 13690 9152 20362 9208
rect 13629 9150 20362 9152
rect 13629 9147 13695 9150
rect 17769 9074 17835 9077
rect 20069 9074 20135 9077
rect 17769 9072 20135 9074
rect 17769 9016 17774 9072
rect 17830 9016 20074 9072
rect 20130 9016 20135 9072
rect 17769 9014 20135 9016
rect 20302 9074 20362 9150
rect 22001 9208 32187 9210
rect 22001 9152 22006 9208
rect 22062 9152 25870 9208
rect 25926 9152 32126 9208
rect 32182 9152 32187 9208
rect 22001 9150 32187 9152
rect 22001 9147 22067 9150
rect 25865 9147 25931 9150
rect 32121 9147 32187 9150
rect 35985 9210 36051 9213
rect 38285 9210 38351 9213
rect 35985 9208 38351 9210
rect 35985 9152 35990 9208
rect 36046 9152 38290 9208
rect 38346 9152 38351 9208
rect 35985 9150 38351 9152
rect 35985 9147 36051 9150
rect 38285 9147 38351 9150
rect 27613 9074 27679 9077
rect 20302 9072 27679 9074
rect 20302 9016 27618 9072
rect 27674 9016 27679 9072
rect 20302 9014 27679 9016
rect 17769 9011 17835 9014
rect 20069 9011 20135 9014
rect 27613 9011 27679 9014
rect 30097 9074 30163 9077
rect 31569 9074 31635 9077
rect 30097 9072 31635 9074
rect 30097 9016 30102 9072
rect 30158 9016 31574 9072
rect 31630 9016 31635 9072
rect 30097 9014 31635 9016
rect 30097 9011 30163 9014
rect 31569 9011 31635 9014
rect 33501 9074 33567 9077
rect 46749 9074 46815 9077
rect 33501 9072 46815 9074
rect 33501 9016 33506 9072
rect 33562 9016 46754 9072
rect 46810 9016 46815 9072
rect 33501 9014 46815 9016
rect 33501 9011 33567 9014
rect 46749 9011 46815 9014
rect 2497 8938 2563 8941
rect 23473 8938 23539 8941
rect 2497 8936 23539 8938
rect 2497 8880 2502 8936
rect 2558 8880 23478 8936
rect 23534 8880 23539 8936
rect 2497 8878 23539 8880
rect 2497 8875 2563 8878
rect 23473 8875 23539 8878
rect 25773 8938 25839 8941
rect 25998 8938 26004 8940
rect 25773 8936 26004 8938
rect 25773 8880 25778 8936
rect 25834 8880 26004 8936
rect 25773 8878 26004 8880
rect 25773 8875 25839 8878
rect 25998 8876 26004 8878
rect 26068 8876 26074 8940
rect 27654 8876 27660 8940
rect 27724 8938 27730 8940
rect 30005 8938 30071 8941
rect 27724 8936 30071 8938
rect 27724 8880 30010 8936
rect 30066 8880 30071 8936
rect 27724 8878 30071 8880
rect 27724 8876 27730 8878
rect 30005 8875 30071 8878
rect 30649 8938 30715 8941
rect 34145 8938 34211 8941
rect 30649 8936 34211 8938
rect 30649 8880 30654 8936
rect 30710 8880 34150 8936
rect 34206 8880 34211 8936
rect 30649 8878 34211 8880
rect 30649 8875 30715 8878
rect 34145 8875 34211 8878
rect 36077 8938 36143 8941
rect 40401 8938 40467 8941
rect 36077 8936 40467 8938
rect 36077 8880 36082 8936
rect 36138 8880 40406 8936
rect 40462 8880 40467 8936
rect 36077 8878 40467 8880
rect 36077 8875 36143 8878
rect 40401 8875 40467 8878
rect 0 8802 800 8832
rect 933 8802 999 8805
rect 0 8800 999 8802
rect 0 8744 938 8800
rect 994 8744 999 8800
rect 0 8742 999 8744
rect 0 8712 800 8742
rect 933 8739 999 8742
rect 20069 8802 20135 8805
rect 26785 8802 26851 8805
rect 20069 8800 26851 8802
rect 20069 8744 20074 8800
rect 20130 8744 26790 8800
rect 26846 8744 26851 8800
rect 20069 8742 26851 8744
rect 20069 8739 20135 8742
rect 26785 8739 26851 8742
rect 29177 8802 29243 8805
rect 32397 8802 32463 8805
rect 29177 8800 32463 8802
rect 29177 8744 29182 8800
rect 29238 8744 32402 8800
rect 32458 8744 32463 8800
rect 29177 8742 32463 8744
rect 29177 8739 29243 8742
rect 32397 8739 32463 8742
rect 32857 8802 32923 8805
rect 33961 8802 34027 8805
rect 38561 8802 38627 8805
rect 32857 8800 38627 8802
rect 32857 8744 32862 8800
rect 32918 8744 33966 8800
rect 34022 8744 38566 8800
rect 38622 8744 38627 8800
rect 32857 8742 38627 8744
rect 32857 8739 32923 8742
rect 33961 8739 34027 8742
rect 38561 8739 38627 8742
rect 58985 8802 59051 8805
rect 59200 8802 60000 8832
rect 58985 8800 60000 8802
rect 58985 8744 58990 8800
rect 59046 8744 60000 8800
rect 58985 8742 60000 8744
rect 58985 8739 59051 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 59200 8712 60000 8742
rect 50290 8671 50606 8672
rect 23381 8666 23447 8669
rect 26325 8666 26391 8669
rect 23381 8664 26391 8666
rect 23381 8608 23386 8664
rect 23442 8608 26330 8664
rect 26386 8608 26391 8664
rect 23381 8606 26391 8608
rect 23381 8603 23447 8606
rect 26325 8603 26391 8606
rect 29913 8666 29979 8669
rect 39113 8666 39179 8669
rect 29913 8664 39179 8666
rect 29913 8608 29918 8664
rect 29974 8608 39118 8664
rect 39174 8608 39179 8664
rect 29913 8606 39179 8608
rect 29913 8603 29979 8606
rect 39113 8603 39179 8606
rect 39297 8666 39363 8669
rect 42333 8666 42399 8669
rect 39297 8664 42399 8666
rect 39297 8608 39302 8664
rect 39358 8608 42338 8664
rect 42394 8608 42399 8664
rect 39297 8606 42399 8608
rect 39297 8603 39363 8606
rect 42333 8603 42399 8606
rect 17125 8530 17191 8533
rect 33041 8530 33107 8533
rect 17125 8528 33107 8530
rect 17125 8472 17130 8528
rect 17186 8472 33046 8528
rect 33102 8472 33107 8528
rect 17125 8470 33107 8472
rect 17125 8467 17191 8470
rect 33041 8467 33107 8470
rect 35709 8530 35775 8533
rect 52361 8530 52427 8533
rect 35709 8528 52427 8530
rect 35709 8472 35714 8528
rect 35770 8472 52366 8528
rect 52422 8472 52427 8528
rect 35709 8470 52427 8472
rect 35709 8467 35775 8470
rect 52361 8467 52427 8470
rect 22921 8394 22987 8397
rect 26509 8394 26575 8397
rect 22921 8392 26575 8394
rect 22921 8336 22926 8392
rect 22982 8336 26514 8392
rect 26570 8336 26575 8392
rect 22921 8334 26575 8336
rect 22921 8331 22987 8334
rect 26509 8331 26575 8334
rect 26877 8394 26943 8397
rect 34145 8394 34211 8397
rect 26877 8392 34211 8394
rect 26877 8336 26882 8392
rect 26938 8336 34150 8392
rect 34206 8336 34211 8392
rect 26877 8334 34211 8336
rect 26877 8331 26943 8334
rect 34145 8331 34211 8334
rect 19333 8258 19399 8261
rect 29545 8258 29611 8261
rect 19333 8256 29611 8258
rect 19333 8200 19338 8256
rect 19394 8200 29550 8256
rect 29606 8200 29611 8256
rect 19333 8198 29611 8200
rect 19333 8195 19399 8198
rect 29545 8195 29611 8198
rect 31385 8258 31451 8261
rect 31661 8258 31727 8261
rect 31385 8256 31727 8258
rect 31385 8200 31390 8256
rect 31446 8200 31666 8256
rect 31722 8200 31727 8256
rect 31385 8198 31727 8200
rect 31385 8195 31451 8198
rect 31661 8195 31727 8198
rect 58985 8258 59051 8261
rect 59200 8258 60000 8288
rect 58985 8256 60000 8258
rect 58985 8200 58990 8256
rect 59046 8200 60000 8256
rect 58985 8198 60000 8200
rect 58985 8195 59051 8198
rect 4210 8192 4526 8193
rect 0 8122 800 8152
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 59200 8168 60000 8198
rect 34930 8127 35246 8128
rect 933 8122 999 8125
rect 0 8120 999 8122
rect 0 8064 938 8120
rect 994 8064 999 8120
rect 0 8062 999 8064
rect 0 8032 800 8062
rect 933 8059 999 8062
rect 14825 8122 14891 8125
rect 17953 8122 18019 8125
rect 14825 8120 18019 8122
rect 14825 8064 14830 8120
rect 14886 8064 17958 8120
rect 18014 8064 18019 8120
rect 14825 8062 18019 8064
rect 14825 8059 14891 8062
rect 17953 8059 18019 8062
rect 24209 8122 24275 8125
rect 25589 8122 25655 8125
rect 26693 8124 26759 8125
rect 26693 8122 26740 8124
rect 24209 8120 25655 8122
rect 24209 8064 24214 8120
rect 24270 8064 25594 8120
rect 25650 8064 25655 8120
rect 24209 8062 25655 8064
rect 26648 8120 26740 8122
rect 26648 8064 26698 8120
rect 26648 8062 26740 8064
rect 24209 8059 24275 8062
rect 25589 8059 25655 8062
rect 26693 8060 26740 8062
rect 26804 8060 26810 8124
rect 39941 8122 40007 8125
rect 48221 8122 48287 8125
rect 39941 8120 48287 8122
rect 39941 8064 39946 8120
rect 40002 8064 48226 8120
rect 48282 8064 48287 8120
rect 39941 8062 48287 8064
rect 26693 8059 26759 8060
rect 39941 8059 40007 8062
rect 48221 8059 48287 8062
rect 7925 7986 7991 7989
rect 36169 7986 36235 7989
rect 36537 7986 36603 7989
rect 7925 7984 36603 7986
rect 7925 7928 7930 7984
rect 7986 7928 36174 7984
rect 36230 7928 36542 7984
rect 36598 7928 36603 7984
rect 7925 7926 36603 7928
rect 7925 7923 7991 7926
rect 36169 7923 36235 7926
rect 36537 7923 36603 7926
rect 24761 7850 24827 7853
rect 28257 7850 28323 7853
rect 24761 7848 28323 7850
rect 24761 7792 24766 7848
rect 24822 7792 28262 7848
rect 28318 7792 28323 7848
rect 24761 7790 28323 7792
rect 24761 7787 24827 7790
rect 28257 7787 28323 7790
rect 30281 7714 30347 7717
rect 33593 7714 33659 7717
rect 30281 7712 33659 7714
rect 30281 7656 30286 7712
rect 30342 7656 33598 7712
rect 33654 7656 33659 7712
rect 30281 7654 33659 7656
rect 30281 7651 30347 7654
rect 33593 7651 33659 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 59200 7624 60000 7744
rect 50290 7583 50606 7584
rect 0 7442 800 7472
rect 933 7442 999 7445
rect 0 7440 999 7442
rect 0 7384 938 7440
rect 994 7384 999 7440
rect 0 7382 999 7384
rect 0 7352 800 7382
rect 933 7379 999 7382
rect 15193 7442 15259 7445
rect 26693 7442 26759 7445
rect 15193 7440 26759 7442
rect 15193 7384 15198 7440
rect 15254 7384 26698 7440
rect 26754 7384 26759 7440
rect 15193 7382 26759 7384
rect 15193 7379 15259 7382
rect 26693 7379 26759 7382
rect 22001 7306 22067 7309
rect 28257 7306 28323 7309
rect 22001 7304 28323 7306
rect 22001 7248 22006 7304
rect 22062 7248 28262 7304
rect 28318 7248 28323 7304
rect 22001 7246 28323 7248
rect 22001 7243 22067 7246
rect 28257 7243 28323 7246
rect 27245 7170 27311 7173
rect 31201 7170 31267 7173
rect 27245 7168 31267 7170
rect 27245 7112 27250 7168
rect 27306 7112 31206 7168
rect 31262 7112 31267 7168
rect 27245 7110 31267 7112
rect 27245 7107 27311 7110
rect 31201 7107 31267 7110
rect 58893 7170 58959 7173
rect 59200 7170 60000 7200
rect 58893 7168 60000 7170
rect 58893 7112 58898 7168
rect 58954 7112 60000 7168
rect 58893 7110 60000 7112
rect 58893 7107 58959 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 59200 7080 60000 7110
rect 34930 7039 35246 7040
rect 22369 7034 22435 7037
rect 25814 7034 25820 7036
rect 22369 7032 25820 7034
rect 22369 6976 22374 7032
rect 22430 6976 25820 7032
rect 22369 6974 25820 6976
rect 22369 6971 22435 6974
rect 25814 6972 25820 6974
rect 25884 7034 25890 7036
rect 30649 7034 30715 7037
rect 25884 7032 30715 7034
rect 25884 6976 30654 7032
rect 30710 6976 30715 7032
rect 25884 6974 30715 6976
rect 25884 6972 25890 6974
rect 30649 6971 30715 6974
rect 15745 6898 15811 6901
rect 17585 6898 17651 6901
rect 26969 6900 27035 6901
rect 15745 6896 17651 6898
rect 15745 6840 15750 6896
rect 15806 6840 17590 6896
rect 17646 6840 17651 6896
rect 15745 6838 17651 6840
rect 15745 6835 15811 6838
rect 17585 6835 17651 6838
rect 26918 6836 26924 6900
rect 26988 6898 27035 6900
rect 27337 6898 27403 6901
rect 40125 6898 40191 6901
rect 26988 6896 27080 6898
rect 27030 6840 27080 6896
rect 26988 6838 27080 6840
rect 27337 6896 40191 6898
rect 27337 6840 27342 6896
rect 27398 6840 40130 6896
rect 40186 6840 40191 6896
rect 27337 6838 40191 6840
rect 26988 6836 27035 6838
rect 26969 6835 27035 6836
rect 27337 6835 27403 6838
rect 40125 6835 40191 6838
rect 0 6762 800 6792
rect 933 6762 999 6765
rect 0 6760 999 6762
rect 0 6704 938 6760
rect 994 6704 999 6760
rect 0 6702 999 6704
rect 0 6672 800 6702
rect 933 6699 999 6702
rect 1853 6762 1919 6765
rect 31201 6762 31267 6765
rect 1853 6760 31267 6762
rect 1853 6704 1858 6760
rect 1914 6704 31206 6760
rect 31262 6704 31267 6760
rect 1853 6702 31267 6704
rect 1853 6699 1919 6702
rect 31201 6699 31267 6702
rect 27797 6626 27863 6629
rect 28717 6626 28783 6629
rect 27797 6624 28783 6626
rect 27797 6568 27802 6624
rect 27858 6568 28722 6624
rect 28778 6568 28783 6624
rect 27797 6566 28783 6568
rect 27797 6563 27863 6566
rect 28717 6563 28783 6566
rect 58065 6626 58131 6629
rect 59200 6626 60000 6656
rect 58065 6624 60000 6626
rect 58065 6568 58070 6624
rect 58126 6568 60000 6624
rect 58065 6566 60000 6568
rect 58065 6563 58131 6566
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 59200 6536 60000 6566
rect 50290 6495 50606 6496
rect 15377 6354 15443 6357
rect 21214 6354 21220 6356
rect 15377 6352 21220 6354
rect 15377 6296 15382 6352
rect 15438 6296 21220 6352
rect 15377 6294 21220 6296
rect 15377 6291 15443 6294
rect 21214 6292 21220 6294
rect 21284 6354 21290 6356
rect 22185 6354 22251 6357
rect 21284 6352 22251 6354
rect 21284 6296 22190 6352
rect 22246 6296 22251 6352
rect 21284 6294 22251 6296
rect 21284 6292 21290 6294
rect 22185 6291 22251 6294
rect 15929 6218 15995 6221
rect 27654 6218 27660 6220
rect 15929 6216 27660 6218
rect 15929 6160 15934 6216
rect 15990 6160 27660 6216
rect 15929 6158 27660 6160
rect 15929 6155 15995 6158
rect 27654 6156 27660 6158
rect 27724 6156 27730 6220
rect 37181 6218 37247 6221
rect 52361 6218 52427 6221
rect 37181 6216 52427 6218
rect 37181 6160 37186 6216
rect 37242 6160 52366 6216
rect 52422 6160 52427 6216
rect 37181 6158 52427 6160
rect 37181 6155 37247 6158
rect 52361 6155 52427 6158
rect 0 6082 800 6112
rect 933 6082 999 6085
rect 0 6080 999 6082
rect 0 6024 938 6080
rect 994 6024 999 6080
rect 0 6022 999 6024
rect 0 5992 800 6022
rect 933 6019 999 6022
rect 19333 6082 19399 6085
rect 27337 6082 27403 6085
rect 19333 6080 27403 6082
rect 19333 6024 19338 6080
rect 19394 6024 27342 6080
rect 27398 6024 27403 6080
rect 19333 6022 27403 6024
rect 19333 6019 19399 6022
rect 27337 6019 27403 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 59200 5992 60000 6112
rect 34930 5951 35246 5952
rect 27705 5810 27771 5813
rect 29494 5810 29500 5812
rect 27705 5808 29500 5810
rect 27705 5752 27710 5808
rect 27766 5752 29500 5808
rect 27705 5750 29500 5752
rect 27705 5747 27771 5750
rect 29494 5748 29500 5750
rect 29564 5810 29570 5812
rect 38377 5810 38443 5813
rect 29564 5808 38443 5810
rect 29564 5752 38382 5808
rect 38438 5752 38443 5808
rect 29564 5750 38443 5752
rect 29564 5748 29570 5750
rect 38377 5747 38443 5750
rect 29637 5674 29703 5677
rect 33317 5674 33383 5677
rect 29637 5672 33383 5674
rect 29637 5616 29642 5672
rect 29698 5616 33322 5672
rect 33378 5616 33383 5672
rect 29637 5614 33383 5616
rect 29637 5611 29703 5614
rect 33317 5611 33383 5614
rect 22369 5540 22435 5541
rect 22318 5538 22324 5540
rect 22278 5478 22324 5538
rect 22388 5536 22435 5540
rect 22430 5480 22435 5536
rect 22318 5476 22324 5478
rect 22388 5476 22435 5480
rect 42558 5476 42564 5540
rect 42628 5538 42634 5540
rect 42701 5538 42767 5541
rect 42628 5536 42767 5538
rect 42628 5480 42706 5536
rect 42762 5480 42767 5536
rect 42628 5478 42767 5480
rect 42628 5476 42634 5478
rect 22369 5475 22435 5476
rect 42701 5475 42767 5478
rect 58985 5538 59051 5541
rect 59200 5538 60000 5568
rect 58985 5536 60000 5538
rect 58985 5480 58990 5536
rect 59046 5480 60000 5536
rect 58985 5478 60000 5480
rect 58985 5475 59051 5478
rect 19570 5472 19886 5473
rect 0 5402 800 5432
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 59200 5448 60000 5478
rect 50290 5407 50606 5408
rect 933 5402 999 5405
rect 28993 5402 29059 5405
rect 0 5400 999 5402
rect 0 5344 938 5400
rect 994 5344 999 5400
rect 0 5342 999 5344
rect 0 5312 800 5342
rect 933 5339 999 5342
rect 22050 5400 29059 5402
rect 22050 5344 28998 5400
rect 29054 5344 29059 5400
rect 22050 5342 29059 5344
rect 14917 5266 14983 5269
rect 22050 5266 22110 5342
rect 28993 5339 29059 5342
rect 41689 5402 41755 5405
rect 45921 5402 45987 5405
rect 41689 5400 45987 5402
rect 41689 5344 41694 5400
rect 41750 5344 45926 5400
rect 45982 5344 45987 5400
rect 41689 5342 45987 5344
rect 41689 5339 41755 5342
rect 45921 5339 45987 5342
rect 14917 5264 22110 5266
rect 14917 5208 14922 5264
rect 14978 5208 22110 5264
rect 14917 5206 22110 5208
rect 25221 5266 25287 5269
rect 35157 5266 35223 5269
rect 36169 5266 36235 5269
rect 25221 5264 31770 5266
rect 25221 5208 25226 5264
rect 25282 5208 31770 5264
rect 25221 5206 31770 5208
rect 14917 5203 14983 5206
rect 25221 5203 25287 5206
rect 18505 5130 18571 5133
rect 31710 5130 31770 5206
rect 35157 5264 36235 5266
rect 35157 5208 35162 5264
rect 35218 5208 36174 5264
rect 36230 5208 36235 5264
rect 35157 5206 36235 5208
rect 35157 5203 35223 5206
rect 36169 5203 36235 5206
rect 42517 5130 42583 5133
rect 18505 5128 26986 5130
rect 18505 5072 18510 5128
rect 18566 5072 26986 5128
rect 18505 5070 26986 5072
rect 31710 5128 42583 5130
rect 31710 5072 42522 5128
rect 42578 5072 42583 5128
rect 31710 5070 42583 5072
rect 18505 5067 18571 5070
rect 5257 4994 5323 4997
rect 23381 4994 23447 4997
rect 5257 4992 23447 4994
rect 5257 4936 5262 4992
rect 5318 4936 23386 4992
rect 23442 4936 23447 4992
rect 5257 4934 23447 4936
rect 26926 4994 26986 5070
rect 42517 5067 42583 5070
rect 32949 4994 33015 4997
rect 26926 4992 33015 4994
rect 26926 4936 32954 4992
rect 33010 4936 33015 4992
rect 26926 4934 33015 4936
rect 5257 4931 5323 4934
rect 23381 4931 23447 4934
rect 32949 4931 33015 4934
rect 58065 4994 58131 4997
rect 59200 4994 60000 5024
rect 58065 4992 60000 4994
rect 58065 4936 58070 4992
rect 58126 4936 60000 4992
rect 58065 4934 60000 4936
rect 58065 4931 58131 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 59200 4904 60000 4934
rect 34930 4863 35246 4864
rect 15285 4858 15351 4861
rect 21633 4858 21699 4861
rect 15285 4856 21699 4858
rect 15285 4800 15290 4856
rect 15346 4800 21638 4856
rect 21694 4800 21699 4856
rect 15285 4798 21699 4800
rect 15285 4795 15351 4798
rect 21633 4795 21699 4798
rect 22737 4858 22803 4861
rect 30741 4858 30807 4861
rect 22737 4856 30807 4858
rect 22737 4800 22742 4856
rect 22798 4800 30746 4856
rect 30802 4800 30807 4856
rect 22737 4798 30807 4800
rect 22737 4795 22803 4798
rect 30741 4795 30807 4798
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 9765 4722 9831 4725
rect 14825 4722 14891 4725
rect 9765 4720 14891 4722
rect 9765 4664 9770 4720
rect 9826 4664 14830 4720
rect 14886 4664 14891 4720
rect 9765 4662 14891 4664
rect 9765 4659 9831 4662
rect 14825 4659 14891 4662
rect 17953 4722 18019 4725
rect 23657 4722 23723 4725
rect 17953 4720 23723 4722
rect 17953 4664 17958 4720
rect 18014 4664 23662 4720
rect 23718 4664 23723 4720
rect 17953 4662 23723 4664
rect 17953 4659 18019 4662
rect 23657 4659 23723 4662
rect 28993 4722 29059 4725
rect 36353 4722 36419 4725
rect 28993 4720 36419 4722
rect 28993 4664 28998 4720
rect 29054 4664 36358 4720
rect 36414 4664 36419 4720
rect 28993 4662 36419 4664
rect 28993 4659 29059 4662
rect 36353 4659 36419 4662
rect 14733 4586 14799 4589
rect 31477 4586 31543 4589
rect 14733 4584 31543 4586
rect 14733 4528 14738 4584
rect 14794 4528 31482 4584
rect 31538 4528 31543 4584
rect 14733 4526 31543 4528
rect 14733 4523 14799 4526
rect 31477 4523 31543 4526
rect 20437 4450 20503 4453
rect 28717 4450 28783 4453
rect 20437 4448 28783 4450
rect 20437 4392 20442 4448
rect 20498 4392 28722 4448
rect 28778 4392 28783 4448
rect 20437 4390 28783 4392
rect 20437 4387 20503 4390
rect 28717 4387 28783 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 59200 4360 60000 4480
rect 50290 4319 50606 4320
rect 22553 4178 22619 4181
rect 28257 4178 28323 4181
rect 33041 4178 33107 4181
rect 22553 4176 33107 4178
rect 22553 4120 22558 4176
rect 22614 4120 28262 4176
rect 28318 4120 33046 4176
rect 33102 4120 33107 4176
rect 22553 4118 33107 4120
rect 22553 4115 22619 4118
rect 28257 4115 28323 4118
rect 33041 4115 33107 4118
rect 34697 4178 34763 4181
rect 36445 4178 36511 4181
rect 38193 4178 38259 4181
rect 34697 4176 34898 4178
rect 34697 4120 34702 4176
rect 34758 4120 34898 4176
rect 34697 4118 34898 4120
rect 34697 4115 34763 4118
rect 0 4042 800 4072
rect 933 4042 999 4045
rect 0 4040 999 4042
rect 0 3984 938 4040
rect 994 3984 999 4040
rect 0 3982 999 3984
rect 0 3952 800 3982
rect 933 3979 999 3982
rect 5717 4042 5783 4045
rect 8937 4042 9003 4045
rect 5717 4040 9003 4042
rect 5717 3984 5722 4040
rect 5778 3984 8942 4040
rect 8998 3984 9003 4040
rect 5717 3982 9003 3984
rect 5717 3979 5783 3982
rect 8937 3979 9003 3982
rect 12893 4042 12959 4045
rect 22645 4044 22711 4045
rect 12893 4040 22110 4042
rect 12893 3984 12898 4040
rect 12954 3984 22110 4040
rect 12893 3982 22110 3984
rect 12893 3979 12959 3982
rect 22050 3906 22110 3982
rect 22645 4040 22692 4044
rect 22756 4042 22762 4044
rect 25773 4042 25839 4045
rect 27286 4042 27292 4044
rect 22645 3984 22650 4040
rect 22645 3980 22692 3984
rect 22756 3982 22802 4042
rect 25773 4040 27292 4042
rect 25773 3984 25778 4040
rect 25834 3984 27292 4040
rect 25773 3982 27292 3984
rect 22756 3980 22762 3982
rect 22645 3979 22711 3980
rect 25773 3979 25839 3982
rect 27286 3980 27292 3982
rect 27356 3980 27362 4044
rect 34838 4042 34898 4118
rect 36445 4176 38259 4178
rect 36445 4120 36450 4176
rect 36506 4120 38198 4176
rect 38254 4120 38259 4176
rect 36445 4118 38259 4120
rect 36445 4115 36511 4118
rect 38193 4115 38259 4118
rect 35893 4044 35959 4045
rect 34838 3982 35450 4042
rect 31477 3906 31543 3909
rect 22050 3904 31543 3906
rect 22050 3848 31482 3904
rect 31538 3848 31543 3904
rect 22050 3846 31543 3848
rect 35390 3906 35450 3982
rect 35893 4040 35940 4044
rect 36004 4042 36010 4044
rect 37089 4042 37155 4045
rect 38193 4042 38259 4045
rect 35893 3984 35898 4040
rect 35893 3980 35940 3984
rect 36004 3982 36050 4042
rect 37089 4040 38259 4042
rect 37089 3984 37094 4040
rect 37150 3984 38198 4040
rect 38254 3984 38259 4040
rect 37089 3982 38259 3984
rect 36004 3980 36010 3982
rect 35893 3979 35959 3980
rect 37089 3979 37155 3982
rect 38193 3979 38259 3982
rect 41781 4044 41847 4045
rect 41781 4040 41828 4044
rect 41892 4042 41898 4044
rect 41781 3984 41786 4040
rect 41781 3980 41828 3984
rect 41892 3982 41938 4042
rect 41892 3980 41898 3982
rect 41781 3979 41847 3980
rect 41321 3906 41387 3909
rect 55305 3906 55371 3909
rect 35390 3904 41387 3906
rect 35390 3848 41326 3904
rect 41382 3848 41387 3904
rect 35390 3846 41387 3848
rect 31477 3843 31543 3846
rect 41321 3843 41387 3846
rect 51030 3904 55371 3906
rect 51030 3848 55310 3904
rect 55366 3848 55371 3904
rect 51030 3846 55371 3848
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 15193 3770 15259 3773
rect 31753 3770 31819 3773
rect 15193 3768 31819 3770
rect 15193 3712 15198 3768
rect 15254 3712 31758 3768
rect 31814 3712 31819 3768
rect 15193 3710 31819 3712
rect 15193 3707 15259 3710
rect 31753 3707 31819 3710
rect 37825 3770 37891 3773
rect 38285 3770 38351 3773
rect 51030 3770 51090 3846
rect 55305 3843 55371 3846
rect 58985 3906 59051 3909
rect 59200 3906 60000 3936
rect 58985 3904 60000 3906
rect 58985 3848 58990 3904
rect 59046 3848 60000 3904
rect 58985 3846 60000 3848
rect 58985 3843 59051 3846
rect 59200 3816 60000 3846
rect 37825 3768 38351 3770
rect 37825 3712 37830 3768
rect 37886 3712 38290 3768
rect 38346 3712 38351 3768
rect 37825 3710 38351 3712
rect 37825 3707 37891 3710
rect 38285 3707 38351 3710
rect 38610 3710 51090 3770
rect 12617 3634 12683 3637
rect 12985 3634 13051 3637
rect 12617 3632 13051 3634
rect 12617 3576 12622 3632
rect 12678 3576 12990 3632
rect 13046 3576 13051 3632
rect 12617 3574 13051 3576
rect 12617 3571 12683 3574
rect 12985 3571 13051 3574
rect 19701 3634 19767 3637
rect 22645 3634 22711 3637
rect 19701 3632 22711 3634
rect 19701 3576 19706 3632
rect 19762 3576 22650 3632
rect 22706 3576 22711 3632
rect 19701 3574 22711 3576
rect 19701 3571 19767 3574
rect 22645 3571 22711 3574
rect 15837 3498 15903 3501
rect 23657 3498 23723 3501
rect 15837 3496 23723 3498
rect 15837 3440 15842 3496
rect 15898 3440 23662 3496
rect 23718 3440 23723 3496
rect 15837 3438 23723 3440
rect 15837 3435 15903 3438
rect 23657 3435 23723 3438
rect 0 3362 800 3392
rect 933 3362 999 3365
rect 0 3360 999 3362
rect 0 3304 938 3360
rect 994 3304 999 3360
rect 0 3302 999 3304
rect 0 3272 800 3302
rect 933 3299 999 3302
rect 20529 3362 20595 3365
rect 37733 3362 37799 3365
rect 38610 3362 38670 3710
rect 39982 3572 39988 3636
rect 40052 3634 40058 3636
rect 40401 3634 40467 3637
rect 40052 3632 40467 3634
rect 40052 3576 40406 3632
rect 40462 3576 40467 3632
rect 40052 3574 40467 3576
rect 40052 3572 40058 3574
rect 40401 3571 40467 3574
rect 43713 3634 43779 3637
rect 43846 3634 43852 3636
rect 43713 3632 43852 3634
rect 43713 3576 43718 3632
rect 43774 3576 43852 3632
rect 43713 3574 43852 3576
rect 43713 3571 43779 3574
rect 43846 3572 43852 3574
rect 43916 3572 43922 3636
rect 20529 3360 38670 3362
rect 20529 3304 20534 3360
rect 20590 3304 37738 3360
rect 37794 3304 38670 3360
rect 20529 3302 38670 3304
rect 58157 3362 58223 3365
rect 59200 3362 60000 3392
rect 58157 3360 60000 3362
rect 58157 3304 58162 3360
rect 58218 3304 60000 3360
rect 58157 3302 60000 3304
rect 20529 3299 20595 3302
rect 37733 3299 37799 3302
rect 58157 3299 58223 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 59200 3272 60000 3302
rect 50290 3231 50606 3232
rect 6913 3226 6979 3229
rect 19333 3226 19399 3229
rect 6913 3224 19399 3226
rect 6913 3168 6918 3224
rect 6974 3168 19338 3224
rect 19394 3168 19399 3224
rect 6913 3166 19399 3168
rect 6913 3163 6979 3166
rect 19333 3163 19399 3166
rect 23657 3226 23723 3229
rect 31017 3226 31083 3229
rect 23657 3224 31083 3226
rect 23657 3168 23662 3224
rect 23718 3168 31022 3224
rect 31078 3168 31083 3224
rect 23657 3166 31083 3168
rect 23657 3163 23723 3166
rect 31017 3163 31083 3166
rect 31150 3164 31156 3228
rect 31220 3226 31226 3228
rect 42609 3226 42675 3229
rect 31220 3224 42675 3226
rect 31220 3168 42614 3224
rect 42670 3168 42675 3224
rect 31220 3166 42675 3168
rect 31220 3164 31226 3166
rect 42609 3163 42675 3166
rect 5809 3090 5875 3093
rect 9305 3090 9371 3093
rect 5809 3088 9371 3090
rect 5809 3032 5814 3088
rect 5870 3032 9310 3088
rect 9366 3032 9371 3088
rect 5809 3030 9371 3032
rect 5809 3027 5875 3030
rect 9305 3027 9371 3030
rect 9489 3090 9555 3093
rect 27521 3090 27587 3093
rect 9489 3088 27587 3090
rect 9489 3032 9494 3088
rect 9550 3032 27526 3088
rect 27582 3032 27587 3088
rect 9489 3030 27587 3032
rect 9489 3027 9555 3030
rect 27521 3027 27587 3030
rect 29126 3028 29132 3092
rect 29196 3090 29202 3092
rect 42609 3090 42675 3093
rect 29196 3088 42675 3090
rect 29196 3032 42614 3088
rect 42670 3032 42675 3088
rect 29196 3030 42675 3032
rect 29196 3028 29202 3030
rect 42609 3027 42675 3030
rect 5993 2954 6059 2957
rect 14825 2954 14891 2957
rect 20713 2954 20779 2957
rect 5993 2952 12450 2954
rect 5993 2896 5998 2952
rect 6054 2896 12450 2952
rect 5993 2894 12450 2896
rect 5993 2891 6059 2894
rect 7649 2818 7715 2821
rect 10317 2818 10383 2821
rect 7649 2816 10383 2818
rect 7649 2760 7654 2816
rect 7710 2760 10322 2816
rect 10378 2760 10383 2816
rect 7649 2758 10383 2760
rect 12390 2818 12450 2894
rect 14825 2952 20779 2954
rect 14825 2896 14830 2952
rect 14886 2896 20718 2952
rect 20774 2896 20779 2952
rect 14825 2894 20779 2896
rect 14825 2891 14891 2894
rect 20713 2891 20779 2894
rect 24117 2818 24183 2821
rect 12390 2816 24183 2818
rect 12390 2760 24122 2816
rect 24178 2760 24183 2816
rect 12390 2758 24183 2760
rect 7649 2755 7715 2758
rect 10317 2755 10383 2758
rect 24117 2755 24183 2758
rect 58985 2818 59051 2821
rect 59200 2818 60000 2848
rect 58985 2816 60000 2818
rect 58985 2760 58990 2816
rect 59046 2760 60000 2816
rect 58985 2758 60000 2760
rect 58985 2755 59051 2758
rect 4210 2752 4526 2753
rect 0 2682 800 2712
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 59200 2728 60000 2758
rect 34930 2687 35246 2688
rect 933 2682 999 2685
rect 0 2680 999 2682
rect 0 2624 938 2680
rect 994 2624 999 2680
rect 0 2622 999 2624
rect 0 2592 800 2622
rect 933 2619 999 2622
rect 27102 2484 27108 2548
rect 27172 2546 27178 2548
rect 44173 2546 44239 2549
rect 27172 2544 44239 2546
rect 27172 2488 44178 2544
rect 44234 2488 44239 2544
rect 27172 2486 44239 2488
rect 27172 2484 27178 2486
rect 44173 2483 44239 2486
rect 25998 2348 26004 2412
rect 26068 2410 26074 2412
rect 52453 2410 52519 2413
rect 26068 2408 52519 2410
rect 26068 2352 52458 2408
rect 52514 2352 52519 2408
rect 26068 2350 52519 2352
rect 26068 2348 26074 2350
rect 52453 2347 52519 2350
rect 58893 2274 58959 2277
rect 59200 2274 60000 2304
rect 58893 2272 60000 2274
rect 58893 2216 58898 2272
rect 58954 2216 60000 2272
rect 58893 2214 60000 2216
rect 58893 2211 58959 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 59200 2184 60000 2214
rect 50290 2143 50606 2144
rect 0 2002 800 2032
rect 933 2002 999 2005
rect 0 2000 999 2002
rect 0 1944 938 2000
rect 994 1944 999 2000
rect 0 1942 999 1944
rect 0 1912 800 1942
rect 933 1939 999 1942
rect 58801 1730 58867 1733
rect 59200 1730 60000 1760
rect 58801 1728 60000 1730
rect 58801 1672 58806 1728
rect 58862 1672 60000 1728
rect 58801 1670 60000 1672
rect 58801 1667 58867 1670
rect 59200 1640 60000 1670
rect 56501 1186 56567 1189
rect 59200 1186 60000 1216
rect 56501 1184 60000 1186
rect 56501 1128 56506 1184
rect 56562 1128 60000 1184
rect 56501 1126 60000 1128
rect 56501 1123 56567 1126
rect 59200 1096 60000 1126
<< via3 >>
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 19576 60956 19640 60960
rect 19576 60900 19580 60956
rect 19580 60900 19636 60956
rect 19636 60900 19640 60956
rect 19576 60896 19640 60900
rect 19656 60956 19720 60960
rect 19656 60900 19660 60956
rect 19660 60900 19716 60956
rect 19716 60900 19720 60956
rect 19656 60896 19720 60900
rect 19736 60956 19800 60960
rect 19736 60900 19740 60956
rect 19740 60900 19796 60956
rect 19796 60900 19800 60956
rect 19736 60896 19800 60900
rect 19816 60956 19880 60960
rect 19816 60900 19820 60956
rect 19820 60900 19876 60956
rect 19876 60900 19880 60956
rect 19816 60896 19880 60900
rect 50296 60956 50360 60960
rect 50296 60900 50300 60956
rect 50300 60900 50356 60956
rect 50356 60900 50360 60956
rect 50296 60896 50360 60900
rect 50376 60956 50440 60960
rect 50376 60900 50380 60956
rect 50380 60900 50436 60956
rect 50436 60900 50440 60956
rect 50376 60896 50440 60900
rect 50456 60956 50520 60960
rect 50456 60900 50460 60956
rect 50460 60900 50516 60956
rect 50516 60900 50520 60956
rect 50456 60896 50520 60900
rect 50536 60956 50600 60960
rect 50536 60900 50540 60956
rect 50540 60900 50596 60956
rect 50596 60900 50600 60956
rect 50536 60896 50600 60900
rect 20484 60692 20548 60756
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 31156 60072 31220 60076
rect 31156 60016 31170 60072
rect 31170 60016 31220 60072
rect 31156 60012 31220 60016
rect 29132 59936 29196 59940
rect 29132 59880 29146 59936
rect 29146 59880 29196 59936
rect 29132 59876 29196 59880
rect 32444 59876 32508 59940
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 21956 59332 22020 59396
rect 42564 59332 42628 59396
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 43852 56612 43916 56676
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 25268 55252 25332 55316
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 25084 52532 25148 52596
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 35940 50220 36004 50284
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 38700 47500 38764 47564
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 37596 44780 37660 44844
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 15884 44236 15948 44300
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 26740 42740 26804 42804
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 39252 38796 39316 38860
rect 22508 38720 22572 38724
rect 22508 38664 22522 38720
rect 22522 38664 22572 38720
rect 22508 38660 22572 38664
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 23428 37708 23492 37772
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 16804 35124 16868 35188
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 17540 34580 17604 34644
rect 24716 34580 24780 34644
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 21220 33356 21284 33420
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 23428 31180 23492 31244
rect 41828 31180 41892 31244
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 21956 29820 22020 29884
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 40540 24108 40604 24172
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 22324 19756 22388 19820
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 27292 18124 27356 18188
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 22692 17852 22756 17916
rect 26188 17852 26252 17916
rect 27108 17640 27172 17644
rect 27108 17584 27122 17640
rect 27122 17584 27172 17640
rect 27108 17580 27172 17584
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 22876 16688 22940 16692
rect 22876 16632 22890 16688
rect 22890 16632 22940 16688
rect 22876 16628 22940 16632
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 25268 15192 25332 15196
rect 25268 15136 25282 15192
rect 25282 15136 25332 15192
rect 25268 15132 25332 15136
rect 25820 15056 25884 15060
rect 25820 15000 25834 15056
rect 25834 15000 25884 15056
rect 25820 14996 25884 15000
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 25084 14452 25148 14516
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 26188 14104 26252 14108
rect 26188 14048 26202 14104
rect 26202 14048 26252 14104
rect 26188 14044 26252 14048
rect 22508 13636 22572 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 32444 13500 32508 13564
rect 29500 13092 29564 13156
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 22876 12684 22940 12748
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 16804 12276 16868 12340
rect 24716 12276 24780 12340
rect 40540 12276 40604 12340
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 20116 11460 20180 11524
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 20484 10916 20548 10980
rect 38700 10976 38764 10980
rect 38700 10920 38714 10976
rect 38714 10920 38764 10976
rect 38700 10916 38764 10920
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 17540 10100 17604 10164
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 20116 9692 20180 9756
rect 15884 9616 15948 9620
rect 26924 9692 26988 9756
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 15884 9560 15898 9616
rect 15898 9560 15948 9616
rect 15884 9556 15948 9560
rect 37596 9284 37660 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 26004 8876 26068 8940
rect 27660 8876 27724 8940
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 26740 8120 26804 8124
rect 26740 8064 26754 8120
rect 26754 8064 26804 8120
rect 26740 8060 26804 8064
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 25820 6972 25884 7036
rect 26924 6896 26988 6900
rect 26924 6840 26974 6896
rect 26974 6840 26988 6896
rect 26924 6836 26988 6840
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 21220 6292 21284 6356
rect 27660 6156 27724 6220
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 29500 5748 29564 5812
rect 22324 5536 22388 5540
rect 22324 5480 22374 5536
rect 22374 5480 22388 5536
rect 22324 5476 22388 5480
rect 42564 5476 42628 5540
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 22692 4040 22756 4044
rect 22692 3984 22706 4040
rect 22706 3984 22756 4040
rect 22692 3980 22756 3984
rect 27292 3980 27356 4044
rect 35940 4040 36004 4044
rect 35940 3984 35954 4040
rect 35954 3984 36004 4040
rect 35940 3980 36004 3984
rect 41828 4040 41892 4044
rect 41828 3984 41842 4040
rect 41842 3984 41892 4040
rect 41828 3980 41892 3984
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 39988 3572 40052 3636
rect 43852 3572 43916 3636
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 31156 3164 31220 3228
rect 29132 3028 29196 3092
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 27108 2484 27172 2548
rect 26004 2348 26068 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 61504 4528 61520
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 19568 60960 19888 61520
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 59872 19888 60896
rect 34928 61504 35248 61520
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 20483 60756 20549 60757
rect 20483 60692 20484 60756
rect 20548 60692 20549 60756
rect 20483 60691 20549 60692
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 58784 19888 59808
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 15883 44300 15949 44301
rect 15883 44236 15884 44300
rect 15948 44236 15949 44300
rect 15883 44235 15949 44236
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 15886 9621 15946 44235
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 16803 35188 16869 35189
rect 16803 35124 16804 35188
rect 16868 35124 16869 35188
rect 16803 35123 16869 35124
rect 16806 12341 16866 35123
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 17539 34644 17605 34645
rect 17539 34580 17540 34644
rect 17604 34580 17605 34644
rect 17539 34579 17605 34580
rect 16803 12340 16869 12341
rect 16803 12276 16804 12340
rect 16868 12276 16869 12340
rect 16803 12275 16869 12276
rect 17542 10165 17602 34579
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 20115 11524 20181 11525
rect 20115 11460 20116 11524
rect 20180 11460 20181 11524
rect 20115 11459 20181 11460
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 17539 10164 17605 10165
rect 17539 10100 17540 10164
rect 17604 10100 17605 10164
rect 17539 10099 17605 10100
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 15883 9620 15949 9621
rect 15883 9556 15884 9620
rect 15948 9556 15949 9620
rect 15883 9555 15949 9556
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 8736 19888 9760
rect 20118 9757 20178 11459
rect 20486 10981 20546 60691
rect 34928 60416 35248 61440
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 31155 60076 31221 60077
rect 31155 60012 31156 60076
rect 31220 60012 31221 60076
rect 31155 60011 31221 60012
rect 29131 59940 29197 59941
rect 29131 59876 29132 59940
rect 29196 59876 29197 59940
rect 29131 59875 29197 59876
rect 21955 59396 22021 59397
rect 21955 59332 21956 59396
rect 22020 59332 22021 59396
rect 21955 59331 22021 59332
rect 21219 33420 21285 33421
rect 21219 33356 21220 33420
rect 21284 33356 21285 33420
rect 21219 33355 21285 33356
rect 20483 10980 20549 10981
rect 20483 10916 20484 10980
rect 20548 10916 20549 10980
rect 20483 10915 20549 10916
rect 20115 9756 20181 9757
rect 20115 9692 20116 9756
rect 20180 9692 20181 9756
rect 20115 9691 20181 9692
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 21222 6357 21282 33355
rect 21958 29885 22018 59331
rect 25267 55316 25333 55317
rect 25267 55252 25268 55316
rect 25332 55252 25333 55316
rect 25267 55251 25333 55252
rect 25083 52596 25149 52597
rect 25083 52532 25084 52596
rect 25148 52532 25149 52596
rect 25083 52531 25149 52532
rect 22507 38724 22573 38725
rect 22507 38660 22508 38724
rect 22572 38660 22573 38724
rect 22507 38659 22573 38660
rect 21955 29884 22021 29885
rect 21955 29820 21956 29884
rect 22020 29820 22021 29884
rect 21955 29819 22021 29820
rect 22323 19820 22389 19821
rect 22323 19756 22324 19820
rect 22388 19756 22389 19820
rect 22323 19755 22389 19756
rect 21219 6356 21285 6357
rect 21219 6292 21220 6356
rect 21284 6292 21285 6356
rect 21219 6291 21285 6292
rect 22326 5541 22386 19755
rect 22510 13701 22570 38659
rect 23427 37772 23493 37773
rect 23427 37708 23428 37772
rect 23492 37708 23493 37772
rect 23427 37707 23493 37708
rect 23430 31245 23490 37707
rect 24715 34644 24781 34645
rect 24715 34580 24716 34644
rect 24780 34580 24781 34644
rect 24715 34579 24781 34580
rect 23427 31244 23493 31245
rect 23427 31180 23428 31244
rect 23492 31180 23493 31244
rect 23427 31179 23493 31180
rect 22691 17916 22757 17917
rect 22691 17852 22692 17916
rect 22756 17852 22757 17916
rect 22691 17851 22757 17852
rect 22507 13700 22573 13701
rect 22507 13636 22508 13700
rect 22572 13636 22573 13700
rect 22507 13635 22573 13636
rect 22323 5540 22389 5541
rect 22323 5476 22324 5540
rect 22388 5476 22389 5540
rect 22323 5475 22389 5476
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 22694 4045 22754 17851
rect 22875 16692 22941 16693
rect 22875 16628 22876 16692
rect 22940 16628 22941 16692
rect 22875 16627 22941 16628
rect 22878 12749 22938 16627
rect 22875 12748 22941 12749
rect 22875 12684 22876 12748
rect 22940 12684 22941 12748
rect 22875 12683 22941 12684
rect 24718 12341 24778 34579
rect 25086 14517 25146 52531
rect 25270 15197 25330 55251
rect 26739 42804 26805 42805
rect 26739 42740 26740 42804
rect 26804 42740 26805 42804
rect 26739 42739 26805 42740
rect 26187 17916 26253 17917
rect 26187 17852 26188 17916
rect 26252 17852 26253 17916
rect 26187 17851 26253 17852
rect 25267 15196 25333 15197
rect 25267 15132 25268 15196
rect 25332 15132 25333 15196
rect 25267 15131 25333 15132
rect 25819 15060 25885 15061
rect 25819 14996 25820 15060
rect 25884 14996 25885 15060
rect 25819 14995 25885 14996
rect 25083 14516 25149 14517
rect 25083 14452 25084 14516
rect 25148 14452 25149 14516
rect 25083 14451 25149 14452
rect 24715 12340 24781 12341
rect 24715 12276 24716 12340
rect 24780 12276 24781 12340
rect 24715 12275 24781 12276
rect 25822 7037 25882 14995
rect 26190 14109 26250 17851
rect 26187 14108 26253 14109
rect 26187 14044 26188 14108
rect 26252 14044 26253 14108
rect 26187 14043 26253 14044
rect 26003 8940 26069 8941
rect 26003 8876 26004 8940
rect 26068 8876 26069 8940
rect 26003 8875 26069 8876
rect 25819 7036 25885 7037
rect 25819 6972 25820 7036
rect 25884 6972 25885 7036
rect 25819 6971 25885 6972
rect 22691 4044 22757 4045
rect 22691 3980 22692 4044
rect 22756 3980 22757 4044
rect 22691 3979 22757 3980
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 26006 2413 26066 8875
rect 26742 8125 26802 42739
rect 27291 18188 27357 18189
rect 27291 18124 27292 18188
rect 27356 18124 27357 18188
rect 27291 18123 27357 18124
rect 27107 17644 27173 17645
rect 27107 17580 27108 17644
rect 27172 17580 27173 17644
rect 27107 17579 27173 17580
rect 26923 9756 26989 9757
rect 26923 9692 26924 9756
rect 26988 9692 26989 9756
rect 26923 9691 26989 9692
rect 26739 8124 26805 8125
rect 26739 8060 26740 8124
rect 26804 8060 26805 8124
rect 26739 8059 26805 8060
rect 26926 6901 26986 9691
rect 26923 6900 26989 6901
rect 26923 6836 26924 6900
rect 26988 6836 26989 6900
rect 26923 6835 26989 6836
rect 27110 2549 27170 17579
rect 27294 4045 27354 18123
rect 27659 8940 27725 8941
rect 27659 8876 27660 8940
rect 27724 8876 27725 8940
rect 27659 8875 27725 8876
rect 27662 6221 27722 8875
rect 27659 6220 27725 6221
rect 27659 6156 27660 6220
rect 27724 6156 27725 6220
rect 27659 6155 27725 6156
rect 27291 4044 27357 4045
rect 27291 3980 27292 4044
rect 27356 3980 27357 4044
rect 27291 3979 27357 3980
rect 29134 3093 29194 59875
rect 29499 13156 29565 13157
rect 29499 13092 29500 13156
rect 29564 13092 29565 13156
rect 29499 13091 29565 13092
rect 29502 5813 29562 13091
rect 29499 5812 29565 5813
rect 29499 5748 29500 5812
rect 29564 5748 29565 5812
rect 29499 5747 29565 5748
rect 31158 3229 31218 60011
rect 32443 59940 32509 59941
rect 32443 59876 32444 59940
rect 32508 59876 32509 59940
rect 32443 59875 32509 59876
rect 32446 13565 32506 59875
rect 34928 59328 35248 60352
rect 50288 60960 50608 61520
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 59872 50608 60896
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 42563 59396 42629 59397
rect 42563 59332 42564 59396
rect 42628 59332 42629 59396
rect 42563 59331 42629 59332
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 57152 35248 58176
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 35939 50284 36005 50285
rect 35939 50220 35940 50284
rect 36004 50220 36005 50284
rect 35939 50219 36005 50220
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 32443 13564 32509 13565
rect 32443 13500 32444 13564
rect 32508 13500 32509 13564
rect 32443 13499 32509 13500
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 35942 4045 36002 50219
rect 38699 47564 38765 47565
rect 38699 47500 38700 47564
rect 38764 47500 38765 47564
rect 38699 47499 38765 47500
rect 37595 44844 37661 44845
rect 37595 44780 37596 44844
rect 37660 44780 37661 44844
rect 37595 44779 37661 44780
rect 37598 9349 37658 44779
rect 38702 10981 38762 47499
rect 39251 38860 39317 38861
rect 39251 38796 39252 38860
rect 39316 38796 39317 38860
rect 39251 38795 39317 38796
rect 39254 22110 39314 38795
rect 41827 31244 41893 31245
rect 41827 31180 41828 31244
rect 41892 31180 41893 31244
rect 41827 31179 41893 31180
rect 40539 24172 40605 24173
rect 40539 24108 40540 24172
rect 40604 24108 40605 24172
rect 40539 24107 40605 24108
rect 39254 22050 40050 22110
rect 38699 10980 38765 10981
rect 38699 10916 38700 10980
rect 38764 10916 38765 10980
rect 38699 10915 38765 10916
rect 37595 9348 37661 9349
rect 37595 9284 37596 9348
rect 37660 9284 37661 9348
rect 37595 9283 37661 9284
rect 35939 4044 36005 4045
rect 35939 3980 35940 4044
rect 36004 3980 36005 4044
rect 35939 3979 36005 3980
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 31155 3228 31221 3229
rect 31155 3164 31156 3228
rect 31220 3164 31221 3228
rect 31155 3163 31221 3164
rect 29131 3092 29197 3093
rect 29131 3028 29132 3092
rect 29196 3028 29197 3092
rect 29131 3027 29197 3028
rect 34928 2752 35248 3776
rect 39990 3637 40050 22050
rect 40542 12341 40602 24107
rect 40539 12340 40605 12341
rect 40539 12276 40540 12340
rect 40604 12276 40605 12340
rect 40539 12275 40605 12276
rect 41830 4045 41890 31179
rect 42566 5541 42626 59331
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 43851 56676 43917 56677
rect 43851 56612 43852 56676
rect 43916 56612 43917 56676
rect 43851 56611 43917 56612
rect 42563 5540 42629 5541
rect 42563 5476 42564 5540
rect 42628 5476 42629 5540
rect 42563 5475 42629 5476
rect 41827 4044 41893 4045
rect 41827 3980 41828 4044
rect 41892 3980 41893 4044
rect 41827 3979 41893 3980
rect 43854 3637 43914 56611
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 39987 3636 40053 3637
rect 39987 3572 39988 3636
rect 40052 3572 40053 3636
rect 39987 3571 40053 3572
rect 43851 3636 43917 3637
rect 43851 3572 43852 3636
rect 43916 3572 43917 3636
rect 43851 3571 43917 3572
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 27107 2548 27173 2549
rect 27107 2484 27108 2548
rect 27172 2484 27173 2548
rect 27107 2483 27173 2484
rect 26003 2412 26069 2413
rect 26003 2348 26004 2412
rect 26068 2348 26069 2412
rect 26003 2347 26069 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20240 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 23368 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 23000 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 27692 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 29072 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 29992 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 29348 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 30636 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 50692 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 22356 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 22632 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 40020 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 27600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 27048 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 35328 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 35604 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 38364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 2300 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 2300 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 2300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 30176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 52440 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 31556 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 32384 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 19688 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform -1 0 30176 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1676037725
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46
timestamp 1676037725
transform 1 0 5336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1676037725
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1676037725
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1676037725
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_102
timestamp 1676037725
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_128
timestamp 1676037725
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1676037725
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1676037725
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1676037725
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1676037725
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_214
timestamp 1676037725
transform 1 0 20792 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_218
timestamp 1676037725
transform 1 0 21160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1676037725
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1676037725
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1676037725
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_268
timestamp 1676037725
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1676037725
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_296
timestamp 1676037725
transform 1 0 28336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1676037725
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_315
timestamp 1676037725
transform 1 0 30084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_322
timestamp 1676037725
transform 1 0 30728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1676037725
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_345
timestamp 1676037725
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1676037725
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1676037725
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1676037725
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_401
timestamp 1676037725
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_411
timestamp 1676037725
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1676037725
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_439
timestamp 1676037725
transform 1 0 41492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1676037725
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_467
timestamp 1676037725
transform 1 0 44068 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_483
timestamp 1676037725
transform 1 0 45540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_487
timestamp 1676037725
transform 1 0 45908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_494
timestamp 1676037725
transform 1 0 46552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1676037725
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_513
timestamp 1676037725
transform 1 0 48300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_523
timestamp 1676037725
transform 1 0 49220 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1676037725
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1676037725
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_539
timestamp 1676037725
transform 1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_547
timestamp 1676037725
transform 1 0 51428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_555
timestamp 1676037725
transform 1 0 52164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1676037725
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_561
timestamp 1676037725
transform 1 0 52716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_569
timestamp 1676037725
transform 1 0 53452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_579
timestamp 1676037725
transform 1 0 54372 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1676037725
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 1676037725
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_597
timestamp 1676037725
transform 1 0 56028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_605
timestamp 1676037725
transform 1 0 56764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1676037725
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1676037725
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_623
timestamp 1676037725
transform 1 0 58420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_23
timestamp 1676037725
transform 1 0 3220 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_31
timestamp 1676037725
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1676037725
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_67
timestamp 1676037725
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1676037725
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_85
timestamp 1676037725
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1676037725
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1676037725
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1676037725
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_126
timestamp 1676037725
transform 1 0 12696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1676037725
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_146
timestamp 1676037725
transform 1 0 14536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1676037725
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1676037725
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1676037725
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1676037725
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_198
timestamp 1676037725
transform 1 0 19320 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1676037725
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_250
timestamp 1676037725
transform 1 0 24104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_254
timestamp 1676037725
transform 1 0 24472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_258
timestamp 1676037725
transform 1 0 24840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_268
timestamp 1676037725
transform 1 0 25760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1676037725
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_316
timestamp 1676037725
transform 1 0 30176 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_322
timestamp 1676037725
transform 1 0 30728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_345
timestamp 1676037725
transform 1 0 32844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_369
timestamp 1676037725
transform 1 0 35052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_379
timestamp 1676037725
transform 1 0 35972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_389
timestamp 1676037725
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_404
timestamp 1676037725
transform 1 0 38272 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_414
timestamp 1676037725
transform 1 0 39192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1676037725
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_434
timestamp 1676037725
transform 1 0 41032 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1676037725
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_465
timestamp 1676037725
transform 1 0 43884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_481
timestamp 1676037725
transform 1 0 45356 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_489
timestamp 1676037725
transform 1 0 46092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1676037725
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_513
timestamp 1676037725
transform 1 0 48300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_523
timestamp 1676037725
transform 1 0 49220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_533
timestamp 1676037725
transform 1 0 50140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_541
timestamp 1676037725
transform 1 0 50876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_549
timestamp 1676037725
transform 1 0 51612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_557
timestamp 1676037725
transform 1 0 52348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1676037725
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_567
timestamp 1676037725
transform 1 0 53268 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_581
timestamp 1676037725
transform 1 0 54556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_591
timestamp 1676037725
transform 1 0 55476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_601
timestamp 1676037725
transform 1 0 56396 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_607
timestamp 1676037725
transform 1 0 56948 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1676037725
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_617
timestamp 1676037725
transform 1 0 57868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_623
timestamp 1676037725
transform 1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_11
timestamp 1676037725
transform 1 0 2116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1676037725
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_46
timestamp 1676037725
transform 1 0 5336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_54
timestamp 1676037725
transform 1 0 6072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_62
timestamp 1676037725
transform 1 0 6808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1676037725
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1676037725
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_107
timestamp 1676037725
transform 1 0 10948 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_115
timestamp 1676037725
transform 1 0 11684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_120
timestamp 1676037725
transform 1 0 12144 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1676037725
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_149
timestamp 1676037725
transform 1 0 14812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_157
timestamp 1676037725
transform 1 0 15548 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_166
timestamp 1676037725
transform 1 0 16376 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_174
timestamp 1676037725
transform 1 0 17112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1676037725
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_201
timestamp 1676037725
transform 1 0 19596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_218
timestamp 1676037725
transform 1 0 21160 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1676037725
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_264
timestamp 1676037725
transform 1 0 25392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_274
timestamp 1676037725
transform 1 0 26312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_278
timestamp 1676037725
transform 1 0 26680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_286
timestamp 1676037725
transform 1 0 27416 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_299
timestamp 1676037725
transform 1 0 28612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1676037725
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_323
timestamp 1676037725
transform 1 0 30820 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_334
timestamp 1676037725
transform 1 0 31832 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_373
timestamp 1676037725
transform 1 0 35420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_386
timestamp 1676037725
transform 1 0 36616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_409
timestamp 1676037725
transform 1 0 38732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_417
timestamp 1676037725
transform 1 0 39468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_438
timestamp 1676037725
transform 1 0 41400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_446
timestamp 1676037725
transform 1 0 42136 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_471
timestamp 1676037725
transform 1 0 44436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_483
timestamp 1676037725
transform 1 0 45540 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_491
timestamp 1676037725
transform 1 0 46276 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_503
timestamp 1676037725
transform 1 0 47380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_511
timestamp 1676037725
transform 1 0 48116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_519
timestamp 1676037725
transform 1 0 48852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_527
timestamp 1676037725
transform 1 0 49588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1676037725
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1676037725
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_539
timestamp 1676037725
transform 1 0 50692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_547
timestamp 1676037725
transform 1 0 51428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_555
timestamp 1676037725
transform 1 0 52164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_563
timestamp 1676037725
transform 1 0 52900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_571
timestamp 1676037725
transform 1 0 53636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_579
timestamp 1676037725
transform 1 0 54372 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1676037725
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_589
timestamp 1676037725
transform 1 0 55292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_595
timestamp 1676037725
transform 1 0 55844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_603
timestamp 1676037725
transform 1 0 56580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_622
timestamp 1676037725
transform 1 0 58328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_11
timestamp 1676037725
transform 1 0 2116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_23
timestamp 1676037725
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1676037725
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_47
timestamp 1676037725
transform 1 0 5428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1676037725
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_63
timestamp 1676037725
transform 1 0 6900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1676037725
transform 1 0 7636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_92
timestamp 1676037725
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_102
timestamp 1676037725
transform 1 0 10488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_119
timestamp 1676037725
transform 1 0 12052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1676037725
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_139
timestamp 1676037725
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_155
timestamp 1676037725
transform 1 0 15364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1676037725
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1676037725
transform 1 0 17572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_189
timestamp 1676037725
transform 1 0 18492 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_199
timestamp 1676037725
transform 1 0 19412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1676037725
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_231
timestamp 1676037725
transform 1 0 22356 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_238
timestamp 1676037725
transform 1 0 23000 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_258
timestamp 1676037725
transform 1 0 24840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_268
timestamp 1676037725
transform 1 0 25760 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_274
timestamp 1676037725
transform 1 0 26312 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1676037725
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_300
timestamp 1676037725
transform 1 0 28704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_307
timestamp 1676037725
transform 1 0 29348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_325
timestamp 1676037725
transform 1 0 31004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1676037725
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_348
timestamp 1676037725
transform 1 0 33120 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_358
timestamp 1676037725
transform 1 0 34040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_368
timestamp 1676037725
transform 1 0 34960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_378
timestamp 1676037725
transform 1 0 35880 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1676037725
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_404
timestamp 1676037725
transform 1 0 38272 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_425
timestamp 1676037725
transform 1 0 40204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_433
timestamp 1676037725
transform 1 0 40940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_465
timestamp 1676037725
transform 1 0 43884 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_481
timestamp 1676037725
transform 1 0 45356 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_489
timestamp 1676037725
transform 1 0 46092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_511
timestamp 1676037725
transform 1 0 48116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_516
timestamp 1676037725
transform 1 0 48576 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_528
timestamp 1676037725
transform 1 0 49680 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_540
timestamp 1676037725
transform 1 0 50784 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_552
timestamp 1676037725
transform 1 0 51888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_558
timestamp 1676037725
transform 1 0 52440 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_561
timestamp 1676037725
transform 1 0 52716 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_567
timestamp 1676037725
transform 1 0 53268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_575
timestamp 1676037725
transform 1 0 54004 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1676037725
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1676037725
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1676037725
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1676037725
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_617
timestamp 1676037725
transform 1 0 57868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_623
timestamp 1676037725
transform 1 0 58420 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_57
timestamp 1676037725
transform 1 0 6348 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_61
timestamp 1676037725
transform 1 0 6716 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_66
timestamp 1676037725
transform 1 0 7176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_74
timestamp 1676037725
transform 1 0 7912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_100
timestamp 1676037725
transform 1 0 10304 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 1676037725
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_114
timestamp 1676037725
transform 1 0 11592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_119
timestamp 1676037725
transform 1 0 12052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_127
timestamp 1676037725
transform 1 0 12788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1676037725
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_149
timestamp 1676037725
transform 1 0 14812 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_161
timestamp 1676037725
transform 1 0 15916 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_169
timestamp 1676037725
transform 1 0 16652 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_174
timestamp 1676037725
transform 1 0 17112 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_184
timestamp 1676037725
transform 1 0 18032 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1676037725
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_208
timestamp 1676037725
transform 1 0 20240 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_229
timestamp 1676037725
transform 1 0 22172 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_237
timestamp 1676037725
transform 1 0 22908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_264
timestamp 1676037725
transform 1 0 25392 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_272
timestamp 1676037725
transform 1 0 26128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_284
timestamp 1676037725
transform 1 0 27232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_293
timestamp 1676037725
transform 1 0 28060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1676037725
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_317
timestamp 1676037725
transform 1 0 30268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_329
timestamp 1676037725
transform 1 0 31372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_337
timestamp 1676037725
transform 1 0 32108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_348
timestamp 1676037725
transform 1 0 33120 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_371
timestamp 1676037725
transform 1 0 35236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_375
timestamp 1676037725
transform 1 0 35604 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_393
timestamp 1676037725
transform 1 0 37260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_402
timestamp 1676037725
transform 1 0 38088 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_408
timestamp 1676037725
transform 1 0 38640 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_414
timestamp 1676037725
transform 1 0 39192 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_427
timestamp 1676037725
transform 1 0 40388 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_435
timestamp 1676037725
transform 1 0 41124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_443
timestamp 1676037725
transform 1 0 41860 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_451
timestamp 1676037725
transform 1 0 42596 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_461
timestamp 1676037725
transform 1 0 43516 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_473
timestamp 1676037725
transform 1 0 44620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_483
timestamp 1676037725
transform 1 0 45540 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_491
timestamp 1676037725
transform 1 0 46276 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_503
timestamp 1676037725
transform 1 0 47380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_515
timestamp 1676037725
transform 1 0 48484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_527
timestamp 1676037725
transform 1 0 49588 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1676037725
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_533
timestamp 1676037725
transform 1 0 50140 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_546
timestamp 1676037725
transform 1 0 51336 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_558
timestamp 1676037725
transform 1 0 52440 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_570
timestamp 1676037725
transform 1 0 53544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_582
timestamp 1676037725
transform 1 0 54648 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1676037725
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1676037725
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_613
timestamp 1676037725
transform 1 0 57500 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_623
timestamp 1676037725
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_11
timestamp 1676037725
transform 1 0 2116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_23
timestamp 1676037725
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1676037725
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1676037725
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_91
timestamp 1676037725
transform 1 0 9476 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1676037725
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1676037725
transform 1 0 12236 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_126
timestamp 1676037725
transform 1 0 12696 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_132
timestamp 1676037725
transform 1 0 13248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1676037725
transform 1 0 13892 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_147
timestamp 1676037725
transform 1 0 14628 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_159
timestamp 1676037725
transform 1 0 15732 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_176
timestamp 1676037725
transform 1 0 17296 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_183
timestamp 1676037725
transform 1 0 17940 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1676037725
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_210
timestamp 1676037725
transform 1 0 20424 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_239
timestamp 1676037725
transform 1 0 23092 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_251
timestamp 1676037725
transform 1 0 24196 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_263
timestamp 1676037725
transform 1 0 25300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_270
timestamp 1676037725
transform 1 0 25944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 1676037725
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_289
timestamp 1676037725
transform 1 0 27692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_301
timestamp 1676037725
transform 1 0 28796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_309
timestamp 1676037725
transform 1 0 29532 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_324
timestamp 1676037725
transform 1 0 30912 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_343
timestamp 1676037725
transform 1 0 32660 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_348
timestamp 1676037725
transform 1 0 33120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_356
timestamp 1676037725
transform 1 0 33856 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_364
timestamp 1676037725
transform 1 0 34592 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_383
timestamp 1676037725
transform 1 0 36340 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_399
timestamp 1676037725
transform 1 0 37812 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_423
timestamp 1676037725
transform 1 0 40020 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_431
timestamp 1676037725
transform 1 0 40756 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_439
timestamp 1676037725
transform 1 0 41492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_455
timestamp 1676037725
transform 1 0 42964 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_463
timestamp 1676037725
transform 1 0 43700 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_471
timestamp 1676037725
transform 1 0 44436 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_479
timestamp 1676037725
transform 1 0 45172 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_489
timestamp 1676037725
transform 1 0 46092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_501
timestamp 1676037725
transform 1 0 47196 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_513
timestamp 1676037725
transform 1 0 48300 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_531
timestamp 1676037725
transform 1 0 49956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_543
timestamp 1676037725
transform 1 0 51060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_555
timestamp 1676037725
transform 1 0 52164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1676037725
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1676037725
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1676037725
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1676037725
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1676037725
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1676037725
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1676037725
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_617
timestamp 1676037725
transform 1 0 57868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_623
timestamp 1676037725
transform 1 0 58420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_11
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1676037725
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_94
timestamp 1676037725
transform 1 0 9752 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_100
timestamp 1676037725
transform 1 0 10304 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_107
timestamp 1676037725
transform 1 0 10948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_119
timestamp 1676037725
transform 1 0 12052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_131
timestamp 1676037725
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_169
timestamp 1676037725
transform 1 0 16652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_219
timestamp 1676037725
transform 1 0 21252 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_236
timestamp 1676037725
transform 1 0 22816 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_246
timestamp 1676037725
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_263
timestamp 1676037725
transform 1 0 25300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_267
timestamp 1676037725
transform 1 0 25668 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_297
timestamp 1676037725
transform 1 0 28428 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1676037725
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_314
timestamp 1676037725
transform 1 0 29992 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_318
timestamp 1676037725
transform 1 0 30360 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_324
timestamp 1676037725
transform 1 0 30912 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_344
timestamp 1676037725
transform 1 0 32752 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_354
timestamp 1676037725
transform 1 0 33672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1676037725
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_371
timestamp 1676037725
transform 1 0 35236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_388
timestamp 1676037725
transform 1 0 36800 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_396
timestamp 1676037725
transform 1 0 37536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_403
timestamp 1676037725
transform 1 0 38180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_407
timestamp 1676037725
transform 1 0 38548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_418
timestamp 1676037725
transform 1 0 39560 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_441
timestamp 1676037725
transform 1 0 41676 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_453
timestamp 1676037725
transform 1 0 42780 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_465
timestamp 1676037725
transform 1 0 43884 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_473
timestamp 1676037725
transform 1 0 44620 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1676037725
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1676037725
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1676037725
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1676037725
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1676037725
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1676037725
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1676037725
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1676037725
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_601
timestamp 1676037725
transform 1 0 56396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_613
timestamp 1676037725
transform 1 0 57500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_623
timestamp 1676037725
transform 1 0 58420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_11
timestamp 1676037725
transform 1 0 2116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_23
timestamp 1676037725
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1676037725
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1676037725
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_94
timestamp 1676037725
transform 1 0 9752 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1676037725
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1676037725
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_143
timestamp 1676037725
transform 1 0 14260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1676037725
transform 1 0 14996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_182
timestamp 1676037725
transform 1 0 17848 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_192
timestamp 1676037725
transform 1 0 18768 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_198
timestamp 1676037725
transform 1 0 19320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1676037725
transform 1 0 20884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_231
timestamp 1676037725
transform 1 0 22356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_247
timestamp 1676037725
transform 1 0 23828 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_255
timestamp 1676037725
transform 1 0 24564 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_294
timestamp 1676037725
transform 1 0 28152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_307
timestamp 1676037725
transform 1 0 29348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_320
timestamp 1676037725
transform 1 0 30544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_369
timestamp 1676037725
transform 1 0 35052 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_379
timestamp 1676037725
transform 1 0 35972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_387
timestamp 1676037725
transform 1 0 36708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_411
timestamp 1676037725
transform 1 0 38916 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_423
timestamp 1676037725
transform 1 0 40020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_435
timestamp 1676037725
transform 1 0 41124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_489
timestamp 1676037725
transform 1 0 46092 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_495
timestamp 1676037725
transform 1 0 46644 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1676037725
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1676037725
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1676037725
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1676037725
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1676037725
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1676037725
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1676037725
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1676037725
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1676037725
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1676037725
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_617
timestamp 1676037725
transform 1 0 57868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_623
timestamp 1676037725
transform 1 0 58420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_11
timestamp 1676037725
transform 1 0 2116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1676037725
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_95
timestamp 1676037725
transform 1 0 9844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_103
timestamp 1676037725
transform 1 0 10580 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_112
timestamp 1676037725
transform 1 0 11408 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_124
timestamp 1676037725
transform 1 0 12512 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_132
timestamp 1676037725
transform 1 0 13248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_149
timestamp 1676037725
transform 1 0 14812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_172
timestamp 1676037725
transform 1 0 16928 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_185
timestamp 1676037725
transform 1 0 18124 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1676037725
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_222
timestamp 1676037725
transform 1 0 21528 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1676037725
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_266
timestamp 1676037725
transform 1 0 25576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_284
timestamp 1676037725
transform 1 0 27232 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_323
timestamp 1676037725
transform 1 0 30820 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_334
timestamp 1676037725
transform 1 0 31832 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_346
timestamp 1676037725
transform 1 0 32936 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_354
timestamp 1676037725
transform 1 0 33672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1676037725
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_376
timestamp 1676037725
transform 1 0 35696 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_388
timestamp 1676037725
transform 1 0 36800 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_400
timestamp 1676037725
transform 1 0 37904 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_412
timestamp 1676037725
transform 1 0 39008 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_495
timestamp 1676037725
transform 1 0 46644 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_505
timestamp 1676037725
transform 1 0 47564 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_517
timestamp 1676037725
transform 1 0 48668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_529
timestamp 1676037725
transform 1 0 49772 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1676037725
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1676037725
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1676037725
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1676037725
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1676037725
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1676037725
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1676037725
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_601
timestamp 1676037725
transform 1 0 56396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_605
timestamp 1676037725
transform 1 0 56764 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_622
timestamp 1676037725
transform 1 0 58328 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1676037725
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_119
timestamp 1676037725
transform 1 0 12052 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_129
timestamp 1676037725
transform 1 0 12972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_141
timestamp 1676037725
transform 1 0 14076 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1676037725
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp 1676037725
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_194
timestamp 1676037725
transform 1 0 18952 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_231
timestamp 1676037725
transform 1 0 22356 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_239
timestamp 1676037725
transform 1 0 23092 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_262
timestamp 1676037725
transform 1 0 25208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_287
timestamp 1676037725
transform 1 0 27508 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_294
timestamp 1676037725
transform 1 0 28152 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_298
timestamp 1676037725
transform 1 0 28520 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_319
timestamp 1676037725
transform 1 0 30452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1676037725
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_357
timestamp 1676037725
transform 1 0 33948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_376
timestamp 1676037725
transform 1 0 35696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_380
timestamp 1676037725
transform 1 0 36064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1676037725
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_398
timestamp 1676037725
transform 1 0 37720 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_410
timestamp 1676037725
transform 1 0 38824 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_422
timestamp 1676037725
transform 1 0 39928 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_434
timestamp 1676037725
transform 1 0 41032 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1676037725
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_469
timestamp 1676037725
transform 1 0 44252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_474
timestamp 1676037725
transform 1 0 44712 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_478
timestamp 1676037725
transform 1 0 45080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_482
timestamp 1676037725
transform 1 0 45448 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_495
timestamp 1676037725
transform 1 0 46644 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1676037725
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1676037725
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1676037725
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1676037725
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1676037725
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1676037725
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_585
timestamp 1676037725
transform 1 0 54924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_593
timestamp 1676037725
transform 1 0 55660 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_598
timestamp 1676037725
transform 1 0 56120 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_611
timestamp 1676037725
transform 1 0 57316 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1676037725
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_617
timestamp 1676037725
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_622
timestamp 1676037725
transform 1 0 58328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_11
timestamp 1676037725
transform 1 0 2116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1676037725
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 1676037725
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1676037725
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1676037725
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_101
timestamp 1676037725
transform 1 0 10396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1676037725
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1676037725
transform 1 0 16100 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_186
timestamp 1676037725
transform 1 0 18216 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_208
timestamp 1676037725
transform 1 0 20240 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_220
timestamp 1676037725
transform 1 0 21344 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_232
timestamp 1676037725
transform 1 0 22448 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_243
timestamp 1676037725
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_262
timestamp 1676037725
transform 1 0 25208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_270
timestamp 1676037725
transform 1 0 25944 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1676037725
transform 1 0 26496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_293
timestamp 1676037725
transform 1 0 28060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1676037725
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_325
timestamp 1676037725
transform 1 0 31004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_338
timestamp 1676037725
transform 1 0 32200 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_349
timestamp 1676037725
transform 1 0 33212 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_362
timestamp 1676037725
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_373
timestamp 1676037725
transform 1 0 35420 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_379
timestamp 1676037725
transform 1 0 35972 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_397
timestamp 1676037725
transform 1 0 37628 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_409
timestamp 1676037725
transform 1 0 38732 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_417
timestamp 1676037725
transform 1 0 39468 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_454
timestamp 1676037725
transform 1 0 42872 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_462
timestamp 1676037725
transform 1 0 43608 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_473
timestamp 1676037725
transform 1 0 44620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_484
timestamp 1676037725
transform 1 0 45632 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_499
timestamp 1676037725
transform 1 0 47012 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_511
timestamp 1676037725
transform 1 0 48116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_523
timestamp 1676037725
transform 1 0 49220 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1676037725
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1676037725
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1676037725
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1676037725
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1676037725
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1676037725
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1676037725
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_589
timestamp 1676037725
transform 1 0 55292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_594
timestamp 1676037725
transform 1 0 55752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_602
timestamp 1676037725
transform 1 0 56488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_622
timestamp 1676037725
transform 1 0 58328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_11
timestamp 1676037725
transform 1 0 2116 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_23
timestamp 1676037725
transform 1 0 3220 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_35
timestamp 1676037725
transform 1 0 4324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_47
timestamp 1676037725
transform 1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_143
timestamp 1676037725
transform 1 0 14260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_153
timestamp 1676037725
transform 1 0 15180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_204
timestamp 1676037725
transform 1 0 19872 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_248
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_257
timestamp 1676037725
transform 1 0 24748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_265
timestamp 1676037725
transform 1 0 25484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1676037725
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_292
timestamp 1676037725
transform 1 0 27968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_321
timestamp 1676037725
transform 1 0 30636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1676037725
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_343
timestamp 1676037725
transform 1 0 32660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_352
timestamp 1676037725
transform 1 0 33488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_364
timestamp 1676037725
transform 1 0 34592 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_381
timestamp 1676037725
transform 1 0 36156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1676037725
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_404
timestamp 1676037725
transform 1 0 38272 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_408
timestamp 1676037725
transform 1 0 38640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_425
timestamp 1676037725
transform 1 0 40204 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_437
timestamp 1676037725
transform 1 0 41308 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_445
timestamp 1676037725
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_476
timestamp 1676037725
transform 1 0 44896 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_486
timestamp 1676037725
transform 1 0 45816 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_498
timestamp 1676037725
transform 1 0 46920 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1676037725
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1676037725
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1676037725
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1676037725
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1676037725
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1676037725
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1676037725
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_597
timestamp 1676037725
transform 1 0 56028 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_604
timestamp 1676037725
transform 1 0 56672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_614
timestamp 1676037725
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1676037725
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_11
timestamp 1676037725
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1676037725
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp 1676037725
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_155
timestamp 1676037725
transform 1 0 15364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_178
timestamp 1676037725
transform 1 0 17480 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1676037725
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_216
timestamp 1676037725
transform 1 0 20976 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_224
timestamp 1676037725
transform 1 0 21712 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_236
timestamp 1676037725
transform 1 0 22816 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_242
timestamp 1676037725
transform 1 0 23368 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_276
timestamp 1676037725
transform 1 0 26496 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_288
timestamp 1676037725
transform 1 0 27600 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_293
timestamp 1676037725
transform 1 0 28060 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_306
timestamp 1676037725
transform 1 0 29256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_322
timestamp 1676037725
transform 1 0 30728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_343
timestamp 1676037725
transform 1 0 32660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_353
timestamp 1676037725
transform 1 0 33580 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_361
timestamp 1676037725
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_386
timestamp 1676037725
transform 1 0 36616 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_399
timestamp 1676037725
transform 1 0 37812 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_407
timestamp 1676037725
transform 1 0 38548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_412
timestamp 1676037725
transform 1 0 39008 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_440
timestamp 1676037725
transform 1 0 41584 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_452
timestamp 1676037725
transform 1 0 42688 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_460
timestamp 1676037725
transform 1 0 43424 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_474
timestamp 1676037725
transform 1 0 44712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_485
timestamp 1676037725
transform 1 0 45724 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_492
timestamp 1676037725
transform 1 0 46368 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_504
timestamp 1676037725
transform 1 0 47472 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_516
timestamp 1676037725
transform 1 0 48576 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_528
timestamp 1676037725
transform 1 0 49680 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1676037725
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1676037725
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1676037725
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1676037725
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1676037725
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1676037725
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_589
timestamp 1676037725
transform 1 0 55292 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_597
timestamp 1676037725
transform 1 0 56028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_602
timestamp 1676037725
transform 1 0 56488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_622
timestamp 1676037725
transform 1 0 58328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_11
timestamp 1676037725
transform 1 0 2116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_23
timestamp 1676037725
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_35
timestamp 1676037725
transform 1 0 4324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1676037725
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_89
timestamp 1676037725
transform 1 0 9292 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_101
timestamp 1676037725
transform 1 0 10396 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1676037725
transform 1 0 12972 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_138
timestamp 1676037725
transform 1 0 13800 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_146
timestamp 1676037725
transform 1 0 14536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1676037725
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_194
timestamp 1676037725
transform 1 0 18952 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_202
timestamp 1676037725
transform 1 0 19688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1676037725
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_245
timestamp 1676037725
transform 1 0 23644 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_252
timestamp 1676037725
transform 1 0 24288 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_289
timestamp 1676037725
transform 1 0 27692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_304
timestamp 1676037725
transform 1 0 29072 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_315
timestamp 1676037725
transform 1 0 30084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1676037725
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_345
timestamp 1676037725
transform 1 0 32844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_356
timestamp 1676037725
transform 1 0 33856 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_368
timestamp 1676037725
transform 1 0 34960 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_376
timestamp 1676037725
transform 1 0 35696 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_382
timestamp 1676037725
transform 1 0 36248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_390
timestamp 1676037725
transform 1 0 36984 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_403
timestamp 1676037725
transform 1 0 38180 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_415
timestamp 1676037725
transform 1 0 39284 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_427
timestamp 1676037725
transform 1 0 40388 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_431
timestamp 1676037725
transform 1 0 40756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_443
timestamp 1676037725
transform 1 0 41860 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_470
timestamp 1676037725
transform 1 0 44344 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_478
timestamp 1676037725
transform 1 0 45080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_495
timestamp 1676037725
transform 1 0 46644 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1676037725
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1676037725
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1676037725
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1676037725
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1676037725
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1676037725
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1676037725
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_597
timestamp 1676037725
transform 1 0 56028 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_605
timestamp 1676037725
transform 1 0 56764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_611
timestamp 1676037725
transform 1 0 57316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1676037725
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1676037725
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_11
timestamp 1676037725
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1676037725
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_105
timestamp 1676037725
transform 1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_114
timestamp 1676037725
transform 1 0 11592 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_126
timestamp 1676037725
transform 1 0 12696 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1676037725
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_152
timestamp 1676037725
transform 1 0 15088 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_156
timestamp 1676037725
transform 1 0 15456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_174
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1676037725
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1676037725
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_232
timestamp 1676037725
transform 1 0 22448 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_244
timestamp 1676037725
transform 1 0 23552 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_264
timestamp 1676037725
transform 1 0 25392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_285
timestamp 1676037725
transform 1 0 27324 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_296
timestamp 1676037725
transform 1 0 28336 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1676037725
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_318
timestamp 1676037725
transform 1 0 30360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_330
timestamp 1676037725
transform 1 0 31464 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_341
timestamp 1676037725
transform 1 0 32476 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_353
timestamp 1676037725
transform 1 0 33580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 1676037725
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_374
timestamp 1676037725
transform 1 0 35512 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_386
timestamp 1676037725
transform 1 0 36616 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_400
timestamp 1676037725
transform 1 0 37904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_412
timestamp 1676037725
transform 1 0 39008 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_446
timestamp 1676037725
transform 1 0 42136 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_458
timestamp 1676037725
transform 1 0 43240 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_464
timestamp 1676037725
transform 1 0 43792 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_473
timestamp 1676037725
transform 1 0 44620 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_483
timestamp 1676037725
transform 1 0 45540 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_490
timestamp 1676037725
transform 1 0 46184 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_496
timestamp 1676037725
transform 1 0 46736 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_517
timestamp 1676037725
transform 1 0 48668 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_529
timestamp 1676037725
transform 1 0 49772 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1676037725
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1676037725
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1676037725
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1676037725
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1676037725
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1676037725
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1676037725
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_601
timestamp 1676037725
transform 1 0 56396 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_613
timestamp 1676037725
transform 1 0 57500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_623
timestamp 1676037725
transform 1 0 58420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_11
timestamp 1676037725
transform 1 0 2116 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_23
timestamp 1676037725
transform 1 0 3220 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_35
timestamp 1676037725
transform 1 0 4324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1676037725
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_96
timestamp 1676037725
transform 1 0 9936 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1676037725
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_121
timestamp 1676037725
transform 1 0 12236 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_127
timestamp 1676037725
transform 1 0 12788 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_145
timestamp 1676037725
transform 1 0 14444 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_154
timestamp 1676037725
transform 1 0 15272 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1676037725
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1676037725
transform 1 0 18032 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_188
timestamp 1676037725
transform 1 0 18400 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_218
timestamp 1676037725
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_236
timestamp 1676037725
transform 1 0 22816 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_245
timestamp 1676037725
transform 1 0 23644 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_261
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_294
timestamp 1676037725
transform 1 0 28152 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_317
timestamp 1676037725
transform 1 0 30268 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1676037725
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_345
timestamp 1676037725
transform 1 0 32844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_356
timestamp 1676037725
transform 1 0 33856 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_367
timestamp 1676037725
transform 1 0 34868 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_377
timestamp 1676037725
transform 1 0 35788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1676037725
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_408
timestamp 1676037725
transform 1 0 38640 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_420
timestamp 1676037725
transform 1 0 39744 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_428
timestamp 1676037725
transform 1 0 40480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_446
timestamp 1676037725
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_467
timestamp 1676037725
transform 1 0 44068 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_488
timestamp 1676037725
transform 1 0 46000 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1676037725
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1676037725
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1676037725
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1676037725
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1676037725
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1676037725
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1676037725
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1676037725
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1676037725
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1676037725
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_612
timestamp 1676037725
transform 1 0 57408 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_617
timestamp 1676037725
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_11
timestamp 1676037725
transform 1 0 2116 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1676037725
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_105
timestamp 1676037725
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_114
timestamp 1676037725
transform 1 0 11592 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_126
timestamp 1676037725
transform 1 0 12696 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1676037725
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_149
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1676037725
transform 1 0 15272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_172
timestamp 1676037725
transform 1 0 16928 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_176
timestamp 1676037725
transform 1 0 17296 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_183
timestamp 1676037725
transform 1 0 17940 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_217
timestamp 1676037725
transform 1 0 21068 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_225
timestamp 1676037725
transform 1 0 21804 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_237
timestamp 1676037725
transform 1 0 22908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1676037725
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_269
timestamp 1676037725
transform 1 0 25852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_277
timestamp 1676037725
transform 1 0 26588 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_323
timestamp 1676037725
transform 1 0 30820 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_327
timestamp 1676037725
transform 1 0 31188 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_332
timestamp 1676037725
transform 1 0 31648 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_339
timestamp 1676037725
transform 1 0 32292 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_345
timestamp 1676037725
transform 1 0 32844 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1676037725
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_380
timestamp 1676037725
transform 1 0 36064 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_392
timestamp 1676037725
transform 1 0 37168 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_411
timestamp 1676037725
transform 1 0 38916 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_429
timestamp 1676037725
transform 1 0 40572 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_446
timestamp 1676037725
transform 1 0 42136 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_464
timestamp 1676037725
transform 1 0 43792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1676037725
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_500
timestamp 1676037725
transform 1 0 47104 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_512
timestamp 1676037725
transform 1 0 48208 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_524
timestamp 1676037725
transform 1 0 49312 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1676037725
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1676037725
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_557
timestamp 1676037725
transform 1 0 52348 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_572
timestamp 1676037725
transform 1 0 53728 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_584
timestamp 1676037725
transform 1 0 54832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_589
timestamp 1676037725
transform 1 0 55292 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_597
timestamp 1676037725
transform 1 0 56028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_602
timestamp 1676037725
transform 1 0 56488 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_622
timestamp 1676037725
transform 1 0 58328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1676037725
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1676037725
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1676037725
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1676037725
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_122
timestamp 1676037725
transform 1 0 12328 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_134
timestamp 1676037725
transform 1 0 13432 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_142
timestamp 1676037725
transform 1 0 14168 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_155
timestamp 1676037725
transform 1 0 15364 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1676037725
transform 1 0 17572 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_187
timestamp 1676037725
transform 1 0 18308 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_199
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_214
timestamp 1676037725
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_222
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_249
timestamp 1676037725
transform 1 0 24012 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_259
timestamp 1676037725
transform 1 0 24932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_272
timestamp 1676037725
transform 1 0 26128 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_299
timestamp 1676037725
transform 1 0 28612 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_314
timestamp 1676037725
transform 1 0 29992 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_320
timestamp 1676037725
transform 1 0 30544 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_324
timestamp 1676037725
transform 1 0 30912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_331
timestamp 1676037725
transform 1 0 31556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_345
timestamp 1676037725
transform 1 0 32844 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_355
timestamp 1676037725
transform 1 0 33764 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_363
timestamp 1676037725
transform 1 0 34500 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_380
timestamp 1676037725
transform 1 0 36064 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_405
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1676037725
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_485
timestamp 1676037725
transform 1 0 45724 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_500
timestamp 1676037725
transform 1 0 47104 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1676037725
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1676037725
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1676037725
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1676037725
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1676037725
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1676037725
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1676037725
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1676037725
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_597
timestamp 1676037725
transform 1 0 56028 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_605
timestamp 1676037725
transform 1 0 56764 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_614
timestamp 1676037725
transform 1 0 57592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1676037725
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1676037725
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_17
timestamp 1676037725
transform 1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1676037725
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_101
timestamp 1676037725
transform 1 0 10396 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_105
timestamp 1676037725
transform 1 0 10764 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_111
timestamp 1676037725
transform 1 0 11316 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_116
timestamp 1676037725
transform 1 0 11776 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_128
timestamp 1676037725
transform 1 0 12880 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_134
timestamp 1676037725
transform 1 0 13432 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_150
timestamp 1676037725
transform 1 0 14904 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_158
timestamp 1676037725
transform 1 0 15640 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_164
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_176
timestamp 1676037725
transform 1 0 17296 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_184
timestamp 1676037725
transform 1 0 18032 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1676037725
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1676037725
transform 1 0 20700 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_230
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_242
timestamp 1676037725
transform 1 0 23368 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_257
timestamp 1676037725
transform 1 0 24748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_263
timestamp 1676037725
transform 1 0 25300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_272
timestamp 1676037725
transform 1 0 26128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_280
timestamp 1676037725
transform 1 0 26864 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_291
timestamp 1676037725
transform 1 0 27876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1676037725
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1676037725
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_313
timestamp 1676037725
transform 1 0 29900 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_320
timestamp 1676037725
transform 1 0 30544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_324
timestamp 1676037725
transform 1 0 30912 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_329
timestamp 1676037725
transform 1 0 31372 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_336
timestamp 1676037725
transform 1 0 32016 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_348
timestamp 1676037725
transform 1 0 33120 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1676037725
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_378
timestamp 1676037725
transform 1 0 35880 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1676037725
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1676037725
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_431
timestamp 1676037725
transform 1 0 40756 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_443
timestamp 1676037725
transform 1 0 41860 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_455
timestamp 1676037725
transform 1 0 42964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_467
timestamp 1676037725
transform 1 0 44068 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1676037725
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1676037725
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1676037725
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1676037725
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1676037725
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1676037725
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1676037725
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1676037725
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1676037725
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1676037725
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1676037725
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_613
timestamp 1676037725
transform 1 0 57500 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_623
timestamp 1676037725
transform 1 0 58420 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_101
timestamp 1676037725
transform 1 0 10396 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_106
timestamp 1676037725
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_119
timestamp 1676037725
transform 1 0 12052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_127
timestamp 1676037725
transform 1 0 12788 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_135
timestamp 1676037725
transform 1 0 13524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_142
timestamp 1676037725
transform 1 0 14168 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_155
timestamp 1676037725
transform 1 0 15364 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1676037725
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_175
timestamp 1676037725
transform 1 0 17204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_189
timestamp 1676037725
transform 1 0 18492 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_201
timestamp 1676037725
transform 1 0 19596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_209
timestamp 1676037725
transform 1 0 20332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_231
timestamp 1676037725
transform 1 0 22356 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_239
timestamp 1676037725
transform 1 0 23092 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_251
timestamp 1676037725
transform 1 0 24196 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_257
timestamp 1676037725
transform 1 0 24748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1676037725
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_287
timestamp 1676037725
transform 1 0 27508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_319
timestamp 1676037725
transform 1 0 30452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1676037725
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_341
timestamp 1676037725
transform 1 0 32476 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_351
timestamp 1676037725
transform 1 0 33396 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_371
timestamp 1676037725
transform 1 0 35236 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_377
timestamp 1676037725
transform 1 0 35788 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1676037725
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1676037725
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1676037725
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_441
timestamp 1676037725
transform 1 0 41676 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_446
timestamp 1676037725
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_458
timestamp 1676037725
transform 1 0 43240 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_470
timestamp 1676037725
transform 1 0 44344 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_482
timestamp 1676037725
transform 1 0 45448 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_494
timestamp 1676037725
transform 1 0 46552 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1676037725
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1676037725
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1676037725
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1676037725
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1676037725
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1676037725
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1676037725
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1676037725
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1676037725
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1676037725
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1676037725
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1676037725
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_11
timestamp 1676037725
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1676037725
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_101
timestamp 1676037725
transform 1 0 10396 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_107
timestamp 1676037725
transform 1 0 10948 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_115
timestamp 1676037725
transform 1 0 11684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_126
timestamp 1676037725
transform 1 0 12696 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_147
timestamp 1676037725
transform 1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_158
timestamp 1676037725
transform 1 0 15640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_168
timestamp 1676037725
transform 1 0 16560 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_172
timestamp 1676037725
transform 1 0 16928 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1676037725
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1676037725
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_203
timestamp 1676037725
transform 1 0 19780 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_212
timestamp 1676037725
transform 1 0 20608 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1676037725
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1676037725
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_260
timestamp 1676037725
transform 1 0 25024 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_268
timestamp 1676037725
transform 1 0 25760 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_291
timestamp 1676037725
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1676037725
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_329
timestamp 1676037725
transform 1 0 31372 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_338
timestamp 1676037725
transform 1 0 32200 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_342
timestamp 1676037725
transform 1 0 32568 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_350
timestamp 1676037725
transform 1 0 33304 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1676037725
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_377
timestamp 1676037725
transform 1 0 35788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_381
timestamp 1676037725
transform 1 0 36156 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_387
timestamp 1676037725
transform 1 0 36708 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_399
timestamp 1676037725
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_412
timestamp 1676037725
transform 1 0 39008 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_445
timestamp 1676037725
transform 1 0 42044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_453
timestamp 1676037725
transform 1 0 42780 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_462
timestamp 1676037725
transform 1 0 43608 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_474
timestamp 1676037725
transform 1 0 44712 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1676037725
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1676037725
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1676037725
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1676037725
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1676037725
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1676037725
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1676037725
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1676037725
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1676037725
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_601
timestamp 1676037725
transform 1 0 56396 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_613
timestamp 1676037725
transform 1 0 57500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_623
timestamp 1676037725
transform 1 0 58420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_11
timestamp 1676037725
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_86
timestamp 1676037725
transform 1 0 9016 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_97
timestamp 1676037725
transform 1 0 10028 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_103
timestamp 1676037725
transform 1 0 10580 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_122
timestamp 1676037725
transform 1 0 12328 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_130
timestamp 1676037725
transform 1 0 13064 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_138
timestamp 1676037725
transform 1 0 13800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_187
timestamp 1676037725
transform 1 0 18308 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_200
timestamp 1676037725
transform 1 0 19504 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_212
timestamp 1676037725
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_221
timestamp 1676037725
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_236
timestamp 1676037725
transform 1 0 22816 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_248
timestamp 1676037725
transform 1 0 23920 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1676037725
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_303
timestamp 1676037725
transform 1 0 28980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_316
timestamp 1676037725
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_348
timestamp 1676037725
transform 1 0 33120 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_360
timestamp 1676037725
transform 1 0 34224 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_372
timestamp 1676037725
transform 1 0 35328 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_384
timestamp 1676037725
transform 1 0 36432 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_407
timestamp 1676037725
transform 1 0 38548 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_414
timestamp 1676037725
transform 1 0 39192 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_426
timestamp 1676037725
transform 1 0 40296 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_438
timestamp 1676037725
transform 1 0 41400 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_446
timestamp 1676037725
transform 1 0 42136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_455
timestamp 1676037725
transform 1 0 42964 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_475
timestamp 1676037725
transform 1 0 44804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_487
timestamp 1676037725
transform 1 0 45908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_499
timestamp 1676037725
transform 1 0 47012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1676037725
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1676037725
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1676037725
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1676037725
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1676037725
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1676037725
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1676037725
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1676037725
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1676037725
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1676037725
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1676037725
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_11
timestamp 1676037725
transform 1 0 2116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1676037725
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_108
timestamp 1676037725
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_129
timestamp 1676037725
transform 1 0 12972 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_163
timestamp 1676037725
transform 1 0 16100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_169
timestamp 1676037725
transform 1 0 16652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1676037725
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_204
timestamp 1676037725
transform 1 0 19872 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_212
timestamp 1676037725
transform 1 0 20608 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_220
timestamp 1676037725
transform 1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_227
timestamp 1676037725
transform 1 0 21988 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_235
timestamp 1676037725
transform 1 0 22724 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_243
timestamp 1676037725
transform 1 0 23460 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_266
timestamp 1676037725
transform 1 0 25576 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1676037725
transform 1 0 26312 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_279
timestamp 1676037725
transform 1 0 26772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_291
timestamp 1676037725
transform 1 0 27876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_299
timestamp 1676037725
transform 1 0 28612 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1676037725
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_328
timestamp 1676037725
transform 1 0 31280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_332
timestamp 1676037725
transform 1 0 31648 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_336
timestamp 1676037725
transform 1 0 32016 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1676037725
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1676037725
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_389
timestamp 1676037725
transform 1 0 36892 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_393
timestamp 1676037725
transform 1 0 37260 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_397
timestamp 1676037725
transform 1 0 37628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1676037725
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_440
timestamp 1676037725
transform 1 0 41584 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_444
timestamp 1676037725
transform 1 0 41952 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_451
timestamp 1676037725
transform 1 0 42596 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1676037725
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1676037725
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1676037725
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1676037725
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1676037725
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1676037725
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1676037725
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1676037725
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1676037725
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1676037725
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_613
timestamp 1676037725
transform 1 0 57500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_623
timestamp 1676037725
transform 1 0 58420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_11
timestamp 1676037725
transform 1 0 2116 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_23
timestamp 1676037725
transform 1 0 3220 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_35
timestamp 1676037725
transform 1 0 4324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1676037725
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1676037725
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1676037725
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_122
timestamp 1676037725
transform 1 0 12328 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_130
timestamp 1676037725
transform 1 0 13064 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_153
timestamp 1676037725
transform 1 0 15180 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_175
timestamp 1676037725
transform 1 0 17204 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1676037725
transform 1 0 18400 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_192
timestamp 1676037725
transform 1 0 18768 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_198
timestamp 1676037725
transform 1 0 19320 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_206
timestamp 1676037725
transform 1 0 20056 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1676037725
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_242
timestamp 1676037725
transform 1 0 23368 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_258
timestamp 1676037725
transform 1 0 24840 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_262
timestamp 1676037725
transform 1 0 25208 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_272
timestamp 1676037725
transform 1 0 26128 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_292
timestamp 1676037725
transform 1 0 27968 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_296
timestamp 1676037725
transform 1 0 28336 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_313
timestamp 1676037725
transform 1 0 29900 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_326
timestamp 1676037725
transform 1 0 31096 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1676037725
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_358
timestamp 1676037725
transform 1 0 34040 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_378
timestamp 1676037725
transform 1 0 35880 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1676037725
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_414
timestamp 1676037725
transform 1 0 39192 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_426
timestamp 1676037725
transform 1 0 40296 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_434
timestamp 1676037725
transform 1 0 41032 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_443
timestamp 1676037725
transform 1 0 41860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_453
timestamp 1676037725
transform 1 0 42780 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_460
timestamp 1676037725
transform 1 0 43424 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_472
timestamp 1676037725
transform 1 0 44528 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_484
timestamp 1676037725
transform 1 0 45632 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_496
timestamp 1676037725
transform 1 0 46736 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_516
timestamp 1676037725
transform 1 0 48576 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_528
timestamp 1676037725
transform 1 0 49680 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_540
timestamp 1676037725
transform 1 0 50784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_552
timestamp 1676037725
transform 1 0 51888 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1676037725
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1676037725
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1676037725
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1676037725
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1676037725
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1676037725
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1676037725
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1676037725
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_101
timestamp 1676037725
transform 1 0 10396 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_107
timestamp 1676037725
transform 1 0 10948 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1676037725
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_129
timestamp 1676037725
transform 1 0 12972 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1676037725
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_147
timestamp 1676037725
transform 1 0 14628 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_158
timestamp 1676037725
transform 1 0 15640 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_162
timestamp 1676037725
transform 1 0 16008 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_167
timestamp 1676037725
transform 1 0 16468 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_175
timestamp 1676037725
transform 1 0 17204 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_183
timestamp 1676037725
transform 1 0 17940 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1676037725
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_206
timestamp 1676037725
transform 1 0 20056 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_214
timestamp 1676037725
transform 1 0 20792 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_226
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_234
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_243
timestamp 1676037725
transform 1 0 23460 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_272
timestamp 1676037725
transform 1 0 26128 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_281
timestamp 1676037725
transform 1 0 26956 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_303
timestamp 1676037725
transform 1 0 28980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1676037725
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1676037725
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1676037725
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_376
timestamp 1676037725
transform 1 0 35696 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_384
timestamp 1676037725
transform 1 0 36432 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1676037725
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1676037725
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1676037725
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_442
timestamp 1676037725
transform 1 0 41768 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_454
timestamp 1676037725
transform 1 0 42872 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_466
timestamp 1676037725
transform 1 0 43976 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_474
timestamp 1676037725
transform 1 0 44712 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_517
timestamp 1676037725
transform 1 0 48668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_529
timestamp 1676037725
transform 1 0 49772 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1676037725
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_545
timestamp 1676037725
transform 1 0 51244 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_564
timestamp 1676037725
transform 1 0 52992 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_576
timestamp 1676037725
transform 1 0 54096 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1676037725
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1676037725
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_613
timestamp 1676037725
transform 1 0 57500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_623
timestamp 1676037725
transform 1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1676037725
transform 1 0 2116 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_99
timestamp 1676037725
transform 1 0 10212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_119
timestamp 1676037725
transform 1 0 12052 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_127
timestamp 1676037725
transform 1 0 12788 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_142
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_154
timestamp 1676037725
transform 1 0 15272 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_158
timestamp 1676037725
transform 1 0 15640 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1676037725
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_189
timestamp 1676037725
transform 1 0 18492 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_201
timestamp 1676037725
transform 1 0 19596 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_213
timestamp 1676037725
transform 1 0 20700 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1676037725
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_231
timestamp 1676037725
transform 1 0 22356 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_244
timestamp 1676037725
transform 1 0 23552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_252
timestamp 1676037725
transform 1 0 24288 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_266
timestamp 1676037725
transform 1 0 25576 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1676037725
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_292
timestamp 1676037725
transform 1 0 27968 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_313
timestamp 1676037725
transform 1 0 29900 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_325
timestamp 1676037725
transform 1 0 31004 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1676037725
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_347
timestamp 1676037725
transform 1 0 33028 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_359
timestamp 1676037725
transform 1 0 34132 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_371
timestamp 1676037725
transform 1 0 35236 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_383
timestamp 1676037725
transform 1 0 36340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_402
timestamp 1676037725
transform 1 0 38088 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_413
timestamp 1676037725
transform 1 0 39100 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_425
timestamp 1676037725
transform 1 0 40204 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_431
timestamp 1676037725
transform 1 0 40756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_446
timestamp 1676037725
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_458
timestamp 1676037725
transform 1 0 43240 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_466
timestamp 1676037725
transform 1 0 43976 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_488
timestamp 1676037725
transform 1 0 46000 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_501
timestamp 1676037725
transform 1 0 47196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_524
timestamp 1676037725
transform 1 0 49312 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_536
timestamp 1676037725
transform 1 0 50416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_541
timestamp 1676037725
transform 1 0 50876 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_550
timestamp 1676037725
transform 1 0 51704 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_558
timestamp 1676037725
transform 1 0 52440 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_561
timestamp 1676037725
transform 1 0 52716 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_566
timestamp 1676037725
transform 1 0 53176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_570
timestamp 1676037725
transform 1 0 53544 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_578
timestamp 1676037725
transform 1 0 54280 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_590
timestamp 1676037725
transform 1 0 55384 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_602
timestamp 1676037725
transform 1 0 56488 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_614
timestamp 1676037725
transform 1 0 57592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1676037725
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_11
timestamp 1676037725
transform 1 0 2116 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1676037725
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_125
timestamp 1676037725
transform 1 0 12604 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_161
timestamp 1676037725
transform 1 0 15916 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_167
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1676037725
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_203
timestamp 1676037725
transform 1 0 19780 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1676037725
transform 1 0 20424 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_230
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_237
timestamp 1676037725
transform 1 0 22908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1676037725
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_269
timestamp 1676037725
transform 1 0 25852 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_286
timestamp 1676037725
transform 1 0 27416 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_290
timestamp 1676037725
transform 1 0 27784 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1676037725
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_342
timestamp 1676037725
transform 1 0 32568 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1676037725
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_377
timestamp 1676037725
transform 1 0 35788 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_381
timestamp 1676037725
transform 1 0 36156 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_391
timestamp 1676037725
transform 1 0 37076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_411
timestamp 1676037725
transform 1 0 38916 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1676037725
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_427
timestamp 1676037725
transform 1 0 40388 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_435
timestamp 1676037725
transform 1 0 41124 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_446
timestamp 1676037725
transform 1 0 42136 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_458
timestamp 1676037725
transform 1 0 43240 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_470
timestamp 1676037725
transform 1 0 44344 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_496
timestamp 1676037725
transform 1 0 46736 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_508
timestamp 1676037725
transform 1 0 47840 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_520
timestamp 1676037725
transform 1 0 48944 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1676037725
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_545
timestamp 1676037725
transform 1 0 51244 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_552
timestamp 1676037725
transform 1 0 51888 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_560
timestamp 1676037725
transform 1 0 52624 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_568
timestamp 1676037725
transform 1 0 53360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_586
timestamp 1676037725
transform 1 0 55016 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1676037725
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_601
timestamp 1676037725
transform 1 0 56396 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_613
timestamp 1676037725
transform 1 0 57500 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_623
timestamp 1676037725
transform 1 0 58420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1676037725
transform 1 0 2116 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1676037725
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1676037725
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1676037725
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_153
timestamp 1676037725
transform 1 0 15180 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_157
timestamp 1676037725
transform 1 0 15548 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_177
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_185
timestamp 1676037725
transform 1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp 1676037725
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_194
timestamp 1676037725
transform 1 0 18952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_202
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_207
timestamp 1676037725
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_211
timestamp 1676037725
transform 1 0 20516 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_231
timestamp 1676037725
transform 1 0 22356 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_243
timestamp 1676037725
transform 1 0 23460 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_255
timestamp 1676037725
transform 1 0 24564 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_265
timestamp 1676037725
transform 1 0 25484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_277
timestamp 1676037725
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_289
timestamp 1676037725
transform 1 0 27692 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_299
timestamp 1676037725
transform 1 0 28612 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_311
timestamp 1676037725
transform 1 0 29716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_323
timestamp 1676037725
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1676037725
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_346
timestamp 1676037725
transform 1 0 32936 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_352
timestamp 1676037725
transform 1 0 33488 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_369
timestamp 1676037725
transform 1 0 35052 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_381
timestamp 1676037725
transform 1 0 36156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1676037725
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_401
timestamp 1676037725
transform 1 0 37996 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_413
timestamp 1676037725
transform 1 0 39100 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_425
timestamp 1676037725
transform 1 0 40204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_438
timestamp 1676037725
transform 1 0 41400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1676037725
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1676037725
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_541
timestamp 1676037725
transform 1 0 50876 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_552
timestamp 1676037725
transform 1 0 51888 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1676037725
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_573
timestamp 1676037725
transform 1 0 53820 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_579
timestamp 1676037725
transform 1 0 54372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_592
timestamp 1676037725
transform 1 0 55568 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_601
timestamp 1676037725
transform 1 0 56396 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_607
timestamp 1676037725
transform 1 0 56948 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_614
timestamp 1676037725
transform 1 0 57592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1676037725
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_11
timestamp 1676037725
transform 1 0 2116 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1676037725
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_63
timestamp 1676037725
transform 1 0 6900 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_91
timestamp 1676037725
transform 1 0 9476 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_98
timestamp 1676037725
transform 1 0 10120 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_110
timestamp 1676037725
transform 1 0 11224 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_122
timestamp 1676037725
transform 1 0 12328 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_134
timestamp 1676037725
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_147
timestamp 1676037725
transform 1 0 14628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_151
timestamp 1676037725
transform 1 0 14996 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_156
timestamp 1676037725
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_164
timestamp 1676037725
transform 1 0 16192 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_172
timestamp 1676037725
transform 1 0 16928 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_184
timestamp 1676037725
transform 1 0 18032 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1676037725
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_202
timestamp 1676037725
transform 1 0 19688 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_210
timestamp 1676037725
transform 1 0 20424 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_219
timestamp 1676037725
transform 1 0 21252 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_231
timestamp 1676037725
transform 1 0 22356 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_243
timestamp 1676037725
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1676037725
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_262
timestamp 1676037725
transform 1 0 25208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_271
timestamp 1676037725
transform 1 0 26036 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_279
timestamp 1676037725
transform 1 0 26772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_289
timestamp 1676037725
transform 1 0 27692 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_293
timestamp 1676037725
transform 1 0 28060 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1676037725
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_320
timestamp 1676037725
transform 1 0 30544 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_337
timestamp 1676037725
transform 1 0 32108 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_346
timestamp 1676037725
transform 1 0 32936 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_350
timestamp 1676037725
transform 1 0 33304 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_360
timestamp 1676037725
transform 1 0 34224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_373
timestamp 1676037725
transform 1 0 35420 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_385
timestamp 1676037725
transform 1 0 36524 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_397
timestamp 1676037725
transform 1 0 37628 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 1676037725
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_441
timestamp 1676037725
transform 1 0 41676 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_453
timestamp 1676037725
transform 1 0 42780 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_465
timestamp 1676037725
transform 1 0 43884 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_473
timestamp 1676037725
transform 1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_516
timestamp 1676037725
transform 1 0 48576 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_528
timestamp 1676037725
transform 1 0 49680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_533
timestamp 1676037725
transform 1 0 50140 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_537
timestamp 1676037725
transform 1 0 50508 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_545
timestamp 1676037725
transform 1 0 51244 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_565
timestamp 1676037725
transform 1 0 53084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_577
timestamp 1676037725
transform 1 0 54188 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_585
timestamp 1676037725
transform 1 0 54924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_589
timestamp 1676037725
transform 1 0 55292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_597
timestamp 1676037725
transform 1 0 56028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_605
timestamp 1676037725
transform 1 0 56764 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_622
timestamp 1676037725
transform 1 0 58328 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_47
timestamp 1676037725
transform 1 0 5428 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1676037725
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_66
timestamp 1676037725
transform 1 0 7176 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_74
timestamp 1676037725
transform 1 0 7912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1676037725
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_104
timestamp 1676037725
transform 1 0 10672 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp 1676037725
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_122
timestamp 1676037725
transform 1 0 12328 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_134
timestamp 1676037725
transform 1 0 13432 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_142
timestamp 1676037725
transform 1 0 14168 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_153
timestamp 1676037725
transform 1 0 15180 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_158
timestamp 1676037725
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1676037725
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_191
timestamp 1676037725
transform 1 0 18676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_197
timestamp 1676037725
transform 1 0 19228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_203
timestamp 1676037725
transform 1 0 19780 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_209
timestamp 1676037725
transform 1 0 20332 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_214
timestamp 1676037725
transform 1 0 20792 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_231
timestamp 1676037725
transform 1 0 22356 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_244
timestamp 1676037725
transform 1 0 23552 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_256
timestamp 1676037725
transform 1 0 24656 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_268
timestamp 1676037725
transform 1 0 25760 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1676037725
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1676037725
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_326
timestamp 1676037725
transform 1 0 31096 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1676037725
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_346
timestamp 1676037725
transform 1 0 32936 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_354
timestamp 1676037725
transform 1 0 33672 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_366
timestamp 1676037725
transform 1 0 34776 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_378
timestamp 1676037725
transform 1 0 35880 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1676037725
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_405
timestamp 1676037725
transform 1 0 38364 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_409
timestamp 1676037725
transform 1 0 38732 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1676037725
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1676037725
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1676037725
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_458
timestamp 1676037725
transform 1 0 43240 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_470
timestamp 1676037725
transform 1 0 44344 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_482
timestamp 1676037725
transform 1 0 45448 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_486
timestamp 1676037725
transform 1 0 45816 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_494
timestamp 1676037725
transform 1 0 46552 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_502
timestamp 1676037725
transform 1 0 47288 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_534
timestamp 1676037725
transform 1 0 50232 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_546
timestamp 1676037725
transform 1 0 51336 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_558
timestamp 1676037725
transform 1 0 52440 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1676037725
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_573
timestamp 1676037725
transform 1 0 53820 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_588
timestamp 1676037725
transform 1 0 55200 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_594
timestamp 1676037725
transform 1 0 55752 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_611
timestamp 1676037725
transform 1 0 57316 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1676037725
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1676037725
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_11
timestamp 1676037725
transform 1 0 2116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1676037725
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_45
timestamp 1676037725
transform 1 0 5244 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_50
timestamp 1676037725
transform 1 0 5704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_71
timestamp 1676037725
transform 1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_94
timestamp 1676037725
transform 1 0 9752 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_105
timestamp 1676037725
transform 1 0 10764 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_111
timestamp 1676037725
transform 1 0 11316 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_115
timestamp 1676037725
transform 1 0 11684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1676037725
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_150
timestamp 1676037725
transform 1 0 14904 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_162
timestamp 1676037725
transform 1 0 16008 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_178
timestamp 1676037725
transform 1 0 17480 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_186
timestamp 1676037725
transform 1 0 18216 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_207
timestamp 1676037725
transform 1 0 20148 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_215
timestamp 1676037725
transform 1 0 20884 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_225
timestamp 1676037725
transform 1 0 21804 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_233
timestamp 1676037725
transform 1 0 22540 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_241
timestamp 1676037725
transform 1 0 23276 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_245
timestamp 1676037725
transform 1 0 23644 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_272
timestamp 1676037725
transform 1 0 26128 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_292
timestamp 1676037725
transform 1 0 27968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1676037725
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_320
timestamp 1676037725
transform 1 0 30544 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_333
timestamp 1676037725
transform 1 0 31740 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_339
timestamp 1676037725
transform 1 0 32292 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_344
timestamp 1676037725
transform 1 0 32752 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_356
timestamp 1676037725
transform 1 0 33856 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_385
timestamp 1676037725
transform 1 0 36524 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_396
timestamp 1676037725
transform 1 0 37536 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_408
timestamp 1676037725
transform 1 0 38640 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_414
timestamp 1676037725
transform 1 0 39192 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_438
timestamp 1676037725
transform 1 0 41400 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_458
timestamp 1676037725
transform 1 0 43240 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_467
timestamp 1676037725
transform 1 0 44068 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_485
timestamp 1676037725
transform 1 0 45724 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_496
timestamp 1676037725
transform 1 0 46736 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_506
timestamp 1676037725
transform 1 0 47656 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_514
timestamp 1676037725
transform 1 0 48392 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_520
timestamp 1676037725
transform 1 0 48944 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1676037725
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1676037725
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1676037725
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1676037725
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1676037725
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1676037725
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_589
timestamp 1676037725
transform 1 0 55292 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_596
timestamp 1676037725
transform 1 0 55936 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_604
timestamp 1676037725
transform 1 0 56672 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_613
timestamp 1676037725
transform 1 0 57500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_623
timestamp 1676037725
transform 1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_11
timestamp 1676037725
transform 1 0 2116 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_23
timestamp 1676037725
transform 1 0 3220 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_35
timestamp 1676037725
transform 1 0 4324 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 1676037725
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_61
timestamp 1676037725
transform 1 0 6716 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_100
timestamp 1676037725
transform 1 0 10304 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_119
timestamp 1676037725
transform 1 0 12052 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_140
timestamp 1676037725
transform 1 0 13984 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_189
timestamp 1676037725
transform 1 0 18492 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_201
timestamp 1676037725
transform 1 0 19596 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_231
timestamp 1676037725
transform 1 0 22356 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_239
timestamp 1676037725
transform 1 0 23092 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_259
timestamp 1676037725
transform 1 0 24932 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_265
timestamp 1676037725
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_270
timestamp 1676037725
transform 1 0 25944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_285
timestamp 1676037725
transform 1 0 27324 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_303
timestamp 1676037725
transform 1 0 28980 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_315
timestamp 1676037725
transform 1 0 30084 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1676037725
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_349
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_362
timestamp 1676037725
transform 1 0 34408 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_374
timestamp 1676037725
transform 1 0 35512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1676037725
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1676037725
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1676037725
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1676037725
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_453
timestamp 1676037725
transform 1 0 42780 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_470
timestamp 1676037725
transform 1 0 44344 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_499
timestamp 1676037725
transform 1 0 47012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_513
timestamp 1676037725
transform 1 0 48300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_536
timestamp 1676037725
transform 1 0 50416 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_542
timestamp 1676037725
transform 1 0 50968 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_550
timestamp 1676037725
transform 1 0 51704 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_558
timestamp 1676037725
transform 1 0 52440 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1676037725
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_573
timestamp 1676037725
transform 1 0 53820 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_586
timestamp 1676037725
transform 1 0 55016 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_598
timestamp 1676037725
transform 1 0 56120 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_610
timestamp 1676037725
transform 1 0 57224 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1676037725
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_11
timestamp 1676037725
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1676037725
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_61
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_68
timestamp 1676037725
transform 1 0 7360 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1676037725
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_91
timestamp 1676037725
transform 1 0 9476 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1676037725
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_107
timestamp 1676037725
transform 1 0 10948 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_118
timestamp 1676037725
transform 1 0 11960 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_147
timestamp 1676037725
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1676037725
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_208
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_212
timestamp 1676037725
transform 1 0 20608 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_229
timestamp 1676037725
transform 1 0 22172 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_237
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_264
timestamp 1676037725
transform 1 0 25392 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_273
timestamp 1676037725
transform 1 0 26220 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_284
timestamp 1676037725
transform 1 0 27232 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_297
timestamp 1676037725
transform 1 0 28428 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1676037725
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_338
timestamp 1676037725
transform 1 0 32200 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_344
timestamp 1676037725
transform 1 0 32752 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_362
timestamp 1676037725
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_394
timestamp 1676037725
transform 1 0 37352 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_407
timestamp 1676037725
transform 1 0 38548 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1676037725
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_427
timestamp 1676037725
transform 1 0 40388 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_433
timestamp 1676037725
transform 1 0 40940 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_454
timestamp 1676037725
transform 1 0 42872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_474
timestamp 1676037725
transform 1 0 44712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_486
timestamp 1676037725
transform 1 0 45816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_507
timestamp 1676037725
transform 1 0 47748 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_516
timestamp 1676037725
transform 1 0 48576 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_528
timestamp 1676037725
transform 1 0 49680 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_533
timestamp 1676037725
transform 1 0 50140 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_553
timestamp 1676037725
transform 1 0 51980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_574
timestamp 1676037725
transform 1 0 53912 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_585
timestamp 1676037725
transform 1 0 54924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_589
timestamp 1676037725
transform 1 0 55292 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_598
timestamp 1676037725
transform 1 0 56120 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_622
timestamp 1676037725
transform 1 0 58328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_11
timestamp 1676037725
transform 1 0 2116 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_23
timestamp 1676037725
transform 1 0 3220 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_35
timestamp 1676037725
transform 1 0 4324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_47
timestamp 1676037725
transform 1 0 5428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_79
timestamp 1676037725
transform 1 0 8372 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_91
timestamp 1676037725
transform 1 0 9476 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_103
timestamp 1676037725
transform 1 0 10580 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_117
timestamp 1676037725
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_122
timestamp 1676037725
transform 1 0 12328 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_126
timestamp 1676037725
transform 1 0 12696 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_134
timestamp 1676037725
transform 1 0 13432 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_144
timestamp 1676037725
transform 1 0 14352 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_152
timestamp 1676037725
transform 1 0 15088 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_158
timestamp 1676037725
transform 1 0 15640 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1676037725
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_190
timestamp 1676037725
transform 1 0 18584 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_199
timestamp 1676037725
transform 1 0 19412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_208
timestamp 1676037725
transform 1 0 20240 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1676037725
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_236
timestamp 1676037725
transform 1 0 22816 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_244
timestamp 1676037725
transform 1 0 23552 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_262
timestamp 1676037725
transform 1 0 25208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1676037725
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1676037725
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_300
timestamp 1676037725
transform 1 0 28704 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_304
timestamp 1676037725
transform 1 0 29072 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_309
timestamp 1676037725
transform 1 0 29532 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1676037725
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_330
timestamp 1676037725
transform 1 0 31464 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_354
timestamp 1676037725
transform 1 0 33672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_367
timestamp 1676037725
transform 1 0 34868 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1676037725
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_400
timestamp 1676037725
transform 1 0 37904 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_425
timestamp 1676037725
transform 1 0 40204 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_437
timestamp 1676037725
transform 1 0 41308 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_443
timestamp 1676037725
transform 1 0 41860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_459
timestamp 1676037725
transform 1 0 43332 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_471
timestamp 1676037725
transform 1 0 44436 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_483
timestamp 1676037725
transform 1 0 45540 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_493
timestamp 1676037725
transform 1 0 46460 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_501
timestamp 1676037725
transform 1 0 47196 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_511
timestamp 1676037725
transform 1 0 48116 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_529
timestamp 1676037725
transform 1 0 49772 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_533
timestamp 1676037725
transform 1 0 50140 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_539
timestamp 1676037725
transform 1 0 50692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_552
timestamp 1676037725
transform 1 0 51888 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_561
timestamp 1676037725
transform 1 0 52716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_581
timestamp 1676037725
transform 1 0 54556 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_601
timestamp 1676037725
transform 1 0 56396 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_613
timestamp 1676037725
transform 1 0 57500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1676037725
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_117
timestamp 1676037725
transform 1 0 11868 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_123
timestamp 1676037725
transform 1 0 12420 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1676037725
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_147
timestamp 1676037725
transform 1 0 14628 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_156
timestamp 1676037725
transform 1 0 15456 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_164
timestamp 1676037725
transform 1 0 16192 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_172
timestamp 1676037725
transform 1 0 16928 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_180
timestamp 1676037725
transform 1 0 17664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_190
timestamp 1676037725
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_203
timestamp 1676037725
transform 1 0 19780 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_211
timestamp 1676037725
transform 1 0 20516 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_219
timestamp 1676037725
transform 1 0 21252 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_227
timestamp 1676037725
transform 1 0 21988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_239
timestamp 1676037725
transform 1 0 23092 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_245
timestamp 1676037725
transform 1 0 23644 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_260
timestamp 1676037725
transform 1 0 25024 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_268
timestamp 1676037725
transform 1 0 25760 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_273
timestamp 1676037725
transform 1 0 26220 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_280
timestamp 1676037725
transform 1 0 26864 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_284
timestamp 1676037725
transform 1 0 27232 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_295
timestamp 1676037725
transform 1 0 28244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1676037725
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_317
timestamp 1676037725
transform 1 0 30268 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_325
timestamp 1676037725
transform 1 0 31004 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1676037725
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1676037725
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1676037725
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1676037725
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_370
timestamp 1676037725
transform 1 0 35144 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_374
timestamp 1676037725
transform 1 0 35512 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_385
timestamp 1676037725
transform 1 0 36524 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_393
timestamp 1676037725
transform 1 0 37260 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_410
timestamp 1676037725
transform 1 0 38824 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_418
timestamp 1676037725
transform 1 0 39560 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_433
timestamp 1676037725
transform 1 0 40940 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_450
timestamp 1676037725
transform 1 0 42504 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_464
timestamp 1676037725
transform 1 0 43792 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_511
timestamp 1676037725
transform 1 0 48116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_523
timestamp 1676037725
transform 1 0 49220 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1676037725
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1676037725
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1676037725
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_557
timestamp 1676037725
transform 1 0 52348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_560
timestamp 1676037725
transform 1 0 52624 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_569
timestamp 1676037725
transform 1 0 53452 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_578
timestamp 1676037725
transform 1 0 54280 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_586
timestamp 1676037725
transform 1 0 55016 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_589
timestamp 1676037725
transform 1 0 55292 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_600
timestamp 1676037725
transform 1 0 56304 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_612
timestamp 1676037725
transform 1 0 57408 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_616
timestamp 1676037725
transform 1 0 57776 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_623
timestamp 1676037725
transform 1 0 58420 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1676037725
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1676037725
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1676037725
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1676037725
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1676037725
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_101
timestamp 1676037725
transform 1 0 10396 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1676037725
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_178
timestamp 1676037725
transform 1 0 17480 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_186
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_191
timestamp 1676037725
transform 1 0 18676 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_199
timestamp 1676037725
transform 1 0 19412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_206
timestamp 1676037725
transform 1 0 20056 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_212
timestamp 1676037725
transform 1 0 20608 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1676037725
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_233
timestamp 1676037725
transform 1 0 22540 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_248
timestamp 1676037725
transform 1 0 23920 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_256
timestamp 1676037725
transform 1 0 24656 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_268
timestamp 1676037725
transform 1 0 25760 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_274
timestamp 1676037725
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_293
timestamp 1676037725
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_303
timestamp 1676037725
transform 1 0 28980 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_315
timestamp 1676037725
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1676037725
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1676037725
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1676037725
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1676037725
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1676037725
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_414
timestamp 1676037725
transform 1 0 39192 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_426
timestamp 1676037725
transform 1 0 40296 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_438
timestamp 1676037725
transform 1 0 41400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1676037725
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_456
timestamp 1676037725
transform 1 0 43056 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_468
timestamp 1676037725
transform 1 0 44160 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_480
timestamp 1676037725
transform 1 0 45264 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_492
timestamp 1676037725
transform 1 0 46368 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1676037725
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1676037725
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1676037725
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1676037725
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1676037725
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1676037725
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1676037725
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1676037725
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1676037725
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1676037725
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1676037725
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_617
timestamp 1676037725
transform 1 0 57868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_623
timestamp 1676037725
transform 1 0 58420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_11
timestamp 1676037725
transform 1 0 2116 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1676037725
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_89
timestamp 1676037725
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_95
timestamp 1676037725
transform 1 0 9844 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_107
timestamp 1676037725
transform 1 0 10948 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_119
timestamp 1676037725
transform 1 0 12052 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_131
timestamp 1676037725
transform 1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_165
timestamp 1676037725
transform 1 0 16284 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_177
timestamp 1676037725
transform 1 0 17388 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_185
timestamp 1676037725
transform 1 0 18124 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1676037725
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1676037725
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1676037725
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1676037725
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1676037725
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1676037725
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1676037725
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1676037725
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1676037725
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1676037725
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1676037725
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1676037725
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1676037725
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1676037725
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1676037725
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1676037725
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1676037725
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1676037725
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1676037725
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1676037725
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1676037725
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1676037725
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1676037725
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1676037725
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1676037725
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1676037725
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1676037725
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1676037725
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_613
timestamp 1676037725
transform 1 0 57500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_623
timestamp 1676037725
transform 1 0 58420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_11
timestamp 1676037725
transform 1 0 2116 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_23
timestamp 1676037725
transform 1 0 3220 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_35
timestamp 1676037725
transform 1 0 4324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_47
timestamp 1676037725
transform 1 0 5428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1676037725
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1676037725
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_178
timestamp 1676037725
transform 1 0 17480 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_190
timestamp 1676037725
transform 1 0 18584 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_202
timestamp 1676037725
transform 1 0 19688 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_214
timestamp 1676037725
transform 1 0 20792 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1676037725
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1676037725
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1676037725
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1676037725
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1676037725
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1676037725
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1676037725
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1676037725
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1676037725
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1676037725
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1676037725
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1676037725
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1676037725
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1676037725
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1676037725
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1676037725
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1676037725
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1676037725
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1676037725
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1676037725
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1676037725
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1676037725
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1676037725
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1676037725
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1676037725
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1676037725
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1676037725
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_617
timestamp 1676037725
transform 1 0 57868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1676037725
transform 1 0 58420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_11
timestamp 1676037725
transform 1 0 2116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 1676037725
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_105
timestamp 1676037725
transform 1 0 10764 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_111
timestamp 1676037725
transform 1 0 11316 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_117
timestamp 1676037725
transform 1 0 11868 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_123
timestamp 1676037725
transform 1 0 12420 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1676037725
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1676037725
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1676037725
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1676037725
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1676037725
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1676037725
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1676037725
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1676037725
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1676037725
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1676037725
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1676037725
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1676037725
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1676037725
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1676037725
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1676037725
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1676037725
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1676037725
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1676037725
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1676037725
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1676037725
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1676037725
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1676037725
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1676037725
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1676037725
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1676037725
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1676037725
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1676037725
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1676037725
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1676037725
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1676037725
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1676037725
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_613
timestamp 1676037725
transform 1 0 57500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_623
timestamp 1676037725
transform 1 0 58420 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1676037725
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1676037725
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_119
timestamp 1676037725
transform 1 0 12052 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_129
timestamp 1676037725
transform 1 0 12972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_141
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_153
timestamp 1676037725
transform 1 0 15180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1676037725
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1676037725
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1676037725
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1676037725
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1676037725
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1676037725
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1676037725
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1676037725
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1676037725
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1676037725
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1676037725
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1676037725
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1676037725
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1676037725
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1676037725
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1676037725
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1676037725
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1676037725
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1676037725
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1676037725
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1676037725
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1676037725
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1676037725
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1676037725
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1676037725
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1676037725
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1676037725
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1676037725
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1676037725
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1676037725
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1676037725
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1676037725
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_11
timestamp 1676037725
transform 1 0 2116 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_22
timestamp 1676037725
transform 1 0 3128 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1676037725
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1676037725
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1676037725
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1676037725
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1676037725
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1676037725
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1676037725
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1676037725
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1676037725
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1676037725
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1676037725
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1676037725
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1676037725
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1676037725
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1676037725
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1676037725
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1676037725
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1676037725
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1676037725
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1676037725
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1676037725
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1676037725
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1676037725
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1676037725
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1676037725
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1676037725
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1676037725
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1676037725
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1676037725
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1676037725
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1676037725
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1676037725
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_11
timestamp 1676037725
transform 1 0 2116 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_23
timestamp 1676037725
transform 1 0 3220 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_35
timestamp 1676037725
transform 1 0 4324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1676037725
transform 1 0 5428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1676037725
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1676037725
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1676037725
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1676037725
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1676037725
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1676037725
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1676037725
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1676037725
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1676037725
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1676037725
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1676037725
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1676037725
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1676037725
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1676037725
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1676037725
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1676037725
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1676037725
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1676037725
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1676037725
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1676037725
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1676037725
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1676037725
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1676037725
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1676037725
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1676037725
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1676037725
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1676037725
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1676037725
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1676037725
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1676037725
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1676037725
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1676037725
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1676037725
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1676037725
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1676037725
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1676037725
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_617
timestamp 1676037725
transform 1 0 57868 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_623
timestamp 1676037725
transform 1 0 58420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1676037725
transform 1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1676037725
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1676037725
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1676037725
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1676037725
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1676037725
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1676037725
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1676037725
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1676037725
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1676037725
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1676037725
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1676037725
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1676037725
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1676037725
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1676037725
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1676037725
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1676037725
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1676037725
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1676037725
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1676037725
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1676037725
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1676037725
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1676037725
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1676037725
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1676037725
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1676037725
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1676037725
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1676037725
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1676037725
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1676037725
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1676037725
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1676037725
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1676037725
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1676037725
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1676037725
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1676037725
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1676037725
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1676037725
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1676037725
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1676037725
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1676037725
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1676037725
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_613
timestamp 1676037725
transform 1 0 57500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_623
timestamp 1676037725
transform 1 0 58420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_11
timestamp 1676037725
transform 1 0 2116 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_23
timestamp 1676037725
transform 1 0 3220 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_35
timestamp 1676037725
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1676037725
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_101
timestamp 1676037725
transform 1 0 10396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_109
timestamp 1676037725
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1676037725
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1676037725
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1676037725
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1676037725
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1676037725
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1676037725
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1676037725
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1676037725
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1676037725
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1676037725
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1676037725
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1676037725
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1676037725
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1676037725
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1676037725
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1676037725
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1676037725
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1676037725
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1676037725
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1676037725
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1676037725
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1676037725
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1676037725
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1676037725
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1676037725
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1676037725
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1676037725
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1676037725
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1676037725
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1676037725
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1676037725
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1676037725
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1676037725
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1676037725
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1676037725
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1676037725
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1676037725
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_617
timestamp 1676037725
transform 1 0 57868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_623
timestamp 1676037725
transform 1 0 58420 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1676037725
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1676037725
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1676037725
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_233
timestamp 1676037725
transform 1 0 22540 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1676037725
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1676037725
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1676037725
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1676037725
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1676037725
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1676037725
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1676037725
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1676037725
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1676037725
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1676037725
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1676037725
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1676037725
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1676037725
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1676037725
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1676037725
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1676037725
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1676037725
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1676037725
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1676037725
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1676037725
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1676037725
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1676037725
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1676037725
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1676037725
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1676037725
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1676037725
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1676037725
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1676037725
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1676037725
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1676037725
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1676037725
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1676037725
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1676037725
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1676037725
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1676037725
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_613
timestamp 1676037725
transform 1 0 57500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_623
timestamp 1676037725
transform 1 0 58420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_11
timestamp 1676037725
transform 1 0 2116 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_20
timestamp 1676037725
transform 1 0 2944 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_32
timestamp 1676037725
transform 1 0 4048 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_44
timestamp 1676037725
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1676037725
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1676037725
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1676037725
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1676037725
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_233
timestamp 1676037725
transform 1 0 22540 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_244
timestamp 1676037725
transform 1 0 23552 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_256
timestamp 1676037725
transform 1 0 24656 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_268
timestamp 1676037725
transform 1 0 25760 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1676037725
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1676037725
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1676037725
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1676037725
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1676037725
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1676037725
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1676037725
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1676037725
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1676037725
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1676037725
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1676037725
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1676037725
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1676037725
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1676037725
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1676037725
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1676037725
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1676037725
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1676037725
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1676037725
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1676037725
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1676037725
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1676037725
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1676037725
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1676037725
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1676037725
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1676037725
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1676037725
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1676037725
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1676037725
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1676037725
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1676037725
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1676037725
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1676037725
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_11
timestamp 1676037725
transform 1 0 2116 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_23
timestamp 1676037725
transform 1 0 3220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1676037725
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1676037725
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1676037725
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1676037725
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1676037725
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1676037725
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1676037725
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1676037725
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1676037725
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1676037725
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1676037725
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1676037725
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1676037725
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1676037725
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1676037725
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1676037725
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1676037725
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1676037725
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1676037725
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1676037725
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1676037725
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1676037725
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1676037725
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1676037725
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1676037725
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1676037725
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1676037725
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1676037725
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1676037725
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1676037725
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1676037725
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1676037725
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1676037725
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1676037725
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1676037725
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1676037725
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1676037725
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_613
timestamp 1676037725
transform 1 0 57500 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_623
timestamp 1676037725
transform 1 0 58420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_11
timestamp 1676037725
transform 1 0 2116 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_23
timestamp 1676037725
transform 1 0 3220 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_35
timestamp 1676037725
transform 1 0 4324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_47
timestamp 1676037725
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1676037725
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1676037725
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1676037725
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1676037725
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1676037725
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1676037725
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1676037725
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1676037725
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1676037725
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1676037725
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1676037725
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1676037725
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1676037725
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1676037725
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1676037725
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1676037725
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1676037725
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1676037725
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1676037725
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1676037725
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1676037725
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1676037725
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1676037725
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1676037725
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1676037725
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1676037725
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1676037725
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1676037725
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1676037725
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1676037725
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1676037725
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1676037725
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1676037725
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1676037725
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1676037725
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1676037725
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1676037725
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1676037725
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1676037725
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1676037725
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1676037725
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1676037725
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_11
timestamp 1676037725
transform 1 0 2116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_20
timestamp 1676037725
transform 1 0 2944 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1676037725
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1676037725
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1676037725
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1676037725
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1676037725
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1676037725
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1676037725
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1676037725
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1676037725
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1676037725
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1676037725
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1676037725
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1676037725
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1676037725
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1676037725
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1676037725
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1676037725
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1676037725
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1676037725
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1676037725
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1676037725
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1676037725
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1676037725
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1676037725
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1676037725
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1676037725
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1676037725
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1676037725
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1676037725
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1676037725
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1676037725
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1676037725
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1676037725
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1676037725
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1676037725
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1676037725
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1676037725
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_613
timestamp 1676037725
transform 1 0 57500 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_623
timestamp 1676037725
transform 1 0 58420 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_89
timestamp 1676037725
transform 1 0 9292 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_95
timestamp 1676037725
transform 1 0 9844 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_107
timestamp 1676037725
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1676037725
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1676037725
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1676037725
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1676037725
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1676037725
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1676037725
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1676037725
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1676037725
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1676037725
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1676037725
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1676037725
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1676037725
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1676037725
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1676037725
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1676037725
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1676037725
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1676037725
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1676037725
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1676037725
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1676037725
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1676037725
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1676037725
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1676037725
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1676037725
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1676037725
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1676037725
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1676037725
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1676037725
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1676037725
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1676037725
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1676037725
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1676037725
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1676037725
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1676037725
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1676037725
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1676037725
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1676037725
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1676037725
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_11
timestamp 1676037725
transform 1 0 2116 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1676037725
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1676037725
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1676037725
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1676037725
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1676037725
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_242
timestamp 1676037725
transform 1 0 23368 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1676037725
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1676037725
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1676037725
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1676037725
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1676037725
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1676037725
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1676037725
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1676037725
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1676037725
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1676037725
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1676037725
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1676037725
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1676037725
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1676037725
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1676037725
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1676037725
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1676037725
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1676037725
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1676037725
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1676037725
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1676037725
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1676037725
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1676037725
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1676037725
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1676037725
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1676037725
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1676037725
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1676037725
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1676037725
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1676037725
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1676037725
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1676037725
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1676037725
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1676037725
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_601
timestamp 1676037725
transform 1 0 56396 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 1676037725
transform 1 0 57500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_623
timestamp 1676037725
transform 1 0 58420 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_11
timestamp 1676037725
transform 1 0 2116 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_23
timestamp 1676037725
transform 1 0 3220 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_35
timestamp 1676037725
transform 1 0 4324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_47
timestamp 1676037725
transform 1 0 5428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1676037725
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1676037725
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1676037725
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1676037725
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_189
timestamp 1676037725
transform 1 0 18492 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_200
timestamp 1676037725
transform 1 0 19504 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_212
timestamp 1676037725
transform 1 0 20608 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_234
timestamp 1676037725
transform 1 0 22632 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_238
timestamp 1676037725
transform 1 0 23000 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_248
timestamp 1676037725
transform 1 0 23920 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_260
timestamp 1676037725
transform 1 0 25024 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_272
timestamp 1676037725
transform 1 0 26128 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1676037725
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1676037725
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1676037725
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1676037725
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1676037725
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1676037725
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1676037725
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1676037725
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1676037725
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1676037725
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1676037725
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1676037725
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1676037725
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1676037725
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1676037725
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1676037725
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1676037725
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1676037725
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1676037725
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1676037725
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1676037725
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1676037725
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1676037725
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1676037725
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1676037725
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1676037725
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1676037725
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1676037725
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1676037725
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1676037725
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1676037725
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1676037725
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1676037725
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1676037725
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1676037725
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1676037725
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1676037725
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1676037725
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_208
timestamp 1676037725
transform 1 0 20240 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_220
timestamp 1676037725
transform 1 0 21344 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_232
timestamp 1676037725
transform 1 0 22448 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_243
timestamp 1676037725
transform 1 0 23460 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1676037725
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1676037725
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1676037725
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1676037725
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1676037725
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1676037725
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1676037725
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1676037725
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1676037725
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1676037725
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1676037725
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1676037725
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1676037725
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1676037725
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1676037725
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1676037725
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1676037725
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1676037725
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1676037725
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1676037725
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1676037725
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1676037725
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1676037725
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1676037725
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1676037725
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1676037725
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1676037725
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1676037725
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1676037725
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1676037725
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1676037725
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1676037725
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1676037725
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1676037725
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1676037725
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1676037725
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_9
timestamp 1676037725
transform 1 0 1932 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_21
timestamp 1676037725
transform 1 0 3036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1676037725
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1676037725
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1676037725
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1676037725
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1676037725
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1676037725
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1676037725
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1676037725
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_249
timestamp 1676037725
transform 1 0 24012 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_259
timestamp 1676037725
transform 1 0 24932 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_271
timestamp 1676037725
transform 1 0 26036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1676037725
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1676037725
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1676037725
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1676037725
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1676037725
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1676037725
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1676037725
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1676037725
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1676037725
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1676037725
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1676037725
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1676037725
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1676037725
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1676037725
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1676037725
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1676037725
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1676037725
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1676037725
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1676037725
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1676037725
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1676037725
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1676037725
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1676037725
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1676037725
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1676037725
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1676037725
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1676037725
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1676037725
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1676037725
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_617
timestamp 1676037725
transform 1 0 57868 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_623
timestamp 1676037725
transform 1 0 58420 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1676037725
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1676037725
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1676037725
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1676037725
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_233
timestamp 1676037725
transform 1 0 22540 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_236
timestamp 1676037725
transform 1 0 22816 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1676037725
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1676037725
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1676037725
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1676037725
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1676037725
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1676037725
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1676037725
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1676037725
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1676037725
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1676037725
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1676037725
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1676037725
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1676037725
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1676037725
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1676037725
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1676037725
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1676037725
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1676037725
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1676037725
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1676037725
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1676037725
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1676037725
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1676037725
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1676037725
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1676037725
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1676037725
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1676037725
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1676037725
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1676037725
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1676037725
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1676037725
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1676037725
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1676037725
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1676037725
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1676037725
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_613
timestamp 1676037725
transform 1 0 57500 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_623
timestamp 1676037725
transform 1 0 58420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1676037725
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1676037725
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1676037725
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1676037725
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1676037725
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1676037725
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1676037725
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1676037725
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1676037725
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1676037725
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1676037725
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1676037725
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1676037725
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_249
timestamp 1676037725
transform 1 0 24012 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_257
timestamp 1676037725
transform 1 0 24748 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_267
timestamp 1676037725
transform 1 0 25668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1676037725
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1676037725
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1676037725
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1676037725
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1676037725
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1676037725
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1676037725
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1676037725
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1676037725
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1676037725
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1676037725
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1676037725
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1676037725
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1676037725
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1676037725
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1676037725
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1676037725
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1676037725
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1676037725
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1676037725
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1676037725
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1676037725
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1676037725
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1676037725
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1676037725
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1676037725
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1676037725
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1676037725
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1676037725
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1676037725
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1676037725
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_9
timestamp 1676037725
transform 1 0 1932 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1676037725
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1676037725
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_221
timestamp 1676037725
transform 1 0 21436 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1676037725
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1676037725
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1676037725
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1676037725
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1676037725
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1676037725
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1676037725
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1676037725
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1676037725
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1676037725
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1676037725
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1676037725
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1676037725
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1676037725
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1676037725
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1676037725
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1676037725
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1676037725
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1676037725
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1676037725
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1676037725
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1676037725
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1676037725
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1676037725
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1676037725
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1676037725
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1676037725
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1676037725
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1676037725
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1676037725
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1676037725
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1676037725
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1676037725
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1676037725
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1676037725
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1676037725
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_601
timestamp 1676037725
transform 1 0 56396 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_613
timestamp 1676037725
transform 1 0 57500 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_623
timestamp 1676037725
transform 1 0 58420 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_9
timestamp 1676037725
transform 1 0 1932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1676037725
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1676037725
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1676037725
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1676037725
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_205
timestamp 1676037725
transform 1 0 19964 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_213
timestamp 1676037725
transform 1 0 20700 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1676037725
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_235
timestamp 1676037725
transform 1 0 22724 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_247
timestamp 1676037725
transform 1 0 23828 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_259
timestamp 1676037725
transform 1 0 24932 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_271
timestamp 1676037725
transform 1 0 26036 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1676037725
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1676037725
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1676037725
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1676037725
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1676037725
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1676037725
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1676037725
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_373
timestamp 1676037725
transform 1 0 35420 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1676037725
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1676037725
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1676037725
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1676037725
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1676037725
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1676037725
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1676037725
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1676037725
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1676037725
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1676037725
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1676037725
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1676037725
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1676037725
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1676037725
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1676037725
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1676037725
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1676037725
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1676037725
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1676037725
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1676037725
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1676037725
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1676037725
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1676037725
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1676037725
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1676037725
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_9
timestamp 1676037725
transform 1 0 1932 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_21
timestamp 1676037725
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1676037725
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1676037725
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_209
timestamp 1676037725
transform 1 0 20332 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_217
timestamp 1676037725
transform 1 0 21068 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_228
timestamp 1676037725
transform 1 0 22080 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_241
timestamp 1676037725
transform 1 0 23276 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_249
timestamp 1676037725
transform 1 0 24012 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_263
timestamp 1676037725
transform 1 0 25300 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_275
timestamp 1676037725
transform 1 0 26404 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_287
timestamp 1676037725
transform 1 0 27508 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_299
timestamp 1676037725
transform 1 0 28612 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1676037725
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1676037725
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1676037725
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1676037725
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1676037725
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1676037725
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1676037725
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1676037725
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1676037725
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1676037725
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1676037725
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1676037725
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1676037725
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1676037725
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1676037725
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1676037725
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1676037725
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1676037725
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1676037725
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1676037725
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1676037725
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1676037725
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1676037725
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1676037725
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1676037725
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1676037725
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1676037725
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1676037725
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1676037725
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1676037725
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1676037725
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1676037725
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1676037725
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1676037725
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1676037725
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1676037725
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1676037725
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1676037725
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1676037725
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1676037725
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1676037725
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1676037725
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1676037725
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1676037725
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1676037725
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1676037725
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1676037725
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1676037725
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1676037725
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1676037725
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1676037725
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1676037725
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1676037725
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1676037725
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1676037725
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1676037725
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1676037725
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1676037725
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1676037725
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1676037725
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1676037725
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1676037725
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1676037725
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1676037725
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1676037725
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_617
timestamp 1676037725
transform 1 0 57868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_623
timestamp 1676037725
transform 1 0 58420 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_9
timestamp 1676037725
transform 1 0 1932 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_21
timestamp 1676037725
transform 1 0 3036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_229
timestamp 1676037725
transform 1 0 22172 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_239
timestamp 1676037725
transform 1 0 23092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1676037725
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1676037725
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1676037725
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1676037725
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1676037725
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1676037725
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1676037725
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1676037725
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1676037725
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1676037725
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1676037725
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1676037725
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1676037725
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1676037725
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1676037725
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1676037725
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_430
timestamp 1676037725
transform 1 0 40664 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_442
timestamp 1676037725
transform 1 0 41768 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_454
timestamp 1676037725
transform 1 0 42872 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_466
timestamp 1676037725
transform 1 0 43976 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_474
timestamp 1676037725
transform 1 0 44712 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1676037725
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1676037725
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1676037725
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1676037725
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1676037725
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1676037725
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1676037725
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1676037725
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1676037725
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1676037725
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1676037725
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1676037725
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1676037725
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1676037725
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1676037725
transform 1 0 57500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_623
timestamp 1676037725
transform 1 0 58420 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_9
timestamp 1676037725
transform 1 0 1932 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_21
timestamp 1676037725
transform 1 0 3036 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_33
timestamp 1676037725
transform 1 0 4140 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_45
timestamp 1676037725
transform 1 0 5244 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1676037725
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1676037725
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1676037725
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1676037725
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1676037725
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_195
timestamp 1676037725
transform 1 0 19044 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_204
timestamp 1676037725
transform 1 0 19872 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_216
timestamp 1676037725
transform 1 0 20976 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_233
timestamp 1676037725
transform 1 0 22540 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_246
timestamp 1676037725
transform 1 0 23736 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_258
timestamp 1676037725
transform 1 0 24840 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_270
timestamp 1676037725
transform 1 0 25944 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1676037725
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1676037725
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1676037725
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1676037725
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1676037725
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1676037725
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1676037725
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1676037725
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1676037725
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1676037725
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1676037725
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1676037725
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_417
timestamp 1676037725
transform 1 0 39468 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_432
timestamp 1676037725
transform 1 0 40848 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_444
timestamp 1676037725
transform 1 0 41952 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1676037725
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1676037725
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1676037725
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1676037725
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1676037725
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1676037725
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1676037725
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1676037725
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1676037725
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1676037725
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1676037725
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1676037725
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1676037725
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1676037725
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1676037725
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1676037725
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1676037725
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1676037725
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_9
timestamp 1676037725
transform 1 0 1932 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_23
timestamp 1676037725
transform 1 0 3220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_205
timestamp 1676037725
transform 1 0 19964 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_216
timestamp 1676037725
transform 1 0 20976 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_228
timestamp 1676037725
transform 1 0 22080 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_237
timestamp 1676037725
transform 1 0 22908 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1676037725
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_262
timestamp 1676037725
transform 1 0 25208 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_274
timestamp 1676037725
transform 1 0 26312 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_286
timestamp 1676037725
transform 1 0 27416 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_298
timestamp 1676037725
transform 1 0 28520 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1676037725
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1676037725
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1676037725
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1676037725
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1676037725
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1676037725
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1676037725
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1676037725
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1676037725
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1676037725
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1676037725
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1676037725
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1676037725
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1676037725
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1676037725
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1676037725
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1676037725
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1676037725
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1676037725
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1676037725
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1676037725
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1676037725
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1676037725
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1676037725
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1676037725
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1676037725
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1676037725
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1676037725
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1676037725
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 1676037725
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_623
timestamp 1676037725
transform 1 0 58420 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_9
timestamp 1676037725
transform 1 0 1932 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_21
timestamp 1676037725
transform 1 0 3036 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_33
timestamp 1676037725
transform 1 0 4140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_45
timestamp 1676037725
transform 1 0 5244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 1676037725
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_196
timestamp 1676037725
transform 1 0 19136 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_212
timestamp 1676037725
transform 1 0 20608 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_221
timestamp 1676037725
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_237
timestamp 1676037725
transform 1 0 22908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_241
timestamp 1676037725
transform 1 0 23276 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_244
timestamp 1676037725
transform 1 0 23552 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_252
timestamp 1676037725
transform 1 0 24288 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_264
timestamp 1676037725
transform 1 0 25392 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1676037725
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1676037725
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1676037725
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1676037725
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1676037725
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1676037725
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1676037725
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1676037725
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1676037725
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1676037725
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1676037725
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1676037725
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1676037725
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1676037725
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1676037725
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1676037725
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1676037725
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1676037725
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1676037725
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1676037725
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1676037725
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1676037725
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1676037725
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1676037725
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1676037725
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1676037725
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1676037725
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_561
timestamp 1676037725
transform 1 0 52716 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_569
timestamp 1676037725
transform 1 0 53452 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_579
timestamp 1676037725
transform 1 0 54372 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_591
timestamp 1676037725
transform 1 0 55476 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_603
timestamp 1676037725
transform 1 0 56580 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1676037725
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1676037725
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_64
timestamp 1676037725
transform 1 0 6992 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_76
timestamp 1676037725
transform 1 0 8096 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_222
timestamp 1676037725
transform 1 0 21528 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_234
timestamp 1676037725
transform 1 0 22632 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_246
timestamp 1676037725
transform 1 0 23736 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1676037725
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1676037725
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1676037725
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1676037725
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1676037725
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1676037725
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1676037725
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1676037725
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1676037725
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1676037725
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1676037725
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1676037725
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1676037725
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1676037725
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1676037725
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1676037725
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1676037725
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1676037725
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1676037725
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1676037725
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1676037725
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1676037725
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1676037725
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1676037725
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1676037725
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1676037725
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1676037725
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_569
timestamp 1676037725
transform 1 0 53452 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_580
timestamp 1676037725
transform 1 0 54464 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1676037725
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1676037725
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_613
timestamp 1676037725
transform 1 0 57500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_623
timestamp 1676037725
transform 1 0 58420 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_9
timestamp 1676037725
transform 1 0 1932 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_21
timestamp 1676037725
transform 1 0 3036 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_33
timestamp 1676037725
transform 1 0 4140 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_45
timestamp 1676037725
transform 1 0 5244 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_53
timestamp 1676037725
transform 1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1676037725
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_180
timestamp 1676037725
transform 1 0 17664 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_192
timestamp 1676037725
transform 1 0 18768 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_206
timestamp 1676037725
transform 1 0 20056 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_210
timestamp 1676037725
transform 1 0 20424 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_218
timestamp 1676037725
transform 1 0 21160 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_233
timestamp 1676037725
transform 1 0 22540 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_242
timestamp 1676037725
transform 1 0 23368 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_255
timestamp 1676037725
transform 1 0 24564 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_266
timestamp 1676037725
transform 1 0 25576 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_278
timestamp 1676037725
transform 1 0 26680 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1676037725
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1676037725
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1676037725
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1676037725
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1676037725
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1676037725
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1676037725
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1676037725
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1676037725
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1676037725
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1676037725
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1676037725
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1676037725
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1676037725
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1676037725
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1676037725
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1676037725
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1676037725
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1676037725
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1676037725
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1676037725
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1676037725
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1676037725
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1676037725
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1676037725
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1676037725
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1676037725
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1676037725
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1676037725
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1676037725
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1676037725
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1676037725
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_617
timestamp 1676037725
transform 1 0 57868 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_623
timestamp 1676037725
transform 1 0 58420 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_9
timestamp 1676037725
transform 1 0 1932 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_17
timestamp 1676037725
transform 1 0 2668 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_26
timestamp 1676037725
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_201
timestamp 1676037725
transform 1 0 19596 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_204
timestamp 1676037725
transform 1 0 19872 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_212
timestamp 1676037725
transform 1 0 20608 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_224
timestamp 1676037725
transform 1 0 21712 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_236
timestamp 1676037725
transform 1 0 22816 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1676037725
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1676037725
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1676037725
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1676037725
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1676037725
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1676037725
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1676037725
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1676037725
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1676037725
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1676037725
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1676037725
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1676037725
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1676037725
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1676037725
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1676037725
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1676037725
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1676037725
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1676037725
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1676037725
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1676037725
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1676037725
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1676037725
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1676037725
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1676037725
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1676037725
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1676037725
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1676037725
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1676037725
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1676037725
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1676037725
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1676037725
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1676037725
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1676037725
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1676037725
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1676037725
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_613
timestamp 1676037725
transform 1 0 57500 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_623
timestamp 1676037725
transform 1 0 58420 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_9
timestamp 1676037725
transform 1 0 1932 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_21
timestamp 1676037725
transform 1 0 3036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_33
timestamp 1676037725
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1676037725
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1676037725
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_236
timestamp 1676037725
transform 1 0 22816 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_240
timestamp 1676037725
transform 1 0 23184 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_252
timestamp 1676037725
transform 1 0 24288 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_264
timestamp 1676037725
transform 1 0 25392 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1676037725
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1676037725
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1676037725
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1676037725
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1676037725
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1676037725
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1676037725
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1676037725
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1676037725
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1676037725
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1676037725
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1676037725
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1676037725
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1676037725
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1676037725
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1676037725
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1676037725
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1676037725
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1676037725
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1676037725
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1676037725
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1676037725
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1676037725
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1676037725
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1676037725
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1676037725
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1676037725
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1676037725
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1676037725
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1676037725
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1676037725
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1676037725
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1676037725
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1676037725
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_9
timestamp 1676037725
transform 1 0 1932 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_21
timestamp 1676037725
transform 1 0 3036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1676037725
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1676037725
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1676037725
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1676037725
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1676037725
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1676037725
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1676037725
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1676037725
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1676037725
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1676037725
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1676037725
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1676037725
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1676037725
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1676037725
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1676037725
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1676037725
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1676037725
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1676037725
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1676037725
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1676037725
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1676037725
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1676037725
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1676037725
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1676037725
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1676037725
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1676037725
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1676037725
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1676037725
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1676037725
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1676037725
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1676037725
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1676037725
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1676037725
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1676037725
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1676037725
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1676037725
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1676037725
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_601
timestamp 1676037725
transform 1 0 56396 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_613
timestamp 1676037725
transform 1 0 57500 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_623
timestamp 1676037725
transform 1 0 58420 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_9
timestamp 1676037725
transform 1 0 1932 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_21
timestamp 1676037725
transform 1 0 3036 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_33
timestamp 1676037725
transform 1 0 4140 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_45
timestamp 1676037725
transform 1 0 5244 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_53
timestamp 1676037725
transform 1 0 5980 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_213
timestamp 1676037725
transform 1 0 20700 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1676037725
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1676037725
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1676037725
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1676037725
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1676037725
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1676037725
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1676037725
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1676037725
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1676037725
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1676037725
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1676037725
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1676037725
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1676037725
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1676037725
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1676037725
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1676037725
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1676037725
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1676037725
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1676037725
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1676037725
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1676037725
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1676037725
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1676037725
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1676037725
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1676037725
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1676037725
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1676037725
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1676037725
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1676037725
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1676037725
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1676037725
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1676037725
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1676037725
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1676037725
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1676037725
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1676037725
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1676037725
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1676037725
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1676037725
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1676037725
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1676037725
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1676037725
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1676037725
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_9
timestamp 1676037725
transform 1 0 1932 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_21
timestamp 1676037725
transform 1 0 3036 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1676037725
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1676037725
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1676037725
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1676037725
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1676037725
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1676037725
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1676037725
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1676037725
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1676037725
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1676037725
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1676037725
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1676037725
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1676037725
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1676037725
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1676037725
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1676037725
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1676037725
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1676037725
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1676037725
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1676037725
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1676037725
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1676037725
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1676037725
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1676037725
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1676037725
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1676037725
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1676037725
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1676037725
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1676037725
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1676037725
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1676037725
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1676037725
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1676037725
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1676037725
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1676037725
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1676037725
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1676037725
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1676037725
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1676037725
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1676037725
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_601
timestamp 1676037725
transform 1 0 56396 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_613
timestamp 1676037725
transform 1 0 57500 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_623
timestamp 1676037725
transform 1 0 58420 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_9
timestamp 1676037725
transform 1 0 1932 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_21
timestamp 1676037725
transform 1 0 3036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_33
timestamp 1676037725
transform 1 0 4140 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_45
timestamp 1676037725
transform 1 0 5244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1676037725
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1676037725
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1676037725
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1676037725
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1676037725
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1676037725
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1676037725
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1676037725
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1676037725
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1676037725
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1676037725
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1676037725
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1676037725
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1676037725
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1676037725
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1676037725
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1676037725
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1676037725
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1676037725
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1676037725
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1676037725
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1676037725
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1676037725
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1676037725
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1676037725
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1676037725
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1676037725
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1676037725
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1676037725
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1676037725
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1676037725
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1676037725
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1676037725
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1676037725
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1676037725
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1676037725
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1676037725
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1676037725
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1676037725
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1676037725
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1676037725
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1676037725
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1676037725
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1676037725
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1676037725
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_11
timestamp 1676037725
transform 1 0 2116 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_23
timestamp 1676037725
transform 1 0 3220 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1676037725
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1676037725
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1676037725
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1676037725
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1676037725
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1676037725
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1676037725
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1676037725
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1676037725
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1676037725
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1676037725
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1676037725
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1676037725
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1676037725
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1676037725
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1676037725
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1676037725
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1676037725
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1676037725
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1676037725
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1676037725
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1676037725
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1676037725
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1676037725
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1676037725
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1676037725
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1676037725
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1676037725
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1676037725
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1676037725
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1676037725
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1676037725
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1676037725
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1676037725
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1676037725
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1676037725
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1676037725
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1676037725
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1676037725
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1676037725
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1676037725
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_601
timestamp 1676037725
transform 1 0 56396 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_613
timestamp 1676037725
transform 1 0 57500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_623
timestamp 1676037725
transform 1 0 58420 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_9
timestamp 1676037725
transform 1 0 1932 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_21
timestamp 1676037725
transform 1 0 3036 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_33
timestamp 1676037725
transform 1 0 4140 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_45
timestamp 1676037725
transform 1 0 5244 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_53
timestamp 1676037725
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1676037725
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1676037725
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1676037725
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1676037725
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1676037725
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1676037725
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1676037725
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1676037725
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1676037725
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1676037725
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1676037725
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1676037725
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1676037725
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1676037725
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1676037725
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1676037725
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1676037725
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1676037725
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1676037725
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1676037725
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1676037725
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1676037725
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1676037725
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1676037725
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1676037725
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1676037725
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1676037725
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1676037725
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1676037725
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1676037725
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1676037725
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1676037725
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1676037725
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1676037725
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1676037725
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1676037725
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1676037725
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1676037725
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1676037725
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1676037725
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1676037725
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1676037725
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1676037725
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1676037725
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1676037725
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1676037725
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1676037725
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1676037725
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1676037725
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1676037725
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1676037725
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1676037725
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1676037725
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1676037725
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1676037725
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1676037725
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1676037725
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1676037725
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1676037725
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1676037725
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1676037725
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1676037725
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1676037725
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1676037725
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1676037725
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1676037725
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1676037725
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1676037725
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1676037725
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_333
timestamp 1676037725
transform 1 0 31740 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_341
timestamp 1676037725
transform 1 0 32476 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_359
timestamp 1676037725
transform 1 0 34132 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1676037725
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1676037725
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1676037725
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_389
timestamp 1676037725
transform 1 0 36892 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_400
timestamp 1676037725
transform 1 0 37904 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_412
timestamp 1676037725
transform 1 0 39008 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1676037725
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1676037725
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1676037725
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1676037725
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1676037725
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1676037725
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1676037725
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1676037725
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1676037725
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1676037725
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1676037725
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1676037725
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1676037725
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1676037725
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1676037725
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1676037725
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1676037725
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1676037725
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1676037725
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_601
timestamp 1676037725
transform 1 0 56396 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_613
timestamp 1676037725
transform 1 0 57500 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_623
timestamp 1676037725
transform 1 0 58420 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_9
timestamp 1676037725
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_21
timestamp 1676037725
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_33
timestamp 1676037725
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1676037725
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1676037725
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1676037725
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1676037725
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1676037725
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1676037725
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1676037725
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1676037725
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1676037725
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1676037725
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1676037725
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1676037725
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1676037725
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1676037725
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1676037725
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1676037725
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1676037725
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1676037725
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1676037725
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1676037725
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1676037725
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_347
timestamp 1676037725
transform 1 0 33028 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_359
timestamp 1676037725
transform 1 0 34132 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_371
timestamp 1676037725
transform 1 0 35236 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_383
timestamp 1676037725
transform 1 0 36340 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1676037725
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1676037725
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1676037725
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1676037725
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1676037725
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1676037725
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1676037725
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1676037725
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1676037725
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1676037725
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1676037725
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1676037725
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1676037725
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1676037725
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1676037725
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1676037725
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1676037725
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1676037725
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1676037725
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1676037725
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1676037725
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1676037725
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1676037725
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1676037725
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1676037725
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_617
timestamp 1676037725
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_9
timestamp 1676037725
transform 1 0 1932 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_21
timestamp 1676037725
transform 1 0 3036 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1676037725
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1676037725
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1676037725
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1676037725
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1676037725
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1676037725
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1676037725
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1676037725
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1676037725
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1676037725
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1676037725
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1676037725
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1676037725
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1676037725
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1676037725
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1676037725
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_345
timestamp 1676037725
transform 1 0 32844 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_353
timestamp 1676037725
transform 1 0 33580 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_362
timestamp 1676037725
transform 1 0 34408 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1676037725
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1676037725
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1676037725
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1676037725
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1676037725
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1676037725
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1676037725
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1676037725
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1676037725
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1676037725
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1676037725
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1676037725
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1676037725
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1676037725
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1676037725
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1676037725
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1676037725
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1676037725
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1676037725
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1676037725
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1676037725
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1676037725
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1676037725
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1676037725
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1676037725
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1676037725
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_613
timestamp 1676037725
transform 1 0 57500 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_623
timestamp 1676037725
transform 1 0 58420 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_9
timestamp 1676037725
transform 1 0 1932 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_21
timestamp 1676037725
transform 1 0 3036 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_33
timestamp 1676037725
transform 1 0 4140 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_45
timestamp 1676037725
transform 1 0 5244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1676037725
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1676037725
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1676037725
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1676037725
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1676037725
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1676037725
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1676037725
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1676037725
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1676037725
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1676037725
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1676037725
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1676037725
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1676037725
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1676037725
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1676037725
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1676037725
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1676037725
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1676037725
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1676037725
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1676037725
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1676037725
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1676037725
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1676037725
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1676037725
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1676037725
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1676037725
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1676037725
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1676037725
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1676037725
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1676037725
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1676037725
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1676037725
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1676037725
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1676037725
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1676037725
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1676037725
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1676037725
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1676037725
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1676037725
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1676037725
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1676037725
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1676037725
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1676037725
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1676037725
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1676037725
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1676037725
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1676037725
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1676037725
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1676037725
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1676037725
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_617
timestamp 1676037725
transform 1 0 57868 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_11
timestamp 1676037725
transform 1 0 2116 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_23
timestamp 1676037725
transform 1 0 3220 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1676037725
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1676037725
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1676037725
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1676037725
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1676037725
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1676037725
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1676037725
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1676037725
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1676037725
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1676037725
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1676037725
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1676037725
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1676037725
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1676037725
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1676037725
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1676037725
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1676037725
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1676037725
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1676037725
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1676037725
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1676037725
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1676037725
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1676037725
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_365
timestamp 1676037725
transform 1 0 34684 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_375
timestamp 1676037725
transform 1 0 35604 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_387
timestamp 1676037725
transform 1 0 36708 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_399
timestamp 1676037725
transform 1 0 37812 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_411
timestamp 1676037725
transform 1 0 38916 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1676037725
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1676037725
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1676037725
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1676037725
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1676037725
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1676037725
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1676037725
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1676037725
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1676037725
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1676037725
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1676037725
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1676037725
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1676037725
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1676037725
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1676037725
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1676037725
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1676037725
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1676037725
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1676037725
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1676037725
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_601
timestamp 1676037725
transform 1 0 56396 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_613
timestamp 1676037725
transform 1 0 57500 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_623
timestamp 1676037725
transform 1 0 58420 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1676037725
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1676037725
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1676037725
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1676037725
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_173
timestamp 1676037725
transform 1 0 17020 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_183
timestamp 1676037725
transform 1 0 17940 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_195
timestamp 1676037725
transform 1 0 19044 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_207
timestamp 1676037725
transform 1 0 20148 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_219
timestamp 1676037725
transform 1 0 21252 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1676037725
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1676037725
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1676037725
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1676037725
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1676037725
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1676037725
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1676037725
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1676037725
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1676037725
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1676037725
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1676037725
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1676037725
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_373
timestamp 1676037725
transform 1 0 35420 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_381
timestamp 1676037725
transform 1 0 36156 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_390
timestamp 1676037725
transform 1 0 36984 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_393
timestamp 1676037725
transform 1 0 37260 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_409
timestamp 1676037725
transform 1 0 38732 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_421
timestamp 1676037725
transform 1 0 39836 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_433
timestamp 1676037725
transform 1 0 40940 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_445
timestamp 1676037725
transform 1 0 42044 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1676037725
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1676037725
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1676037725
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1676037725
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1676037725
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1676037725
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1676037725
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1676037725
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1676037725
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1676037725
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1676037725
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1676037725
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1676037725
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1676037725
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1676037725
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1676037725
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1676037725
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1676037725
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_617
timestamp 1676037725
transform 1 0 57868 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_623
timestamp 1676037725
transform 1 0 58420 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_9
timestamp 1676037725
transform 1 0 1932 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1676037725
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1676037725
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1676037725
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1676037725
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1676037725
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1676037725
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1676037725
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1676037725
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1676037725
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1676037725
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1676037725
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1676037725
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1676037725
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1676037725
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1676037725
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1676037725
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1676037725
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1676037725
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1676037725
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1676037725
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1676037725
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1676037725
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1676037725
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1676037725
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1676037725
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1676037725
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1676037725
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1676037725
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1676037725
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1676037725
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1676037725
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1676037725
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1676037725
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1676037725
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1676037725
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1676037725
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1676037725
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1676037725
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1676037725
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1676037725
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1676037725
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1676037725
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1676037725
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1676037725
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1676037725
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1676037725
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1676037725
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1676037725
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1676037725
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1676037725
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_613
timestamp 1676037725
transform 1 0 57500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_623
timestamp 1676037725
transform 1 0 58420 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_9
timestamp 1676037725
transform 1 0 1932 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_21
timestamp 1676037725
transform 1 0 3036 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_33
timestamp 1676037725
transform 1 0 4140 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_45
timestamp 1676037725
transform 1 0 5244 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_53
timestamp 1676037725
transform 1 0 5980 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1676037725
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1676037725
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1676037725
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1676037725
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1676037725
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1676037725
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1676037725
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1676037725
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1676037725
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1676037725
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1676037725
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1676037725
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1676037725
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1676037725
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1676037725
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1676037725
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1676037725
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1676037725
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1676037725
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1676037725
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1676037725
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1676037725
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1676037725
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1676037725
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1676037725
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1676037725
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1676037725
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1676037725
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1676037725
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1676037725
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1676037725
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1676037725
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1676037725
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1676037725
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1676037725
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1676037725
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1676037725
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1676037725
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1676037725
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1676037725
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1676037725
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1676037725
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1676037725
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1676037725
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1676037725
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1676037725
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_9
timestamp 1676037725
transform 1 0 1932 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1676037725
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1676037725
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1676037725
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1676037725
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1676037725
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1676037725
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1676037725
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1676037725
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1676037725
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1676037725
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1676037725
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1676037725
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1676037725
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1676037725
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1676037725
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1676037725
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1676037725
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1676037725
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1676037725
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1676037725
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1676037725
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1676037725
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1676037725
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1676037725
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1676037725
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1676037725
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1676037725
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1676037725
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1676037725
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1676037725
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1676037725
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1676037725
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1676037725
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1676037725
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1676037725
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1676037725
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1676037725
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1676037725
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1676037725
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1676037725
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1676037725
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1676037725
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1676037725
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1676037725
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_9
timestamp 1676037725
transform 1 0 1932 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_21
timestamp 1676037725
transform 1 0 3036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_33
timestamp 1676037725
transform 1 0 4140 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_45
timestamp 1676037725
transform 1 0 5244 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_53
timestamp 1676037725
transform 1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1676037725
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1676037725
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1676037725
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1676037725
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1676037725
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1676037725
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1676037725
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1676037725
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1676037725
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1676037725
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1676037725
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1676037725
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1676037725
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1676037725
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1676037725
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1676037725
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1676037725
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1676037725
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1676037725
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1676037725
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1676037725
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1676037725
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1676037725
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1676037725
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1676037725
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1676037725
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1676037725
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1676037725
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1676037725
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1676037725
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1676037725
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1676037725
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1676037725
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1676037725
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1676037725
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1676037725
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1676037725
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1676037725
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1676037725
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1676037725
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1676037725
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1676037725
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1676037725
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1676037725
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_617
timestamp 1676037725
transform 1 0 57868 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_623
timestamp 1676037725
transform 1 0 58420 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_9
timestamp 1676037725
transform 1 0 1932 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_18
timestamp 1676037725
transform 1 0 2760 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_26
timestamp 1676037725
transform 1 0 3496 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1676037725
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1676037725
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1676037725
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1676037725
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1676037725
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1676037725
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1676037725
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1676037725
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1676037725
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1676037725
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1676037725
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1676037725
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1676037725
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1676037725
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1676037725
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1676037725
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1676037725
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1676037725
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1676037725
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1676037725
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1676037725
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1676037725
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1676037725
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1676037725
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1676037725
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1676037725
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1676037725
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1676037725
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1676037725
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1676037725
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1676037725
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1676037725
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1676037725
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1676037725
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1676037725
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1676037725
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1676037725
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1676037725
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1676037725
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_613
timestamp 1676037725
transform 1 0 57500 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_623
timestamp 1676037725
transform 1 0 58420 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_9
timestamp 1676037725
transform 1 0 1932 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_21
timestamp 1676037725
transform 1 0 3036 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_33
timestamp 1676037725
transform 1 0 4140 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_45
timestamp 1676037725
transform 1 0 5244 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_53
timestamp 1676037725
transform 1 0 5980 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1676037725
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1676037725
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1676037725
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1676037725
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1676037725
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1676037725
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1676037725
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1676037725
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1676037725
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1676037725
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1676037725
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1676037725
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1676037725
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1676037725
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1676037725
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1676037725
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1676037725
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1676037725
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1676037725
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1676037725
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1676037725
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1676037725
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1676037725
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1676037725
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1676037725
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1676037725
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1676037725
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1676037725
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1676037725
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1676037725
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1676037725
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1676037725
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1676037725
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1676037725
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1676037725
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1676037725
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1676037725
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1676037725
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1676037725
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_617
timestamp 1676037725
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_9
timestamp 1676037725
transform 1 0 1932 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1676037725
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1676037725
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1676037725
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1676037725
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1676037725
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1676037725
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1676037725
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1676037725
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1676037725
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1676037725
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1676037725
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1676037725
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1676037725
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1676037725
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1676037725
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1676037725
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1676037725
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1676037725
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1676037725
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1676037725
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1676037725
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1676037725
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1676037725
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1676037725
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1676037725
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1676037725
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1676037725
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1676037725
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1676037725
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1676037725
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1676037725
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1676037725
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1676037725
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1676037725
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1676037725
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1676037725
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1676037725
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1676037725
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1676037725
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1676037725
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1676037725
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_613
timestamp 1676037725
transform 1 0 57500 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_623
timestamp 1676037725
transform 1 0 58420 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_9
timestamp 1676037725
transform 1 0 1932 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_21
timestamp 1676037725
transform 1 0 3036 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_33
timestamp 1676037725
transform 1 0 4140 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_45
timestamp 1676037725
transform 1 0 5244 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_53
timestamp 1676037725
transform 1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1676037725
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1676037725
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1676037725
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1676037725
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1676037725
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1676037725
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1676037725
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1676037725
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1676037725
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1676037725
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1676037725
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1676037725
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1676037725
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1676037725
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1676037725
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1676037725
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1676037725
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1676037725
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1676037725
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1676037725
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1676037725
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1676037725
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1676037725
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1676037725
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1676037725
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1676037725
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1676037725
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1676037725
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1676037725
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1676037725
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1676037725
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1676037725
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1676037725
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1676037725
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1676037725
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1676037725
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1676037725
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1676037725
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1676037725
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1676037725
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_9
timestamp 1676037725
transform 1 0 1932 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_21
timestamp 1676037725
transform 1 0 3036 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1676037725
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1676037725
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1676037725
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1676037725
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1676037725
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1676037725
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1676037725
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1676037725
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1676037725
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1676037725
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1676037725
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1676037725
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1676037725
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1676037725
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1676037725
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1676037725
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1676037725
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1676037725
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1676037725
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1676037725
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1676037725
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1676037725
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1676037725
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1676037725
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1676037725
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1676037725
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1676037725
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1676037725
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1676037725
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1676037725
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1676037725
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1676037725
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1676037725
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1676037725
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1676037725
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1676037725
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1676037725
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1676037725
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1676037725
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1676037725
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1676037725
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1676037725
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1676037725
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1676037725
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_613
timestamp 1676037725
transform 1 0 57500 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_623
timestamp 1676037725
transform 1 0 58420 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1676037725
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_27
timestamp 1676037725
transform 1 0 3588 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_36
timestamp 1676037725
transform 1 0 4416 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_48
timestamp 1676037725
transform 1 0 5520 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1676037725
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1676037725
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1676037725
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1676037725
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1676037725
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1676037725
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1676037725
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1676037725
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1676037725
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1676037725
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1676037725
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1676037725
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1676037725
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1676037725
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1676037725
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1676037725
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1676037725
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1676037725
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1676037725
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1676037725
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1676037725
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1676037725
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1676037725
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1676037725
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1676037725
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1676037725
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1676037725
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1676037725
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1676037725
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1676037725
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1676037725
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1676037725
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1676037725
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1676037725
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1676037725
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1676037725
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1676037725
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1676037725
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1676037725
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1676037725
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_9
timestamp 1676037725
transform 1 0 1932 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_21
timestamp 1676037725
transform 1 0 3036 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1676037725
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1676037725
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1676037725
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1676037725
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1676037725
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1676037725
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1676037725
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1676037725
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1676037725
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1676037725
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1676037725
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1676037725
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1676037725
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1676037725
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1676037725
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1676037725
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1676037725
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1676037725
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1676037725
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1676037725
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1676037725
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1676037725
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1676037725
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1676037725
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1676037725
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1676037725
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1676037725
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1676037725
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1676037725
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1676037725
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1676037725
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1676037725
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1676037725
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1676037725
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1676037725
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1676037725
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1676037725
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1676037725
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1676037725
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1676037725
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1676037725
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1676037725
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1676037725
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_613
timestamp 1676037725
transform 1 0 57500 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_619
timestamp 1676037725
transform 1 0 58052 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_623
timestamp 1676037725
transform 1 0 58420 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_9
timestamp 1676037725
transform 1 0 1932 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_21
timestamp 1676037725
transform 1 0 3036 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_33
timestamp 1676037725
transform 1 0 4140 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_45
timestamp 1676037725
transform 1 0 5244 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_53
timestamp 1676037725
transform 1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_69
timestamp 1676037725
transform 1 0 7452 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_79
timestamp 1676037725
transform 1 0 8372 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_91
timestamp 1676037725
transform 1 0 9476 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_103
timestamp 1676037725
transform 1 0 10580 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1676037725
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_91_220
timestamp 1676037725
transform 1 0 21344 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1676037725
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1676037725
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1676037725
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1676037725
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1676037725
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1676037725
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1676037725
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1676037725
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1676037725
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1676037725
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1676037725
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1676037725
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1676037725
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1676037725
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1676037725
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1676037725
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1676037725
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1676037725
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1676037725
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1676037725
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1676037725
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1676037725
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1676037725
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1676037725
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1676037725
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1676037725
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1676037725
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1676037725
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1676037725
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1676037725
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1676037725
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1676037725
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1676037725
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1676037725
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1676037725
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1676037725
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1676037725
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1676037725
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1676037725
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_11
timestamp 1676037725
transform 1 0 2116 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_23
timestamp 1676037725
transform 1 0 3220 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1676037725
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1676037725
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1676037725
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1676037725
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1676037725
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1676037725
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1676037725
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1676037725
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1676037725
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1676037725
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1676037725
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1676037725
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1676037725
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1676037725
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_261
timestamp 1676037725
transform 1 0 25116 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_273
timestamp 1676037725
transform 1 0 26220 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_285
timestamp 1676037725
transform 1 0 27324 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_297
timestamp 1676037725
transform 1 0 28428 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_305
timestamp 1676037725
transform 1 0 29164 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1676037725
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1676037725
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1676037725
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1676037725
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1676037725
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1676037725
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1676037725
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1676037725
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1676037725
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1676037725
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1676037725
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1676037725
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1676037725
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1676037725
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1676037725
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1676037725
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1676037725
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1676037725
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1676037725
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1676037725
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1676037725
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1676037725
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1676037725
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1676037725
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1676037725
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1676037725
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1676037725
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1676037725
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1676037725
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1676037725
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1676037725
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1676037725
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1676037725
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_9
timestamp 1676037725
transform 1 0 1932 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_21
timestamp 1676037725
transform 1 0 3036 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_33
timestamp 1676037725
transform 1 0 4140 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_45
timestamp 1676037725
transform 1 0 5244 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_53
timestamp 1676037725
transform 1 0 5980 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1676037725
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1676037725
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1676037725
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1676037725
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1676037725
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1676037725
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1676037725
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1676037725
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1676037725
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_237
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_243
timestamp 1676037725
transform 1 0 23460 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_251
timestamp 1676037725
transform 1 0 24196 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1676037725
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1676037725
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1676037725
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1676037725
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1676037725
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1676037725
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1676037725
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1676037725
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1676037725
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1676037725
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1676037725
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1676037725
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1676037725
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1676037725
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1676037725
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1676037725
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1676037725
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1676037725
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1676037725
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1676037725
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1676037725
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1676037725
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1676037725
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1676037725
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1676037725
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1676037725
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1676037725
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1676037725
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1676037725
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1676037725
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1676037725
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1676037725
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1676037725
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1676037725
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1676037725
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1676037725
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1676037725
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1676037725
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1676037725
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_93_617
timestamp 1676037725
transform 1 0 57868 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_623
timestamp 1676037725
transform 1 0 58420 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1676037725
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1676037725
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1676037725
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1676037725
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1676037725
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1676037725
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1676037725
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1676037725
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1676037725
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1676037725
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1676037725
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1676037725
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1676037725
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1676037725
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1676037725
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1676037725
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1676037725
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1676037725
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1676037725
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1676037725
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1676037725
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1676037725
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1676037725
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1676037725
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1676037725
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1676037725
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1676037725
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1676037725
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1676037725
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1676037725
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1676037725
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1676037725
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1676037725
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1676037725
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_421
timestamp 1676037725
transform 1 0 39836 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_425
timestamp 1676037725
transform 1 0 40204 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_435
timestamp 1676037725
transform 1 0 41124 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_447
timestamp 1676037725
transform 1 0 42228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_459
timestamp 1676037725
transform 1 0 43332 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_471
timestamp 1676037725
transform 1 0 44436 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1676037725
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1676037725
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1676037725
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1676037725
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1676037725
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1676037725
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1676037725
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1676037725
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1676037725
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1676037725
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1676037725
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1676037725
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1676037725
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1676037725
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1676037725
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1676037725
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_21
timestamp 1676037725
transform 1 0 3036 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_33
timestamp 1676037725
transform 1 0 4140 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_45
timestamp 1676037725
transform 1 0 5244 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_53
timestamp 1676037725
transform 1 0 5980 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1676037725
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1676037725
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1676037725
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1676037725
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1676037725
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1676037725
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1676037725
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1676037725
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1676037725
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1676037725
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1676037725
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1676037725
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1676037725
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1676037725
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1676037725
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1676037725
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1676037725
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1676037725
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1676037725
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1676037725
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1676037725
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1676037725
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1676037725
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1676037725
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1676037725
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1676037725
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1676037725
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1676037725
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1676037725
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1676037725
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1676037725
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1676037725
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1676037725
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1676037725
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1676037725
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1676037725
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1676037725
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1676037725
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1676037725
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1676037725
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1676037725
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1676037725
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1676037725
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1676037725
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1676037725
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1676037725
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1676037725
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1676037725
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1676037725
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1676037725
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1676037725
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1676037725
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1676037725
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1676037725
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1676037725
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_617
timestamp 1676037725
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_96_3
timestamp 1676037725
transform 1 0 1380 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_9
timestamp 1676037725
transform 1 0 1932 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_21
timestamp 1676037725
transform 1 0 3036 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1676037725
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1676037725
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1676037725
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1676037725
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1676037725
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1676037725
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1676037725
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1676037725
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1676037725
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1676037725
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1676037725
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1676037725
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1676037725
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1676037725
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1676037725
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1676037725
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1676037725
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1676037725
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1676037725
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1676037725
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1676037725
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1676037725
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_233
timestamp 1676037725
transform 1 0 22540 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_250
timestamp 1676037725
transform 1 0 24104 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1676037725
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1676037725
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1676037725
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1676037725
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1676037725
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1676037725
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1676037725
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1676037725
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1676037725
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1676037725
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1676037725
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1676037725
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1676037725
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1676037725
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1676037725
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1676037725
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1676037725
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1676037725
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1676037725
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1676037725
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1676037725
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1676037725
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1676037725
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1676037725
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1676037725
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1676037725
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1676037725
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1676037725
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1676037725
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1676037725
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1676037725
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1676037725
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1676037725
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1676037725
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1676037725
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1676037725
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1676037725
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1676037725
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_613
timestamp 1676037725
transform 1 0 57500 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_619
timestamp 1676037725
transform 1 0 58052 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_623
timestamp 1676037725
transform 1 0 58420 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_3
timestamp 1676037725
transform 1 0 1380 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_9
timestamp 1676037725
transform 1 0 1932 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_21
timestamp 1676037725
transform 1 0 3036 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_33
timestamp 1676037725
transform 1 0 4140 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_45
timestamp 1676037725
transform 1 0 5244 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_53
timestamp 1676037725
transform 1 0 5980 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1676037725
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1676037725
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1676037725
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1676037725
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1676037725
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1676037725
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1676037725
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1676037725
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1676037725
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1676037725
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1676037725
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1676037725
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1676037725
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1676037725
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1676037725
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1676037725
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1676037725
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1676037725
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1676037725
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_237
timestamp 1676037725
transform 1 0 22908 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_245
timestamp 1676037725
transform 1 0 23644 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_260
timestamp 1676037725
transform 1 0 25024 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_272
timestamp 1676037725
transform 1 0 26128 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1676037725
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1676037725
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1676037725
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1676037725
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1676037725
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1676037725
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1676037725
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1676037725
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1676037725
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1676037725
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1676037725
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1676037725
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1676037725
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1676037725
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1676037725
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_429
timestamp 1676037725
transform 1 0 40572 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_97_440
timestamp 1676037725
transform 1 0 41584 0 -1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1676037725
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1676037725
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1676037725
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1676037725
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1676037725
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1676037725
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1676037725
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1676037725
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1676037725
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1676037725
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1676037725
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1676037725
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1676037725
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1676037725
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1676037725
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1676037725
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1676037725
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1676037725
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_617
timestamp 1676037725
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_3
timestamp 1676037725
transform 1 0 1380 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_9
timestamp 1676037725
transform 1 0 1932 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_21
timestamp 1676037725
transform 1 0 3036 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1676037725
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1676037725
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1676037725
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1676037725
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1676037725
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1676037725
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1676037725
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1676037725
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1676037725
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1676037725
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1676037725
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1676037725
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1676037725
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1676037725
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1676037725
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1676037725
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1676037725
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1676037725
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1676037725
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1676037725
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1676037725
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1676037725
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1676037725
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1676037725
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1676037725
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_253
timestamp 1676037725
transform 1 0 24380 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_269
timestamp 1676037725
transform 1 0 25852 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_281
timestamp 1676037725
transform 1 0 26956 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_293
timestamp 1676037725
transform 1 0 28060 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_305
timestamp 1676037725
transform 1 0 29164 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_98_309
timestamp 1676037725
transform 1 0 29532 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_325
timestamp 1676037725
transform 1 0 31004 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_337
timestamp 1676037725
transform 1 0 32108 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_349
timestamp 1676037725
transform 1 0 33212 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_361
timestamp 1676037725
transform 1 0 34316 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1676037725
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1676037725
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1676037725
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1676037725
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1676037725
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1676037725
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1676037725
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1676037725
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1676037725
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1676037725
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1676037725
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1676037725
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1676037725
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1676037725
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1676037725
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1676037725
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1676037725
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1676037725
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1676037725
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1676037725
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1676037725
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1676037725
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1676037725
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1676037725
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1676037725
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1676037725
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_613
timestamp 1676037725
transform 1 0 57500 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_619
timestamp 1676037725
transform 1 0 58052 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_623
timestamp 1676037725
transform 1 0 58420 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1676037725
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1676037725
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1676037725
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1676037725
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1676037725
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1676037725
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1676037725
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1676037725
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1676037725
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1676037725
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1676037725
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1676037725
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1676037725
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1676037725
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1676037725
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1676037725
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1676037725
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1676037725
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1676037725
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1676037725
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1676037725
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1676037725
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1676037725
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1676037725
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1676037725
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1676037725
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1676037725
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1676037725
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1676037725
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1676037725
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1676037725
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1676037725
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1676037725
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1676037725
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1676037725
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1676037725
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1676037725
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1676037725
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1676037725
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1676037725
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1676037725
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1676037725
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1676037725
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1676037725
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1676037725
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_429
timestamp 1676037725
transform 1 0 40572 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_446
timestamp 1676037725
transform 1 0 42136 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1676037725
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1676037725
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1676037725
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1676037725
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1676037725
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1676037725
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1676037725
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1676037725
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1676037725
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1676037725
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1676037725
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1676037725
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1676037725
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1676037725
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1676037725
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1676037725
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1676037725
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1676037725
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_617
timestamp 1676037725
transform 1 0 57868 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1676037725
transform 1 0 58420 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_3
timestamp 1676037725
transform 1 0 1380 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_11
timestamp 1676037725
transform 1 0 2116 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_23
timestamp 1676037725
transform 1 0 3220 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1676037725
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1676037725
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1676037725
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1676037725
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1676037725
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1676037725
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1676037725
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1676037725
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1676037725
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1676037725
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1676037725
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1676037725
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1676037725
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1676037725
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1676037725
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1676037725
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1676037725
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1676037725
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1676037725
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1676037725
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1676037725
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1676037725
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1676037725
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1676037725
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1676037725
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1676037725
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1676037725
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1676037725
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1676037725
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1676037725
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1676037725
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1676037725
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1676037725
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_333
timestamp 1676037725
transform 1 0 31740 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_339
timestamp 1676037725
transform 1 0 32292 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_354
timestamp 1676037725
transform 1 0 33672 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_362
timestamp 1676037725
transform 1 0 34408 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1676037725
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1676037725
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1676037725
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1676037725
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1676037725
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1676037725
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1676037725
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1676037725
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1676037725
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1676037725
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1676037725
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1676037725
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1676037725
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1676037725
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1676037725
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1676037725
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1676037725
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1676037725
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1676037725
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1676037725
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1676037725
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1676037725
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1676037725
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1676037725
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1676037725
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1676037725
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_613
timestamp 1676037725
transform 1 0 57500 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_623
timestamp 1676037725
transform 1 0 58420 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_3
timestamp 1676037725
transform 1 0 1380 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_9
timestamp 1676037725
transform 1 0 1932 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_21
timestamp 1676037725
transform 1 0 3036 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_33
timestamp 1676037725
transform 1 0 4140 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_45
timestamp 1676037725
transform 1 0 5244 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1676037725
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1676037725
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1676037725
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_81
timestamp 1676037725
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_93
timestamp 1676037725
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1676037725
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1676037725
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1676037725
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1676037725
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_137
timestamp 1676037725
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_149
timestamp 1676037725
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_161
timestamp 1676037725
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_167
timestamp 1676037725
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1676037725
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1676037725
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_193
timestamp 1676037725
transform 1 0 18860 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_205
timestamp 1676037725
transform 1 0 19964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_217
timestamp 1676037725
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1676037725
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1676037725
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1676037725
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_249
timestamp 1676037725
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_261
timestamp 1676037725
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_273
timestamp 1676037725
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1676037725
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1676037725
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1676037725
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_305
timestamp 1676037725
transform 1 0 29164 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_317
timestamp 1676037725
transform 1 0 30268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_329
timestamp 1676037725
transform 1 0 31372 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_335
timestamp 1676037725
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1676037725
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1676037725
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_361
timestamp 1676037725
transform 1 0 34316 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_373
timestamp 1676037725
transform 1 0 35420 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_385
timestamp 1676037725
transform 1 0 36524 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_391
timestamp 1676037725
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1676037725
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1676037725
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_417
timestamp 1676037725
transform 1 0 39468 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_429
timestamp 1676037725
transform 1 0 40572 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_441
timestamp 1676037725
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1676037725
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1676037725
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1676037725
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_473
timestamp 1676037725
transform 1 0 44620 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_485
timestamp 1676037725
transform 1 0 45724 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1676037725
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1676037725
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1676037725
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1676037725
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_529
timestamp 1676037725
transform 1 0 49772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_541
timestamp 1676037725
transform 1 0 50876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_553
timestamp 1676037725
transform 1 0 51980 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1676037725
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1676037725
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1676037725
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_585
timestamp 1676037725
transform 1 0 54924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_597
timestamp 1676037725
transform 1 0 56028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_609
timestamp 1676037725
transform 1 0 57132 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1676037725
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_617
timestamp 1676037725
transform 1 0 57868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_102_3
timestamp 1676037725
transform 1 0 1380 0 1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_11
timestamp 1676037725
transform 1 0 2116 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_23
timestamp 1676037725
transform 1 0 3220 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1676037725
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1676037725
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1676037725
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1676037725
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_65
timestamp 1676037725
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1676037725
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1676037725
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_85
timestamp 1676037725
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_97
timestamp 1676037725
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_109
timestamp 1676037725
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_121
timestamp 1676037725
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1676037725
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1676037725
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_141
timestamp 1676037725
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_153
timestamp 1676037725
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_165
timestamp 1676037725
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_177
timestamp 1676037725
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_189
timestamp 1676037725
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_195
timestamp 1676037725
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_197
timestamp 1676037725
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_209
timestamp 1676037725
transform 1 0 20332 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_221
timestamp 1676037725
transform 1 0 21436 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_233
timestamp 1676037725
transform 1 0 22540 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_245
timestamp 1676037725
transform 1 0 23644 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_251
timestamp 1676037725
transform 1 0 24196 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_253
timestamp 1676037725
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_265
timestamp 1676037725
transform 1 0 25484 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_277
timestamp 1676037725
transform 1 0 26588 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_289
timestamp 1676037725
transform 1 0 27692 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_301
timestamp 1676037725
transform 1 0 28796 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_307
timestamp 1676037725
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_309
timestamp 1676037725
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_321
timestamp 1676037725
transform 1 0 30636 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_333
timestamp 1676037725
transform 1 0 31740 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_345
timestamp 1676037725
transform 1 0 32844 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_357
timestamp 1676037725
transform 1 0 33948 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_363
timestamp 1676037725
transform 1 0 34500 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_365
timestamp 1676037725
transform 1 0 34684 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_369
timestamp 1676037725
transform 1 0 35052 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_387
timestamp 1676037725
transform 1 0 36708 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_399
timestamp 1676037725
transform 1 0 37812 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_411
timestamp 1676037725
transform 1 0 38916 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_102_419
timestamp 1676037725
transform 1 0 39652 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_421
timestamp 1676037725
transform 1 0 39836 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_433
timestamp 1676037725
transform 1 0 40940 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_445
timestamp 1676037725
transform 1 0 42044 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_457
timestamp 1676037725
transform 1 0 43148 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_469
timestamp 1676037725
transform 1 0 44252 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_475
timestamp 1676037725
transform 1 0 44804 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_477
timestamp 1676037725
transform 1 0 44988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_489
timestamp 1676037725
transform 1 0 46092 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_501
timestamp 1676037725
transform 1 0 47196 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_513
timestamp 1676037725
transform 1 0 48300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_525
timestamp 1676037725
transform 1 0 49404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_531
timestamp 1676037725
transform 1 0 49956 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_533
timestamp 1676037725
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_545
timestamp 1676037725
transform 1 0 51244 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_557
timestamp 1676037725
transform 1 0 52348 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_569
timestamp 1676037725
transform 1 0 53452 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_581
timestamp 1676037725
transform 1 0 54556 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_587
timestamp 1676037725
transform 1 0 55108 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_589
timestamp 1676037725
transform 1 0 55292 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_601
timestamp 1676037725
transform 1 0 56396 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_613
timestamp 1676037725
transform 1 0 57500 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_102_623
timestamp 1676037725
transform 1 0 58420 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_3
timestamp 1676037725
transform 1 0 1380 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_11
timestamp 1676037725
transform 1 0 2116 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_23
timestamp 1676037725
transform 1 0 3220 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_35
timestamp 1676037725
transform 1 0 4324 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_47
timestamp 1676037725
transform 1 0 5428 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1676037725
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1676037725
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_69
timestamp 1676037725
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_81
timestamp 1676037725
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_93
timestamp 1676037725
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1676037725
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1676037725
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_113
timestamp 1676037725
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_125
timestamp 1676037725
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_137
timestamp 1676037725
transform 1 0 13708 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_149
timestamp 1676037725
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_161
timestamp 1676037725
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_167
timestamp 1676037725
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_169
timestamp 1676037725
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_181
timestamp 1676037725
transform 1 0 17756 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_193
timestamp 1676037725
transform 1 0 18860 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_205
timestamp 1676037725
transform 1 0 19964 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_217
timestamp 1676037725
transform 1 0 21068 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_223
timestamp 1676037725
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_225
timestamp 1676037725
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_237
timestamp 1676037725
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_249
timestamp 1676037725
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_261
timestamp 1676037725
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_273
timestamp 1676037725
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_279
timestamp 1676037725
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_281
timestamp 1676037725
transform 1 0 26956 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_293
timestamp 1676037725
transform 1 0 28060 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_305
timestamp 1676037725
transform 1 0 29164 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_317
timestamp 1676037725
transform 1 0 30268 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_329
timestamp 1676037725
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_335
timestamp 1676037725
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_337
timestamp 1676037725
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_349
timestamp 1676037725
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_361
timestamp 1676037725
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_103_373
timestamp 1676037725
transform 1 0 35420 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_103_384
timestamp 1676037725
transform 1 0 36432 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_103_393
timestamp 1676037725
transform 1 0 37260 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_412
timestamp 1676037725
transform 1 0 39008 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_424
timestamp 1676037725
transform 1 0 40112 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_103_446
timestamp 1676037725
transform 1 0 42136 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_449
timestamp 1676037725
transform 1 0 42412 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_461
timestamp 1676037725
transform 1 0 43516 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_473
timestamp 1676037725
transform 1 0 44620 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_485
timestamp 1676037725
transform 1 0 45724 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_497
timestamp 1676037725
transform 1 0 46828 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_503
timestamp 1676037725
transform 1 0 47380 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_505
timestamp 1676037725
transform 1 0 47564 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_517
timestamp 1676037725
transform 1 0 48668 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_529
timestamp 1676037725
transform 1 0 49772 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_541
timestamp 1676037725
transform 1 0 50876 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_553
timestamp 1676037725
transform 1 0 51980 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_559
timestamp 1676037725
transform 1 0 52532 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_561
timestamp 1676037725
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_573
timestamp 1676037725
transform 1 0 53820 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_585
timestamp 1676037725
transform 1 0 54924 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_597
timestamp 1676037725
transform 1 0 56028 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_609
timestamp 1676037725
transform 1 0 57132 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_615
timestamp 1676037725
transform 1 0 57684 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_103_617
timestamp 1676037725
transform 1 0 57868 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_623
timestamp 1676037725
transform 1 0 58420 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_104_3
timestamp 1676037725
transform 1 0 1380 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_9
timestamp 1676037725
transform 1 0 1932 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_21
timestamp 1676037725
transform 1 0 3036 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1676037725
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1676037725
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1676037725
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1676037725
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_65
timestamp 1676037725
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1676037725
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1676037725
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_85
timestamp 1676037725
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_97
timestamp 1676037725
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_109
timestamp 1676037725
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_121
timestamp 1676037725
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_133
timestamp 1676037725
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_139
timestamp 1676037725
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_141
timestamp 1676037725
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_153
timestamp 1676037725
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_165
timestamp 1676037725
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_177
timestamp 1676037725
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_189
timestamp 1676037725
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_195
timestamp 1676037725
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_104_197
timestamp 1676037725
transform 1 0 19228 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_207
timestamp 1676037725
transform 1 0 20148 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_219
timestamp 1676037725
transform 1 0 21252 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_231
timestamp 1676037725
transform 1 0 22356 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_243
timestamp 1676037725
transform 1 0 23460 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_251
timestamp 1676037725
transform 1 0 24196 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_253
timestamp 1676037725
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_265
timestamp 1676037725
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_277
timestamp 1676037725
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_289
timestamp 1676037725
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_301
timestamp 1676037725
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_307
timestamp 1676037725
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_309
timestamp 1676037725
transform 1 0 29532 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_321
timestamp 1676037725
transform 1 0 30636 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_333
timestamp 1676037725
transform 1 0 31740 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_345
timestamp 1676037725
transform 1 0 32844 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_357
timestamp 1676037725
transform 1 0 33948 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_363
timestamp 1676037725
transform 1 0 34500 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_365
timestamp 1676037725
transform 1 0 34684 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_377
timestamp 1676037725
transform 1 0 35788 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_389
timestamp 1676037725
transform 1 0 36892 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_401
timestamp 1676037725
transform 1 0 37996 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_413
timestamp 1676037725
transform 1 0 39100 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_419
timestamp 1676037725
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_421
timestamp 1676037725
transform 1 0 39836 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_104_429
timestamp 1676037725
transform 1 0 40572 0 1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_104_446
timestamp 1676037725
transform 1 0 42136 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_458
timestamp 1676037725
transform 1 0 43240 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_470
timestamp 1676037725
transform 1 0 44344 0 1 58752
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_104_477
timestamp 1676037725
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_489
timestamp 1676037725
transform 1 0 46092 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_501
timestamp 1676037725
transform 1 0 47196 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_513
timestamp 1676037725
transform 1 0 48300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_525
timestamp 1676037725
transform 1 0 49404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_531
timestamp 1676037725
transform 1 0 49956 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_533
timestamp 1676037725
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_545
timestamp 1676037725
transform 1 0 51244 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_557
timestamp 1676037725
transform 1 0 52348 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_569
timestamp 1676037725
transform 1 0 53452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_581
timestamp 1676037725
transform 1 0 54556 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_587
timestamp 1676037725
transform 1 0 55108 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_589
timestamp 1676037725
transform 1 0 55292 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_601
timestamp 1676037725
transform 1 0 56396 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_104_613
timestamp 1676037725
transform 1 0 57500 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_104_623
timestamp 1676037725
transform 1 0 58420 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_3
timestamp 1676037725
transform 1 0 1380 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_105_11
timestamp 1676037725
transform 1 0 2116 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_105_19
timestamp 1676037725
transform 1 0 2852 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_31
timestamp 1676037725
transform 1 0 3956 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_43
timestamp 1676037725
transform 1 0 5060 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1676037725
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_57
timestamp 1676037725
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_69
timestamp 1676037725
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_81
timestamp 1676037725
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_93
timestamp 1676037725
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1676037725
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1676037725
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_113
timestamp 1676037725
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_125
timestamp 1676037725
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_137
timestamp 1676037725
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_149
timestamp 1676037725
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_161
timestamp 1676037725
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_167
timestamp 1676037725
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_169
timestamp 1676037725
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_181
timestamp 1676037725
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_193
timestamp 1676037725
transform 1 0 18860 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_205
timestamp 1676037725
transform 1 0 19964 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_213
timestamp 1676037725
transform 1 0 20700 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_222
timestamp 1676037725
transform 1 0 21528 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_105_225
timestamp 1676037725
transform 1 0 21804 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_236
timestamp 1676037725
transform 1 0 22816 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_105_248
timestamp 1676037725
transform 1 0 23920 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_260
timestamp 1676037725
transform 1 0 25024 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_272
timestamp 1676037725
transform 1 0 26128 0 -1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_105_281
timestamp 1676037725
transform 1 0 26956 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_105_293
timestamp 1676037725
transform 1 0 28060 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_302
timestamp 1676037725
transform 1 0 28888 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_306
timestamp 1676037725
transform 1 0 29256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_309
timestamp 1676037725
transform 1 0 29532 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_319
timestamp 1676037725
transform 1 0 30452 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_323
timestamp 1676037725
transform 1 0 30820 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_335
timestamp 1676037725
transform 1 0 31924 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_337
timestamp 1676037725
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_349
timestamp 1676037725
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_361
timestamp 1676037725
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_373
timestamp 1676037725
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_385
timestamp 1676037725
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_391
timestamp 1676037725
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_393
timestamp 1676037725
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_405
timestamp 1676037725
transform 1 0 38364 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_417
timestamp 1676037725
transform 1 0 39468 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_429
timestamp 1676037725
transform 1 0 40572 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_441
timestamp 1676037725
transform 1 0 41676 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_447
timestamp 1676037725
transform 1 0 42228 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_449
timestamp 1676037725
transform 1 0 42412 0 -1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_105_465
timestamp 1676037725
transform 1 0 43884 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_477
timestamp 1676037725
transform 1 0 44988 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_489
timestamp 1676037725
transform 1 0 46092 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_105_501
timestamp 1676037725
transform 1 0 47196 0 -1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_105_505
timestamp 1676037725
transform 1 0 47564 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_517
timestamp 1676037725
transform 1 0 48668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_529
timestamp 1676037725
transform 1 0 49772 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_541
timestamp 1676037725
transform 1 0 50876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_553
timestamp 1676037725
transform 1 0 51980 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_559
timestamp 1676037725
transform 1 0 52532 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_561
timestamp 1676037725
transform 1 0 52716 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_573
timestamp 1676037725
transform 1 0 53820 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_585
timestamp 1676037725
transform 1 0 54924 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_597
timestamp 1676037725
transform 1 0 56028 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_609
timestamp 1676037725
transform 1 0 57132 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_614
timestamp 1676037725
transform 1 0 57592 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_617
timestamp 1676037725
transform 1 0 57868 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_623
timestamp 1676037725
transform 1 0 58420 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_3
timestamp 1676037725
transform 1 0 1380 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_106_11
timestamp 1676037725
transform 1 0 2116 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_106_19
timestamp 1676037725
transform 1 0 2852 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1676037725
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1676037725
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1676037725
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_53
timestamp 1676037725
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_65
timestamp 1676037725
transform 1 0 7084 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_106_75
timestamp 1676037725
transform 1 0 8004 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1676037725
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_85
timestamp 1676037725
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_97
timestamp 1676037725
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_109
timestamp 1676037725
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_121
timestamp 1676037725
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_133
timestamp 1676037725
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_139
timestamp 1676037725
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_141
timestamp 1676037725
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_153
timestamp 1676037725
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_165
timestamp 1676037725
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_191
timestamp 1676037725
transform 1 0 18676 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_195
timestamp 1676037725
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_106_197
timestamp 1676037725
transform 1 0 19228 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_106_207
timestamp 1676037725
transform 1 0 20148 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_211
timestamp 1676037725
transform 1 0 20516 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_220
timestamp 1676037725
transform 1 0 21344 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_241
timestamp 1676037725
transform 1 0 23276 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_249
timestamp 1676037725
transform 1 0 24012 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_253
timestamp 1676037725
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_265
timestamp 1676037725
transform 1 0 25484 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_277
timestamp 1676037725
transform 1 0 26588 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_291
timestamp 1676037725
transform 1 0 27876 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_302
timestamp 1676037725
transform 1 0 28888 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_306
timestamp 1676037725
transform 1 0 29256 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_106_309
timestamp 1676037725
transform 1 0 29532 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_313
timestamp 1676037725
transform 1 0 29900 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_106_316
timestamp 1676037725
transform 1 0 30176 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_106_327
timestamp 1676037725
transform 1 0 31188 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_333
timestamp 1676037725
transform 1 0 31740 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_349
timestamp 1676037725
transform 1 0 33212 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_361
timestamp 1676037725
transform 1 0 34316 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_365
timestamp 1676037725
transform 1 0 34684 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_377
timestamp 1676037725
transform 1 0 35788 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_389
timestamp 1676037725
transform 1 0 36892 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_401
timestamp 1676037725
transform 1 0 37996 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_413
timestamp 1676037725
transform 1 0 39100 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_419
timestamp 1676037725
transform 1 0 39652 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_421
timestamp 1676037725
transform 1 0 39836 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_429
timestamp 1676037725
transform 1 0 40572 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_438
timestamp 1676037725
transform 1 0 41400 0 1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_106_456
timestamp 1676037725
transform 1 0 43056 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_468
timestamp 1676037725
transform 1 0 44160 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_106_477
timestamp 1676037725
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_489
timestamp 1676037725
transform 1 0 46092 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_501
timestamp 1676037725
transform 1 0 47196 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_513
timestamp 1676037725
transform 1 0 48300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_525
timestamp 1676037725
transform 1 0 49404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_531
timestamp 1676037725
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_533
timestamp 1676037725
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_545
timestamp 1676037725
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_557
timestamp 1676037725
transform 1 0 52348 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_569
timestamp 1676037725
transform 1 0 53452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_581
timestamp 1676037725
transform 1 0 54556 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_587
timestamp 1676037725
transform 1 0 55108 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_589
timestamp 1676037725
transform 1 0 55292 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_605
timestamp 1676037725
transform 1 0 56764 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_613
timestamp 1676037725
transform 1 0 57500 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_623
timestamp 1676037725
transform 1 0 58420 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_3
timestamp 1676037725
transform 1 0 1380 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_107_11
timestamp 1676037725
transform 1 0 2116 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_19
timestamp 1676037725
transform 1 0 2852 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_26
timestamp 1676037725
transform 1 0 3496 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_34
timestamp 1676037725
transform 1 0 4232 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_46
timestamp 1676037725
transform 1 0 5336 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_54
timestamp 1676037725
transform 1 0 6072 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1676037725
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_69
timestamp 1676037725
transform 1 0 7452 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_77
timestamp 1676037725
transform 1 0 8188 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_82
timestamp 1676037725
transform 1 0 8648 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_90
timestamp 1676037725
transform 1 0 9384 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_102
timestamp 1676037725
transform 1 0 10488 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_110
timestamp 1676037725
transform 1 0 11224 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_113
timestamp 1676037725
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_125
timestamp 1676037725
transform 1 0 12604 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_133
timestamp 1676037725
transform 1 0 13340 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_138
timestamp 1676037725
transform 1 0 13800 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_146
timestamp 1676037725
transform 1 0 14536 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_162
timestamp 1676037725
transform 1 0 16008 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_169
timestamp 1676037725
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_181
timestamp 1676037725
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_193
timestamp 1676037725
transform 1 0 18860 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_197
timestamp 1676037725
transform 1 0 19228 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_202
timestamp 1676037725
transform 1 0 19688 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_214
timestamp 1676037725
transform 1 0 20792 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_222
timestamp 1676037725
transform 1 0 21528 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_225
timestamp 1676037725
transform 1 0 21804 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_107_233
timestamp 1676037725
transform 1 0 22540 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_239
timestamp 1676037725
transform 1 0 23092 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_247
timestamp 1676037725
transform 1 0 23828 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_253
timestamp 1676037725
transform 1 0 24380 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_258
timestamp 1676037725
transform 1 0 24840 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_270
timestamp 1676037725
transform 1 0 25944 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_278
timestamp 1676037725
transform 1 0 26680 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_107_281
timestamp 1676037725
transform 1 0 26956 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_285
timestamp 1676037725
transform 1 0 27324 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_290
timestamp 1676037725
transform 1 0 27784 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_306
timestamp 1676037725
transform 1 0 29256 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_316
timestamp 1676037725
transform 1 0 30176 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_322
timestamp 1676037725
transform 1 0 30728 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_334
timestamp 1676037725
transform 1 0 31832 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_337
timestamp 1676037725
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_349
timestamp 1676037725
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_361
timestamp 1676037725
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_373
timestamp 1676037725
transform 1 0 35420 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_381
timestamp 1676037725
transform 1 0 36156 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_386
timestamp 1676037725
transform 1 0 36616 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_393
timestamp 1676037725
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_405
timestamp 1676037725
transform 1 0 38364 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_417
timestamp 1676037725
transform 1 0 39468 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_429
timestamp 1676037725
transform 1 0 40572 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_437
timestamp 1676037725
transform 1 0 41308 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_442
timestamp 1676037725
transform 1 0 41768 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_449
timestamp 1676037725
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_461
timestamp 1676037725
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_473
timestamp 1676037725
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_485
timestamp 1676037725
transform 1 0 45724 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_493
timestamp 1676037725
transform 1 0 46460 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_498
timestamp 1676037725
transform 1 0 46920 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_505
timestamp 1676037725
transform 1 0 47564 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_517
timestamp 1676037725
transform 1 0 48668 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_529
timestamp 1676037725
transform 1 0 49772 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_533
timestamp 1676037725
transform 1 0 50140 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_538
timestamp 1676037725
transform 1 0 50600 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_550
timestamp 1676037725
transform 1 0 51704 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_558
timestamp 1676037725
transform 1 0 52440 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_561
timestamp 1676037725
transform 1 0 52716 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_567
timestamp 1676037725
transform 1 0 53268 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_107_579
timestamp 1676037725
transform 1 0 54372 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_586
timestamp 1676037725
transform 1 0 55016 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_594
timestamp 1676037725
transform 1 0 55752 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_602
timestamp 1676037725
transform 1 0 56488 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_107_610
timestamp 1676037725
transform 1 0 57224 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_107_617
timestamp 1676037725
transform 1 0 57868 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_623
timestamp 1676037725
transform 1 0 58420 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_3
timestamp 1676037725
transform 1 0 1380 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_14
timestamp 1676037725
transform 1 0 2392 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_24
timestamp 1676037725
transform 1 0 3312 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_29
timestamp 1676037725
transform 1 0 3772 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_33
timestamp 1676037725
transform 1 0 4140 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_38
timestamp 1676037725
transform 1 0 4600 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_46
timestamp 1676037725
transform 1 0 5336 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_54
timestamp 1676037725
transform 1 0 6072 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_108_57
timestamp 1676037725
transform 1 0 6348 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_66
timestamp 1676037725
transform 1 0 7176 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_76
timestamp 1676037725
transform 1 0 8096 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_108_85
timestamp 1676037725
transform 1 0 8924 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_89
timestamp 1676037725
transform 1 0 9292 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_94
timestamp 1676037725
transform 1 0 9752 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_102
timestamp 1676037725
transform 1 0 10488 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_110
timestamp 1676037725
transform 1 0 11224 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_113
timestamp 1676037725
transform 1 0 11500 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_117
timestamp 1676037725
transform 1 0 11868 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_122
timestamp 1676037725
transform 1 0 12328 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_132
timestamp 1676037725
transform 1 0 13248 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_108_141
timestamp 1676037725
transform 1 0 14076 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_149
timestamp 1676037725
transform 1 0 14812 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_156
timestamp 1676037725
transform 1 0 15456 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_108_166
timestamp 1676037725
transform 1 0 16376 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_169
timestamp 1676037725
transform 1 0 16652 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_173
timestamp 1676037725
transform 1 0 17020 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_178
timestamp 1676037725
transform 1 0 17480 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_186
timestamp 1676037725
transform 1 0 18216 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_194
timestamp 1676037725
transform 1 0 18952 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_197
timestamp 1676037725
transform 1 0 19228 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_201
timestamp 1676037725
transform 1 0 19596 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_206
timestamp 1676037725
transform 1 0 20056 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_214
timestamp 1676037725
transform 1 0 20792 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_222
timestamp 1676037725
transform 1 0 21528 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_225
timestamp 1676037725
transform 1 0 21804 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_229
timestamp 1676037725
transform 1 0 22172 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_236
timestamp 1676037725
transform 1 0 22816 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_244
timestamp 1676037725
transform 1 0 23552 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_250
timestamp 1676037725
transform 1 0 24104 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_253
timestamp 1676037725
transform 1 0 24380 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_261
timestamp 1676037725
transform 1 0 25116 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_268
timestamp 1676037725
transform 1 0 25760 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_276
timestamp 1676037725
transform 1 0 26496 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_281
timestamp 1676037725
transform 1 0 26956 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_289
timestamp 1676037725
transform 1 0 27692 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_293
timestamp 1676037725
transform 1 0 28060 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_300
timestamp 1676037725
transform 1 0 28704 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_309
timestamp 1676037725
transform 1 0 29532 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_317
timestamp 1676037725
transform 1 0 30268 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_325
timestamp 1676037725
transform 1 0 31004 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_332
timestamp 1676037725
transform 1 0 31648 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_337
timestamp 1676037725
transform 1 0 32108 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_345
timestamp 1676037725
transform 1 0 32844 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_353
timestamp 1676037725
transform 1 0 33580 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_108_361
timestamp 1676037725
transform 1 0 34316 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_108_365
timestamp 1676037725
transform 1 0 34684 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_371
timestamp 1676037725
transform 1 0 35236 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_379
timestamp 1676037725
transform 1 0 35972 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_387
timestamp 1676037725
transform 1 0 36708 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_391
timestamp 1676037725
transform 1 0 37076 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_393
timestamp 1676037725
transform 1 0 37260 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_399
timestamp 1676037725
transform 1 0 37812 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_407
timestamp 1676037725
transform 1 0 38548 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_415
timestamp 1676037725
transform 1 0 39284 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_419
timestamp 1676037725
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_421
timestamp 1676037725
transform 1 0 39836 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_427
timestamp 1676037725
transform 1 0 40388 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_435
timestamp 1676037725
transform 1 0 41124 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_443
timestamp 1676037725
transform 1 0 41860 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_447
timestamp 1676037725
transform 1 0 42228 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_449
timestamp 1676037725
transform 1 0 42412 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_457
timestamp 1676037725
transform 1 0 43148 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_465
timestamp 1676037725
transform 1 0 43884 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_108_473
timestamp 1676037725
transform 1 0 44620 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_108_477
timestamp 1676037725
transform 1 0 44988 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_483
timestamp 1676037725
transform 1 0 45540 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_491
timestamp 1676037725
transform 1 0 46276 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_499
timestamp 1676037725
transform 1 0 47012 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_503
timestamp 1676037725
transform 1 0 47380 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_505
timestamp 1676037725
transform 1 0 47564 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_511
timestamp 1676037725
transform 1 0 48116 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_519
timestamp 1676037725
transform 1 0 48852 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_527
timestamp 1676037725
transform 1 0 49588 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_531
timestamp 1676037725
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_533
timestamp 1676037725
transform 1 0 50140 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_541
timestamp 1676037725
transform 1 0 50876 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_549
timestamp 1676037725
transform 1 0 51612 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_108_557
timestamp 1676037725
transform 1 0 52348 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_561
timestamp 1676037725
transform 1 0 52716 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_565
timestamp 1676037725
transform 1 0 53084 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_572
timestamp 1676037725
transform 1 0 53728 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_580
timestamp 1676037725
transform 1 0 54464 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_589
timestamp 1676037725
transform 1 0 55292 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_597
timestamp 1676037725
transform 1 0 56028 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_607
timestamp 1676037725
transform 1 0 56948 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_615
timestamp 1676037725
transform 1 0 57684 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_617
timestamp 1676037725
transform 1 0 57868 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_623
timestamp 1676037725
transform 1 0 58420 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1676037725
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1676037725
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1676037725
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1676037725
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1676037725
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1676037725
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1676037725
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1676037725
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1676037725
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1676037725
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1676037725
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1676037725
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1676037725
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1676037725
transform -1 0 58880 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1676037725
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1676037725
transform -1 0 58880 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1676037725
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1676037725
transform -1 0 58880 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1676037725
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1676037725
transform -1 0 58880 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1676037725
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1676037725
transform -1 0 58880 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1676037725
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1676037725
transform -1 0 58880 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1676037725
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1676037725
transform -1 0 58880 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1676037725
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1676037725
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1676037725
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1676037725
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1676037725
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1676037725
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1676037725
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1676037725
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1676037725
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1676037725
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1676037725
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1676037725
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1676037725
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1676037725
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1676037725
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1676037725
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1676037725
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1676037725
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1676037725
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1676037725
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1676037725
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1676037725
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1676037725
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1676037725
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1676037725
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1676037725
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1676037725
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1676037725
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1676037725
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1676037725
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1676037725
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1676037725
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1676037725
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1676037725
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1676037725
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1676037725
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1676037725
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1676037725
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1676037725
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1676037725
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1676037725
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1676037725
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1676037725
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1676037725
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1676037725
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1676037725
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1676037725
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1676037725
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1676037725
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1676037725
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1676037725
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1676037725
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1676037725
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1676037725
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1676037725
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1676037725
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1676037725
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1676037725
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1676037725
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1676037725
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1676037725
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1676037725
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1676037725
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1676037725
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1676037725
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1676037725
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1676037725
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1676037725
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1676037725
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1676037725
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1676037725
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1676037725
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1676037725
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1676037725
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1676037725
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1676037725
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1676037725
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1676037725
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1676037725
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1676037725
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1676037725
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1676037725
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1676037725
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1676037725
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1676037725
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1676037725
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1676037725
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1676037725
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1676037725
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1676037725
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1676037725
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1676037725
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1676037725
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1676037725
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1676037725
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1676037725
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1676037725
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1676037725
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1676037725
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1676037725
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1676037725
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1676037725
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1676037725
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1676037725
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1676037725
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1676037725
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1676037725
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1676037725
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1676037725
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1676037725
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1676037725
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1676037725
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1676037725
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1676037725
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1676037725
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1676037725
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1676037725
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1676037725
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1676037725
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1676037725
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1676037725
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1676037725
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1676037725
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1676037725
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1676037725
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1676037725
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1676037725
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1676037725
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1676037725
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1676037725
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1676037725
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1676037725
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1676037725
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1676037725
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1676037725
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1676037725
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1676037725
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1676037725
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1676037725
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1676037725
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1676037725
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1676037725
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1676037725
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1676037725
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1676037725
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1676037725
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1676037725
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1676037725
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1676037725
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1676037725
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1676037725
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1676037725
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1676037725
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1676037725
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1676037725
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1676037725
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1676037725
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1676037725
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1676037725
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1676037725
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1676037725
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1676037725
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1676037725
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1676037725
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1676037725
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1676037725
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1676037725
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1676037725
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1676037725
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1676037725
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1676037725
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1676037725
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1676037725
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1676037725
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1676037725
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1676037725
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1676037725
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1676037725
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1676037725
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1676037725
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1676037725
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1676037725
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1676037725
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1676037725
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1676037725
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1676037725
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1676037725
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1676037725
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1676037725
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1676037725
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1676037725
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1676037725
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1676037725
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1676037725
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1676037725
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1676037725
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1676037725
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1676037725
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1676037725
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1676037725
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1676037725
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1676037725
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1676037725
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1676037725
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1676037725
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1676037725
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1676037725
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1676037725
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1676037725
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1676037725
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1676037725
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1676037725
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1676037725
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1676037725
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1676037725
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1676037725
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1676037725
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1676037725
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1676037725
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1676037725
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1676037725
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1676037725
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1676037725
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1676037725
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1676037725
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1676037725
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1676037725
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1676037725
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1676037725
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1676037725
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1676037725
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1676037725
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1676037725
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1676037725
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1676037725
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1676037725
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1676037725
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1676037725
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1676037725
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1676037725
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1676037725
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1676037725
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1676037725
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1676037725
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1676037725
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1676037725
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1676037725
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1676037725
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1676037725
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1676037725
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1676037725
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1676037725
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1676037725
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1676037725
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1676037725
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1676037725
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1676037725
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1676037725
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1676037725
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1676037725
transform 1 0 6256 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1676037725
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1676037725
transform 1 0 11408 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1676037725
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1676037725
transform 1 0 16560 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1676037725
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1676037725
transform 1 0 21712 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1676037725
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1676037725
transform 1 0 26864 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1676037725
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1676037725
transform 1 0 32016 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1676037725
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1676037725
transform 1 0 37168 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1676037725
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1676037725
transform 1 0 42320 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1676037725
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1676037725
transform 1 0 47472 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1676037725
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1676037725
transform 1 0 52624 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1676037725
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1676037725
transform 1 0 57776 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0449_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 40480 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1676037725
transform 1 0 23828 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0451_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0452_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0453_
timestamp 1676037725
transform 1 0 44436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1676037725
transform 1 0 41860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0455_
timestamp 1676037725
transform 1 0 42596 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0456_
timestamp 1676037725
transform 1 0 14904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457_
timestamp 1676037725
transform 1 0 13984 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0458_
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor4b_4  _0459_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15732 0 1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_4  _0460_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2b_1  _0461_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2668 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0462_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor4b_4  _0463_
timestamp 1676037725
transform 1 0 18124 0 -1 8704
box -38 -48 1786 592
use sky130_fd_sc_hd__or3_4  _0464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 12880 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_4  _0465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14996 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0466_
timestamp 1676037725
transform 1 0 9384 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0467_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26496 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor4b_4  _0468_
timestamp 1676037725
transform 1 0 16468 0 1 7616
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_1  _0469_
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0470_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0471_
timestamp 1676037725
transform 1 0 10672 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0472_
timestamp 1676037725
transform 1 0 16836 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0473_
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_2  _0474_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15272 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _0475_
timestamp 1676037725
transform 1 0 11960 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15456 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_4  _0477_
timestamp 1676037725
transform 1 0 16744 0 1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_1  _0478_
timestamp 1676037725
transform 1 0 10672 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0479_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25576 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_4  _0480_
timestamp 1676037725
transform 1 0 15180 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0481_
timestamp 1676037725
transform 1 0 10856 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _0482_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or3_4  _0483_
timestamp 1676037725
transform 1 0 12788 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_4  _0484_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17848 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_2  _0485_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0486_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2b_1  _0487_
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_4  _0488_
timestamp 1676037725
transform 1 0 15916 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_1  _0489_
timestamp 1676037725
transform 1 0 9384 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_4  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25852 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 1 56576
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 37260 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0493_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32568 0 1 42432
box -38 -48 1602 592
use sky130_fd_sc_hd__a221o_1  _0494_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33120 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0495_
timestamp 1676037725
transform 1 0 32936 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29348 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28520 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0498_
timestamp 1676037725
transform 1 0 27324 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0499_
timestamp 1676037725
transform 1 0 29716 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28428 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _0501_
timestamp 1676037725
transform 1 0 27600 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _0502_
timestamp 1676037725
transform 1 0 32292 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0503_
timestamp 1676037725
transform 1 0 43884 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0504_
timestamp 1676037725
transform 1 0 31924 0 1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0505_
timestamp 1676037725
transform 1 0 31556 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0506_
timestamp 1676037725
transform 1 0 35236 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0507_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32752 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _0508_
timestamp 1676037725
transform 1 0 32568 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0509_
timestamp 1676037725
transform 1 0 37996 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0510_
timestamp 1676037725
transform 1 0 38272 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_4  _0511_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0512_
timestamp 1676037725
transform 1 0 53084 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0513_
timestamp 1676037725
transform 1 0 33672 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0514_
timestamp 1676037725
transform 1 0 34224 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0515_
timestamp 1676037725
transform 1 0 35236 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0516_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35052 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0517_
timestamp 1676037725
transform 1 0 37168 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0518_
timestamp 1676037725
transform 1 0 17388 0 1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0519_
timestamp 1676037725
transform 1 0 35880 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0520_
timestamp 1676037725
transform 1 0 37444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0521_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35696 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0522_
timestamp 1676037725
transform 1 0 37444 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0523_
timestamp 1676037725
transform 1 0 37996 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0524_
timestamp 1676037725
transform 1 0 34868 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0525_
timestamp 1676037725
transform 1 0 17112 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0526_
timestamp 1676037725
transform 1 0 18768 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _0527_
timestamp 1676037725
transform 1 0 35144 0 1 57664
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_4  _0528_
timestamp 1676037725
transform 1 0 19412 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_2  _0529_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14720 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0530_
timestamp 1676037725
transform 1 0 31372 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0531_
timestamp 1676037725
transform 1 0 27968 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_2  _0532_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9752 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0533_
timestamp 1676037725
transform 1 0 36340 0 -1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0534_
timestamp 1676037725
transform 1 0 37444 0 -1 58752
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0535_
timestamp 1676037725
transform 1 0 23184 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0536_
timestamp 1676037725
transform 1 0 24564 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0537_
timestamp 1676037725
transform 1 0 24196 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0538_
timestamp 1676037725
transform 1 0 24840 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0539_
timestamp 1676037725
transform 1 0 23000 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0540_
timestamp 1676037725
transform 1 0 21988 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0541_
timestamp 1676037725
transform 1 0 20884 0 -1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0542_
timestamp 1676037725
transform 1 0 21712 0 1 59840
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0543_
timestamp 1676037725
transform 1 0 22816 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0544_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23092 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0545_
timestamp 1676037725
transform 1 0 22540 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0546_
timestamp 1676037725
transform 1 0 19412 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0547_
timestamp 1676037725
transform 1 0 19320 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0548_
timestamp 1676037725
transform 1 0 53636 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0549_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20608 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0550_
timestamp 1676037725
transform 1 0 19228 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0551_
timestamp 1676037725
transform 1 0 18492 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0552_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20976 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0553_
timestamp 1676037725
transform 1 0 20148 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0554_
timestamp 1676037725
transform 1 0 20884 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0555_
timestamp 1676037725
transform 1 0 21988 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0556_
timestamp 1676037725
transform 1 0 53728 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0557_
timestamp 1676037725
transform 1 0 2024 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0558_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3036 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__nor4_4  _0559_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15548 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0560_
timestamp 1676037725
transform 1 0 19412 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0561_
timestamp 1676037725
transform 1 0 20056 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _0562_
timestamp 1676037725
transform 1 0 21712 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_4  _0563_
timestamp 1676037725
transform 1 0 14720 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0564_
timestamp 1676037725
transform 1 0 20608 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0565_
timestamp 1676037725
transform 1 0 22264 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0566_
timestamp 1676037725
transform 1 0 21252 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0567_
timestamp 1676037725
transform 1 0 40020 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0568_
timestamp 1676037725
transform 1 0 2300 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _0569_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22448 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0570_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22448 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1676037725
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _0572_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _0573_
timestamp 1676037725
transform 1 0 22080 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0574_
timestamp 1676037725
transform 1 0 22908 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0575_
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0576_
timestamp 1676037725
transform 1 0 23276 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0577_
timestamp 1676037725
transform 1 0 40204 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0578_
timestamp 1676037725
transform 1 0 23736 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0579_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0580_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25944 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0581_
timestamp 1676037725
transform 1 0 20884 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0582_
timestamp 1676037725
transform 1 0 40112 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _0583_
timestamp 1676037725
transform 1 0 2024 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0584_
timestamp 1676037725
transform 1 0 40664 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _0585_
timestamp 1676037725
transform 1 0 20516 0 -1 52224
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0586_
timestamp 1676037725
transform 1 0 21988 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0587_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0588_
timestamp 1676037725
transform 1 0 30636 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0589_
timestamp 1676037725
transform 1 0 32108 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0590_
timestamp 1676037725
transform 1 0 3680 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _0591_
timestamp 1676037725
transform 1 0 5428 0 1 36992
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0592_
timestamp 1676037725
transform 1 0 27048 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0593_
timestamp 1676037725
transform 1 0 28152 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0594_
timestamp 1676037725
transform 1 0 29716 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0595_
timestamp 1676037725
transform 1 0 31280 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1676037725
transform 1 0 32016 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0597_
timestamp 1676037725
transform 1 0 23092 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0598_
timestamp 1676037725
transform 1 0 23920 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0599_
timestamp 1676037725
transform 1 0 7360 0 1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0600_
timestamp 1676037725
transform 1 0 7728 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0601_
timestamp 1676037725
transform 1 0 22724 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _0602_
timestamp 1676037725
transform 1 0 27140 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_4  _0603_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25760 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0604_
timestamp 1676037725
transform 1 0 23184 0 -1 60928
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0605_
timestamp 1676037725
transform 1 0 23736 0 -1 55488
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0606_
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _0607_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0608_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1676037725
transform 1 0 24748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0610_
timestamp 1676037725
transform 1 0 23552 0 -1 53312
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0611_
timestamp 1676037725
transform 1 0 24932 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0612_
timestamp 1676037725
transform 1 0 22724 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0613_
timestamp 1676037725
transform 1 0 23736 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0614_
timestamp 1676037725
transform 1 0 40388 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0615_
timestamp 1676037725
transform 1 0 42596 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0616_
timestamp 1676037725
transform 1 0 40480 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0617_
timestamp 1676037725
transform 1 0 38456 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0618_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _0619_
timestamp 1676037725
transform 1 0 42596 0 -1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0620_
timestamp 1676037725
transform 1 0 28060 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0621_
timestamp 1676037725
transform 1 0 22816 0 1 54400
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0622_
timestamp 1676037725
transform 1 0 41216 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0623_
timestamp 1676037725
transform 1 0 40848 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0624_
timestamp 1676037725
transform 1 0 41492 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0625_
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0626_
timestamp 1676037725
transform 1 0 42596 0 -1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0627_
timestamp 1676037725
transform -1 0 31188 0 1 59840
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0628_
timestamp 1676037725
transform 1 0 24564 0 1 55488
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0629_
timestamp 1676037725
transform 1 0 40848 0 -1 56576
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0630_
timestamp 1676037725
transform 1 0 41032 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0631_
timestamp 1676037725
transform 1 0 40848 0 -1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0632_
timestamp 1676037725
transform 1 0 42780 0 1 2176
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0633_
timestamp 1676037725
transform 1 0 29716 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0634_
timestamp 1676037725
transform 1 0 29716 0 1 55488
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_4  _0635_
timestamp 1676037725
transform 1 0 32292 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  _0636_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31188 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0637_
timestamp 1676037725
transform 1 0 42596 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0638_
timestamp 1676037725
transform 1 0 42504 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_2  _0639_
timestamp 1676037725
transform 1 0 29164 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0640_
timestamp 1676037725
transform 1 0 41768 0 1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0641_
timestamp 1676037725
transform 1 0 42688 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_2  _0642_
timestamp 1676037725
transform 1 0 32292 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0643_
timestamp 1676037725
transform 1 0 40848 0 1 58752
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0644_
timestamp 1676037725
transform 1 0 40020 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0645_
timestamp 1676037725
transform 1 0 42504 0 1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0646_
timestamp 1676037725
transform 1 0 40848 0 -1 58752
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0647_
timestamp 1676037725
transform 1 0 41124 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0648_
timestamp 1676037725
transform 1 0 40848 0 1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0649_
timestamp 1676037725
transform 1 0 42596 0 -1 59840
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_4  _0650_
timestamp 1676037725
transform 1 0 42872 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__a211o_4  _0651_
timestamp 1676037725
transform 1 0 30544 0 -1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0652_
timestamp 1676037725
transform 1 0 15640 0 1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_2  _0653_
timestamp 1676037725
transform 1 0 13064 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18676 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0655_
timestamp 1676037725
transform 1 0 17572 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0656_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10304 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0657_
timestamp 1676037725
transform 1 0 26772 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0658_
timestamp 1676037725
transform 1 0 8004 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9292 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0660_
timestamp 1676037725
transform 1 0 8372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0661_
timestamp 1676037725
transform 1 0 9384 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0662_
timestamp 1676037725
transform 1 0 7176 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0663_
timestamp 1676037725
transform 1 0 8924 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0664_
timestamp 1676037725
transform 1 0 8096 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0665_
timestamp 1676037725
transform 1 0 9660 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0666_
timestamp 1676037725
transform 1 0 10396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0667_
timestamp 1676037725
transform 1 0 10212 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0668_
timestamp 1676037725
transform 1 0 8924 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0669_
timestamp 1676037725
transform 1 0 9108 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0670_
timestamp 1676037725
transform 1 0 9936 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0671_
timestamp 1676037725
transform 1 0 9108 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0672_
timestamp 1676037725
transform 1 0 10672 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0673_
timestamp 1676037725
transform 1 0 10764 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0674_
timestamp 1676037725
transform 1 0 10396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0675_
timestamp 1676037725
transform 1 0 10580 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0676_
timestamp 1676037725
transform 1 0 12420 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0677_
timestamp 1676037725
transform 1 0 25852 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0678_
timestamp 1676037725
transform 1 0 12788 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0679_
timestamp 1676037725
transform 1 0 29716 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0680_
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0681_
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0682_
timestamp 1676037725
transform 1 0 12604 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0683_
timestamp 1676037725
transform 1 0 24288 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0684_
timestamp 1676037725
transform 1 0 11040 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0685_
timestamp 1676037725
transform 1 0 10948 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0686_
timestamp 1676037725
transform 1 0 11684 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0687_
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0688_
timestamp 1676037725
transform 1 0 12420 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0689_
timestamp 1676037725
transform 1 0 31004 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0690_
timestamp 1676037725
transform 1 0 13156 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0691_
timestamp 1676037725
transform 1 0 23460 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0692_
timestamp 1676037725
transform 1 0 14260 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0693_
timestamp 1676037725
transform 1 0 31096 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0694_
timestamp 1676037725
transform 1 0 13340 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0695_
timestamp 1676037725
transform 1 0 23276 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0696_
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0697_
timestamp 1676037725
transform 1 0 31188 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0698_
timestamp 1676037725
transform 1 0 13340 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0699_
timestamp 1676037725
transform 1 0 13064 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0700_
timestamp 1676037725
transform 1 0 14260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0701_
timestamp 1676037725
transform 1 0 28428 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0702_
timestamp 1676037725
transform 1 0 13064 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0703_
timestamp 1676037725
transform 1 0 13156 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0704_
timestamp 1676037725
transform 1 0 15456 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0705_
timestamp 1676037725
transform 1 0 29440 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _0706_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15732 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_4  _0707_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29716 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_1  _0708_
timestamp 1676037725
transform 1 0 13248 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0709_
timestamp 1676037725
transform 1 0 13524 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0710_
timestamp 1676037725
transform 1 0 8740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0711_
timestamp 1676037725
transform 1 0 9292 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0712_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 57040 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _0713_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43792 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0714_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36156 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1676037725
transform 1 0 36524 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0716_
timestamp 1676037725
transform 1 0 46184 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0717_
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0718_
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0719_
timestamp 1676037725
transform 1 0 34868 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0720_
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1676037725
transform 1 0 35972 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0722_
timestamp 1676037725
transform 1 0 34960 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0723_
timestamp 1676037725
transform 1 0 38732 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0724_
timestamp 1676037725
transform 1 0 38732 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0725_
timestamp 1676037725
transform 1 0 30820 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0726_
timestamp 1676037725
transform 1 0 30912 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0727_
timestamp 1676037725
transform 1 0 25300 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0728_
timestamp 1676037725
transform 1 0 25668 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0729_
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0730_
timestamp 1676037725
transform 1 0 45172 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0731_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43700 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0732_
timestamp 1676037725
transform 1 0 28428 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0733_
timestamp 1676037725
transform 1 0 27692 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0734_
timestamp 1676037725
transform 1 0 32292 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0735_
timestamp 1676037725
transform 1 0 31372 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0736_
timestamp 1676037725
transform 1 0 32292 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0737_
timestamp 1676037725
transform 1 0 33488 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0738_
timestamp 1676037725
transform 1 0 37444 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0739_
timestamp 1676037725
transform 1 0 37628 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 1676037725
transform 1 0 27784 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0741_
timestamp 1676037725
transform 1 0 27600 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1676037725
transform 1 0 29348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0743_
timestamp 1676037725
transform 1 0 28796 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1676037725
transform 1 0 25300 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0745_
timestamp 1676037725
transform 1 0 26496 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0746_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0747_
timestamp 1676037725
transform 1 0 20148 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0749_
timestamp 1676037725
transform 1 0 20976 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0750_
timestamp 1676037725
transform 1 0 20700 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0751_
timestamp 1676037725
transform 1 0 20792 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1676037725
transform 1 0 27968 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0753_
timestamp 1676037725
transform 1 0 27508 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 1676037725
transform 1 0 41676 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0755_
timestamp 1676037725
transform 1 0 41400 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1676037725
transform 1 0 38364 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0757_
timestamp 1676037725
transform 1 0 38364 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 1676037725
transform 1 0 27416 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0759_
timestamp 1676037725
transform 1 0 26404 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1676037725
transform 1 0 27600 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0761_
timestamp 1676037725
transform 1 0 26772 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0762_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0763_
timestamp 1676037725
transform 1 0 20976 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0764_
timestamp 1676037725
transform 1 0 35880 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0765_
timestamp 1676037725
transform 1 0 37444 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0767_
timestamp 1676037725
transform 1 0 25760 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1676037725
transform 1 0 35696 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0769_
timestamp 1676037725
transform 1 0 34408 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0770_
timestamp 1676037725
transform 1 0 25576 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0771_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0772_
timestamp 1676037725
transform 1 0 38732 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0773_
timestamp 1676037725
transform 1 0 38732 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0774_
timestamp 1676037725
transform 1 0 30636 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0775_
timestamp 1676037725
transform 1 0 30544 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 1676037725
transform 1 0 30912 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0777_
timestamp 1676037725
transform 1 0 30084 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 1676037725
transform 1 0 33580 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0779_
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0780_
timestamp 1676037725
transform 1 0 50876 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0781_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1676037725
transform 1 0 27968 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp 1676037725
transform 1 0 23276 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp 1676037725
transform 1 0 18124 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1676037725
transform 1 0 19964 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 1676037725
transform 1 0 20608 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 1676037725
transform 1 0 21988 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1676037725
transform 1 0 20700 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1676037725
transform 1 0 20240 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0790_
timestamp 1676037725
transform 1 0 21620 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1676037725
transform 1 0 41308 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0794_
timestamp 1676037725
transform 1 0 35236 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1676037725
transform 1 0 27232 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0796_
timestamp 1676037725
transform 1 0 25760 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1676037725
transform 1 0 20976 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0798_
timestamp 1676037725
transform 1 0 34500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0799_
timestamp 1676037725
transform 1 0 36248 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp 1676037725
transform 1 0 34868 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1676037725
transform 1 0 33396 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0802_
timestamp 1676037725
transform 1 0 38272 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0803_
timestamp 1676037725
transform 1 0 29072 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0804_
timestamp 1676037725
transform 1 0 40572 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1676037725
transform 1 0 33948 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0806_
timestamp 1676037725
transform 1 0 45816 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp 1676037725
transform 1 0 47748 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1676037725
transform 1 0 46368 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1676037725
transform 1 0 46276 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0810_
timestamp 1676037725
transform 1 0 19412 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0811_
timestamp 1676037725
transform 1 0 19596 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0812_
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 1676037725
transform 1 0 23276 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1676037725
transform 1 0 25760 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp 1676037725
transform 1 0 24748 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1676037725
transform 1 0 23000 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0817_
timestamp 1676037725
transform 1 0 22632 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0818_
timestamp 1676037725
transform 1 0 44252 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0819_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0820_
timestamp 1676037725
transform 1 0 58052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0821_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27508 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0822_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _0823_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 33028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0824_
timestamp 1676037725
transform 1 0 32568 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0825_
timestamp 1676037725
transform 1 0 55752 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1676037725
transform 1 0 55476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0827_
timestamp 1676037725
transform 1 0 30636 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0828_
timestamp 1676037725
transform 1 0 32752 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0829_
timestamp 1676037725
transform 1 0 35972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _0830_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0831_
timestamp 1676037725
transform 1 0 56120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0832_
timestamp 1676037725
transform 1 0 57040 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0833_
timestamp 1676037725
transform 1 0 33856 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0834_
timestamp 1676037725
transform 1 0 34132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _0835_
timestamp 1676037725
transform 1 0 35328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0836_
timestamp 1676037725
transform 1 0 56120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0837_
timestamp 1676037725
transform 1 0 37444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0838_
timestamp 1676037725
transform 1 0 52900 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0839_
timestamp 1676037725
transform 1 0 38272 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0840_
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0841_
timestamp 1676037725
transform 1 0 39836 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0842_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0843_
timestamp 1676037725
transform 1 0 57132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0844_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1676037725
transform 1 0 31280 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _0846_
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0847_
timestamp 1676037725
transform 1 0 31832 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0848_
timestamp 1676037725
transform 1 0 56120 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0849_
timestamp 1676037725
transform 1 0 24288 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0850_
timestamp 1676037725
transform 1 0 23368 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0851_
timestamp 1676037725
transform 1 0 31004 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0853_
timestamp 1676037725
transform 1 0 45632 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43884 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0855_
timestamp 1676037725
transform 1 0 24104 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0856_
timestamp 1676037725
transform 1 0 51060 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0857_
timestamp 1676037725
transform 1 0 51428 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0858_
timestamp 1676037725
transform 1 0 22724 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0859_
timestamp 1676037725
transform 1 0 53636 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0860_
timestamp 1676037725
transform 1 0 53912 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1676037725
transform 1 0 23828 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0862_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23092 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0863_
timestamp 1676037725
transform 1 0 22632 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0864_
timestamp 1676037725
transform 1 0 37812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0865_
timestamp 1676037725
transform 1 0 37352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22816 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0867_
timestamp 1676037725
transform 1 0 38456 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0868_
timestamp 1676037725
transform 1 0 38916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0869_
timestamp 1676037725
transform 1 0 27600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0870_
timestamp 1676037725
transform 1 0 27876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0871_
timestamp 1676037725
transform 1 0 54924 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0872_
timestamp 1676037725
transform 1 0 55936 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0873_
timestamp 1676037725
transform 1 0 30820 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1676037725
transform 1 0 43608 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0875_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 43700 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0876_
timestamp 1676037725
transform 1 0 42596 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0877_
timestamp 1676037725
transform 1 0 29992 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 1676037725
transform 1 0 40480 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0879_
timestamp 1676037725
transform 1 0 42596 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0880_
timestamp 1676037725
transform 1 0 41676 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0881_
timestamp 1676037725
transform 1 0 27232 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0882_
timestamp 1676037725
transform 1 0 28336 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0883_
timestamp 1676037725
transform 1 0 54280 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0884_
timestamp 1676037725
transform 1 0 54556 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0885_
timestamp 1676037725
transform 1 0 25576 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0886_
timestamp 1676037725
transform 1 0 24840 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0887_
timestamp 1676037725
transform 1 0 50600 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0888_
timestamp 1676037725
transform 1 0 51428 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0889_
timestamp 1676037725
transform 1 0 23092 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_2  _0890_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0891_
timestamp 1676037725
transform 1 0 54556 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0892_
timestamp 1676037725
transform 1 0 55476 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0893_
timestamp 1676037725
transform 1 0 37720 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0894_
timestamp 1676037725
transform 1 0 47472 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0895_
timestamp 1676037725
transform 1 0 48116 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _0896_
timestamp 1676037725
transform 1 0 23000 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0897_
timestamp 1676037725
transform 1 0 55476 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0898_
timestamp 1676037725
transform 1 0 55844 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 1676037725
transform 1 0 36708 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0900_
timestamp 1676037725
transform 1 0 49772 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0901_
timestamp 1676037725
transform 1 0 50232 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0902_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0903_
timestamp 1676037725
transform 1 0 52808 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0904_
timestamp 1676037725
transform 1 0 53820 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0905_
timestamp 1676037725
transform 1 0 40572 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0906_
timestamp 1676037725
transform 1 0 45908 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0907_
timestamp 1676037725
transform 1 0 45264 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0908_
timestamp 1676037725
transform 1 0 31648 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0909_
timestamp 1676037725
transform 1 0 32292 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0910_
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0911_
timestamp 1676037725
transform 1 0 45356 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0912_
timestamp 1676037725
transform 1 0 30268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0913_
timestamp 1676037725
transform 1 0 51060 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0914_
timestamp 1676037725
transform 1 0 51428 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0915_
timestamp 1676037725
transform 1 0 32476 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0916_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0917_
timestamp 1676037725
transform 1 0 47932 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0918_
timestamp 1676037725
transform 1 0 48484 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _0919_
timestamp 1676037725
transform 1 0 38180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0920_
timestamp 1676037725
transform 1 0 42136 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0921_
timestamp 1676037725
transform 1 0 43148 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0922_
timestamp 1676037725
transform 1 0 41492 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0923_
timestamp 1676037725
transform 1 0 42780 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a32oi_4  _0924_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32384 0 1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0926_
timestamp 1676037725
transform 1 0 35880 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0927_
timestamp 1676037725
transform 1 0 36248 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0928_
timestamp 1676037725
transform 1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13156 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0930_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _0931_
timestamp 1676037725
transform 1 0 14536 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0932_
timestamp 1676037725
transform 1 0 14996 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0933_
timestamp 1676037725
transform 1 0 16008 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 1676037725
transform 1 0 10488 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0935_
timestamp 1676037725
transform 1 0 10488 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0936_
timestamp 1676037725
transform 1 0 9936 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0937_
timestamp 1676037725
transform 1 0 9384 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _0938_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11868 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0939_
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0940_
timestamp 1676037725
transform 1 0 10672 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0941_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0942_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0943_
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0944_
timestamp 1676037725
transform 1 0 18032 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0945_
timestamp 1676037725
transform 1 0 17296 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0946_
timestamp 1676037725
transform 1 0 17020 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1676037725
transform 1 0 22632 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0948_
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0949_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0950_
timestamp 1676037725
transform 1 0 18308 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and4_2  _0951_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1676037725
transform 1 0 20148 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1676037725
transform 1 0 19872 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0954_
timestamp 1676037725
transform 1 0 18032 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0955_
timestamp 1676037725
transform 1 0 17204 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0956_
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0957_
timestamp 1676037725
transform 1 0 16836 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0958_
timestamp 1676037725
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0959_
timestamp 1676037725
transform 1 0 18952 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1676037725
transform 1 0 19780 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0961_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0962_
timestamp 1676037725
transform 1 0 19320 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0963_
timestamp 1676037725
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0964_
timestamp 1676037725
transform 1 0 19596 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0965_
timestamp 1676037725
transform 1 0 19780 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0966_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _0967_
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0968_
timestamp 1676037725
transform 1 0 16192 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0969_
timestamp 1676037725
transform 1 0 15272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0970_
timestamp 1676037725
transform 1 0 11408 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0971_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0972_
timestamp 1676037725
transform 1 0 11316 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0973_
timestamp 1676037725
transform 1 0 12696 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0974_
timestamp 1676037725
transform 1 0 12788 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0975_
timestamp 1676037725
transform 1 0 10672 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0976_
timestamp 1676037725
transform 1 0 9844 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0977_
timestamp 1676037725
transform 1 0 8004 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0978_
timestamp 1676037725
transform 1 0 10120 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0979_
timestamp 1676037725
transform 1 0 9108 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0980_
timestamp 1676037725
transform 1 0 8004 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0981_
timestamp 1676037725
transform 1 0 7728 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0982_
timestamp 1676037725
transform 1 0 6532 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_2  _0983_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 36064 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0984_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0985_
timestamp 1676037725
transform 1 0 34132 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0986_
timestamp 1676037725
transform 1 0 35696 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0987_
timestamp 1676037725
transform 1 0 38456 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1676037725
transform 1 0 31280 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1676037725
transform 1 0 27140 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1676037725
transform 1 0 19688 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1676037725
transform 1 0 48484 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _0992_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28520 0 -1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0993_
timestamp 1676037725
transform 1 0 32200 0 1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0994_
timestamp 1676037725
transform 1 0 33304 0 -1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0995_
timestamp 1676037725
transform 1 0 36984 0 1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0996_
timestamp 1676037725
transform 1 0 28428 0 -1 3264
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _0997_
timestamp 1676037725
transform 1 0 29716 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0998_
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1676037725
transform 1 0 20792 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1000_
timestamp 1676037725
transform 1 0 20976 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1676037725
transform 1 0 20792 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1676037725
transform 1 0 27508 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1003_
timestamp 1676037725
transform 1 0 41308 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1004_
timestamp 1676037725
transform 1 0 38456 0 -1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1005_
timestamp 1676037725
transform 1 0 27140 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1006_
timestamp 1676037725
transform 1 0 27416 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1676037725
transform 1 0 20700 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1008_
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1009_
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1010_
timestamp 1676037725
transform 1 0 35236 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1676037725
transform 1 0 23736 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1012_
timestamp 1676037725
transform 1 0 38824 0 -1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1013_
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1014_
timestamp 1676037725
transform 1 0 30268 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1015_
timestamp 1676037725
transform 1 0 32844 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1676037725
transform 1 0 56856 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1676037725
transform 1 0 27232 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1676037725
transform 1 0 22632 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1676037725
transform 1 0 19688 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1676037725
transform 1 0 19688 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1676037725
transform 1 0 19780 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1676037725
transform 1 0 19780 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1676037725
transform 1 0 20056 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1676037725
transform 1 0 19504 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1676037725
transform 1 0 19780 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1676037725
transform 1 0 25944 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1676037725
transform 1 0 40664 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1676037725
transform 1 0 34592 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1676037725
transform 1 0 26496 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1676037725
transform 1 0 33764 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1676037725
transform 1 0 36524 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1676037725
transform 1 0 34408 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1676037725
transform 1 0 32936 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1676037725
transform 1 0 37444 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1676037725
transform 1 0 28428 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1676037725
transform 1 0 40204 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1676037725
transform 1 0 33580 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1676037725
transform 1 0 45172 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1042_
timestamp 1676037725
transform 1 0 47748 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1043_
timestamp 1676037725
transform 1 0 45172 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1044_
timestamp 1676037725
transform 1 0 45540 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1676037725
transform 1 0 19412 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1676037725
transform 1 0 23368 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1676037725
transform 1 0 24748 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1676037725
transform 1 0 22448 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1676037725
transform 1 0 56856 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1676037725
transform 1 0 56856 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1051_
timestamp 1676037725
transform 1 0 56856 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1052_
timestamp 1676037725
transform 1 0 40020 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1676037725
transform 1 0 56856 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1676037725
transform 1 0 45172 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1676037725
transform 1 0 51520 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1676037725
transform 1 0 53544 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1057_
timestamp 1676037725
transform 1 0 37996 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1058_
timestamp 1676037725
transform 1 0 40020 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1676037725
transform 1 0 56856 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1676037725
transform 1 0 43240 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1676037725
transform 1 0 42872 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1676037725
transform 1 0 54924 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1676037725
transform 1 0 51612 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1676037725
transform 1 0 55844 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1065_
timestamp 1676037725
transform 1 0 48208 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1676037725
transform 1 0 56856 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1067_
timestamp 1676037725
transform 1 0 50416 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1676037725
transform 1 0 53084 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1069_
timestamp 1676037725
transform 1 0 45448 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1070_
timestamp 1676037725
transform 1 0 46184 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1071_
timestamp 1676037725
transform 1 0 52348 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1072_
timestamp 1676037725
transform 1 0 48668 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1073_
timestamp 1676037725
transform 1 0 42964 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1074_
timestamp 1676037725
transform 1 0 43056 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1075_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1076_
timestamp 1676037725
transform 1 0 36248 0 1 11968
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1077_
timestamp 1676037725
transform 1 0 13432 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1078_
timestamp 1676037725
transform 1 0 14352 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1079_
timestamp 1676037725
transform 1 0 14168 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1080_
timestamp 1676037725
transform 1 0 9384 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1081_
timestamp 1676037725
transform 1 0 9292 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1082_
timestamp 1676037725
transform 1 0 11408 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1083_
timestamp 1676037725
transform 1 0 11040 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1085_
timestamp 1676037725
transform 1 0 16744 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1676037725
transform 1 0 17020 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1676037725
transform 1 0 16836 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1088_
timestamp 1676037725
transform 1 0 14996 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1089_
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1090_
timestamp 1676037725
transform 1 0 16928 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1091_
timestamp 1676037725
transform 1 0 17112 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1093_
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1094_
timestamp 1676037725
transform 1 0 12420 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1095_
timestamp 1676037725
transform 1 0 12052 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1676037725
transform 1 0 12328 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1097_
timestamp 1676037725
transform 1 0 8188 0 -1 18496
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1098_
timestamp 1676037725
transform 1 0 8740 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1099_
timestamp 1676037725
transform 1 0 6808 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1100_
timestamp 1676037725
transform 1 0 6072 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  _1121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 29900 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1676037725
transform 1 0 29900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1123_
timestamp 1676037725
transform 1 0 30636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1676037725
transform 1 0 31464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1125_
timestamp 1676037725
transform 1 0 32752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1126_
timestamp 1676037725
transform 1 0 33488 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1127_
timestamp 1676037725
transform 1 0 34224 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1128_
timestamp 1676037725
transform 1 0 34868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1129_
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1130_
timestamp 1676037725
transform 1 0 34868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1131_
timestamp 1676037725
transform 1 0 33304 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1132_
timestamp 1676037725
transform 1 0 34040 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1133_
timestamp 1676037725
transform 1 0 37444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 38732 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1676037725
transform 1 0 23368 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1676037725
transform 1 0 28612 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1676037725
transform 1 0 26036 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1676037725
transform 1 0 28612 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1676037725
transform 1 0 44160 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1676037725
transform 1 0 46828 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1676037725
transform 1 0 44160 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1676037725
transform 1 0 46828 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout411 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 55476 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout412 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 52072 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout413 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 30820 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout414
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout415
timestamp 1676037725
transform 1 0 45172 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout416
timestamp 1676037725
transform 1 0 44160 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout417
timestamp 1676037725
transform 1 0 47748 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout418
timestamp 1676037725
transform 1 0 52256 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout419
timestamp 1676037725
transform 1 0 47104 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout420 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 28428 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout421
timestamp 1676037725
transform 1 0 34868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout422
timestamp 1676037725
transform 1 0 46184 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout423
timestamp 1676037725
transform 1 0 46368 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout424
timestamp 1676037725
transform 1 0 30268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout425
timestamp 1676037725
transform 1 0 28704 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout426
timestamp 1676037725
transform 1 0 38640 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  fanout427 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 32936 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  fanout429
timestamp 1676037725
transform 1 0 14260 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout430
timestamp 1676037725
transform 1 0 37352 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  fanout431
timestamp 1676037725
transform 1 0 16836 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  fanout432 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 22632 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout433
timestamp 1676037725
transform 1 0 24564 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout434
timestamp 1676037725
transform 1 0 20700 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout435
timestamp 1676037725
transform 1 0 15548 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout436
timestamp 1676037725
transform 1 0 37444 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout437
timestamp 1676037725
transform 1 0 28520 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout438
timestamp 1676037725
transform 1 0 29716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout439
timestamp 1676037725
transform 1 0 28336 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout440
timestamp 1676037725
transform 1 0 32108 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout441
timestamp 1676037725
transform 1 0 15640 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout442
timestamp 1676037725
transform 1 0 17480 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout443
timestamp 1676037725
transform 1 0 12144 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout444
timestamp 1676037725
transform 1 0 19504 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout445
timestamp 1676037725
transform 1 0 28336 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout446
timestamp 1676037725
transform 1 0 29532 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout447
timestamp 1676037725
transform 1 0 24748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_12  fanout448
timestamp 1676037725
transform 1 0 27324 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  fanout449
timestamp 1676037725
transform 1 0 21988 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  fanout450
timestamp 1676037725
transform 1 0 10764 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  fanout451
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  fanout452
timestamp 1676037725
transform 1 0 25484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout453
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout454
timestamp 1676037725
transform 1 0 35604 0 -1 58752
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout455
timestamp 1676037725
transform 1 0 24564 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout456
timestamp 1676037725
transform 1 0 19504 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout457
timestamp 1676037725
transform 1 0 29716 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout458
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout459
timestamp 1676037725
transform 1 0 18400 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout460
timestamp 1676037725
transform 1 0 23184 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout461 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 -1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout462
timestamp 1676037725
transform 1 0 18216 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout463
timestamp 1676037725
transform 1 0 25576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout464
timestamp 1676037725
transform 1 0 17296 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout465
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout466
timestamp 1676037725
transform 1 0 19504 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout467
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout468
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout469
timestamp 1676037725
transform 1 0 8188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout470
timestamp 1676037725
transform 1 0 9476 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout471
timestamp 1676037725
transform 1 0 11684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout472
timestamp 1676037725
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout473
timestamp 1676037725
transform 1 0 13432 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout474
timestamp 1676037725
transform 1 0 14260 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout475
timestamp 1676037725
transform 1 0 21988 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  fanout476
timestamp 1676037725
transform 1 0 29716 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout477
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout478
timestamp 1676037725
transform 1 0 33304 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout479
timestamp 1676037725
transform 1 0 30820 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout480
timestamp 1676037725
transform 1 0 43700 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout481
timestamp 1676037725
transform 1 0 25024 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout482
timestamp 1676037725
transform 1 0 34500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout483
timestamp 1676037725
transform 1 0 28612 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout484
timestamp 1676037725
transform 1 0 34868 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout485
timestamp 1676037725
transform 1 0 42044 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout486
timestamp 1676037725
transform 1 0 45908 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout487
timestamp 1676037725
transform 1 0 47012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout488
timestamp 1676037725
transform 1 0 42872 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout489
timestamp 1676037725
transform 1 0 45264 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout490
timestamp 1676037725
transform 1 0 42688 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout491
timestamp 1676037725
transform 1 0 43240 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout492
timestamp 1676037725
transform 1 0 56488 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  hold1
timestamp 1676037725
transform 1 0 18584 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold2
timestamp 1676037725
transform 1 0 5704 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold3
timestamp 1676037725
transform 1 0 21160 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold4
timestamp 1676037725
transform 1 0 10304 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold5
timestamp 1676037725
transform 1 0 28612 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold6
timestamp 1676037725
transform 1 0 17756 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold7
timestamp 1676037725
transform 1 0 24288 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold8
timestamp 1676037725
transform 1 0 12788 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold9
timestamp 1676037725
transform 1 0 24288 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold10
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold11
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold12
timestamp 1676037725
transform 1 0 16100 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold13
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold14
timestamp 1676037725
transform 1 0 13432 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold15
timestamp 1676037725
transform 1 0 16836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold16
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold17
timestamp 1676037725
transform 1 0 21344 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold18
timestamp 1676037725
transform 1 0 8280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold19
timestamp 1676037725
transform 1 0 17848 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold20
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold21
timestamp 1676037725
transform 1 0 25576 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold22
timestamp 1676037725
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold23
timestamp 1676037725
transform 1 0 25760 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold24
timestamp 1676037725
transform 1 0 15272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold25
timestamp 1676037725
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold26
timestamp 1676037725
transform 1 0 29164 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold27
timestamp 1676037725
transform 1 0 16008 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold28
timestamp 1676037725
transform 1 0 15272 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold29
timestamp 1676037725
transform 1 0 23736 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold30
timestamp 1676037725
transform 1 0 18584 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold31
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold32
timestamp 1676037725
transform 1 0 23920 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold33
timestamp 1676037725
transform 1 0 17020 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold34
timestamp 1676037725
transform 1 0 16008 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold35
timestamp 1676037725
transform 1 0 20424 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold36
timestamp 1676037725
transform 1 0 18400 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold37
timestamp 1676037725
transform 1 0 23552 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold38
timestamp 1676037725
transform 1 0 19044 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold39
timestamp 1676037725
transform 1 0 17296 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold40
timestamp 1676037725
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold41
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold42
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold43
timestamp 1676037725
transform 1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold44
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold45
timestamp 1676037725
transform 1 0 6992 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold46
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold47
timestamp 1676037725
transform 1 0 18400 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold48
timestamp 1676037725
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold49
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold50
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold51
timestamp 1676037725
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold52
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold53
timestamp 1676037725
transform 1 0 20424 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold54
timestamp 1676037725
transform 1 0 17572 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold55
timestamp 1676037725
transform 1 0 23920 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold56
timestamp 1676037725
transform 1 0 10488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold57
timestamp 1676037725
transform 1 0 9844 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold58
timestamp 1676037725
transform 1 0 18492 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold59
timestamp 1676037725
transform 1 0 11960 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold60
timestamp 1676037725
transform 1 0 10580 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold61
timestamp 1676037725
transform 1 0 25576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold62
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold63
timestamp 1676037725
transform 1 0 5336 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold64
timestamp 1676037725
transform 1 0 6532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold65
timestamp 1676037725
transform 1 0 26312 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold66
timestamp 1676037725
transform 1 0 16008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold67
timestamp 1676037725
transform 1 0 10212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold68
timestamp 1676037725
transform 1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold69
timestamp 1676037725
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold70
timestamp 1676037725
transform 1 0 15272 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold71
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold72
timestamp 1676037725
transform 1 0 12420 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold73
timestamp 1676037725
transform 1 0 29900 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold74
timestamp 1676037725
transform 1 0 16560 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold75
timestamp 1676037725
transform 1 0 12052 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold76
timestamp 1676037725
transform 1 0 11960 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold77
timestamp 1676037725
transform 1 0 34776 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold78
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold79
timestamp 1676037725
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold80
timestamp 1676037725
transform 1 0 15824 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold81
timestamp 1676037725
transform 1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold82
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold83
timestamp 1676037725
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold84
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold85
timestamp 1676037725
transform 1 0 26220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold86
timestamp 1676037725
transform 1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold87
timestamp 1676037725
transform 1 0 12696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold88
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold89
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold90
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold91
timestamp 1676037725
transform 1 0 17112 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold92
timestamp 1676037725
transform 1 0 16376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold93
timestamp 1676037725
transform 1 0 29624 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold94
timestamp 1676037725
transform 1 0 18584 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold95
timestamp 1676037725
transform 1 0 14444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold96
timestamp 1676037725
transform 1 0 13432 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold97
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold98
timestamp 1676037725
transform 1 0 15640 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold99
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold100
timestamp 1676037725
transform 1 0 13984 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold101
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold102
timestamp 1676037725
transform 1 0 14904 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold103
timestamp 1676037725
transform 1 0 8648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold104
timestamp 1676037725
transform 1 0 9660 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold105
timestamp 1676037725
transform 1 0 32384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold106
timestamp 1676037725
transform 1 0 15824 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold107
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold108
timestamp 1676037725
transform 1 0 26312 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold109
timestamp 1676037725
transform 1 0 22908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold110
timestamp 1676037725
transform 1 0 19320 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold111
timestamp 1676037725
transform 1 0 17664 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold112
timestamp 1676037725
transform 1 0 31372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold113
timestamp 1676037725
transform 1 0 22172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold114
timestamp 1676037725
transform 1 0 16560 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold115
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold116
timestamp 1676037725
transform 1 0 26312 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold117
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold118
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold119
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold120
timestamp 1676037725
transform 1 0 23736 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold121
timestamp 1676037725
transform 1 0 25852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold122
timestamp 1676037725
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold123
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold124
timestamp 1676037725
transform 1 0 20148 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold125
timestamp 1676037725
transform 1 0 22724 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold126
timestamp 1676037725
transform 1 0 19228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold127
timestamp 1676037725
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold128
timestamp 1676037725
transform 1 0 16008 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold129
timestamp 1676037725
transform 1 0 25944 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold130
timestamp 1676037725
transform 1 0 14444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold131
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold132
timestamp 1676037725
transform 1 0 26404 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold133
timestamp 1676037725
transform 1 0 16008 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold134
timestamp 1676037725
transform 1 0 12420 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold135
timestamp 1676037725
transform 1 0 30544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold136
timestamp 1676037725
transform 1 0 17940 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold137
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold138
timestamp 1676037725
transform 1 0 20332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold139
timestamp 1676037725
transform 1 0 19688 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold140
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold141
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold142
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold143
timestamp 1676037725
transform 1 0 20884 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold144
timestamp 1676037725
transform 1 0 16008 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1676037725
transform 1 0 40020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1676037725
transform 1 0 40480 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1676037725
transform 1 0 41124 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1676037725
transform 1 0 45172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1676037725
transform 1 0 44988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1676037725
transform 1 0 41308 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1676037725
transform 1 0 41584 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform 1 0 42596 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1676037725
transform 1 0 44252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform 1 0 46920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1676037725
transform 1 0 45172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1676037725
transform 1 0 41768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform 1 0 43332 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1676037725
transform 1 0 44988 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1676037725
transform 1 0 44068 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1676037725
transform 1 0 45172 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1676037725
transform 1 0 44804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1676037725
transform 1 0 41308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1676037725
transform 1 0 40756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1676037725
transform 1 0 38548 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1676037725
transform 1 0 40388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1676037725
transform 1 0 41492 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1676037725
transform 1 0 39560 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1676037725
transform 1 0 44252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1676037725
transform 1 0 54096 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1676037725
transform 1 0 54648 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input30
timestamp 1676037725
transform 1 0 55476 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input31
timestamp 1676037725
transform 1 0 56396 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1676037725
transform 1 0 56856 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1676037725
transform 1 0 58052 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input34
timestamp 1676037725
transform 1 0 57868 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1676037725
transform 1 0 57132 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1676037725
transform 1 0 46460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 1676037725
transform 1 0 48484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1676037725
transform 1 0 50324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 1676037725
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1676037725
transform 1 0 49220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input42
timestamp 1676037725
transform 1 0 49588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1676037725
transform 1 0 50508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 50324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1676037725
transform 1 0 51796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1676037725
transform 1 0 45908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1676037725
transform 1 0 51244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1676037725
transform 1 0 51060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1676037725
transform 1 0 51980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1676037725
transform 1 0 51796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1676037725
transform 1 0 52900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1676037725
transform 1 0 52532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1676037725
transform 1 0 52072 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1676037725
transform 1 0 47748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input57
timestamp 1676037725
transform 1 0 46000 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input58
timestamp 1676037725
transform 1 0 46276 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input59
timestamp 1676037725
transform 1 0 47748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input60
timestamp 1676037725
transform 1 0 46828 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input61
timestamp 1676037725
transform 1 0 47748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1676037725
transform 1 0 48668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1676037725
transform 1 0 13432 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1676037725
transform 1 0 20424 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1676037725
transform 1 0 21160 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input66
timestamp 1676037725
transform 1 0 22264 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input67
timestamp 1676037725
transform 1 0 23644 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 23736 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1676037725
transform 1 0 24472 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1676037725
transform 1 0 25208 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1676037725
transform 1 0 26128 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input72
timestamp 1676037725
transform 1 0 27140 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1676037725
transform 1 0 27416 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1676037725
transform 1 0 14168 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input75
timestamp 1676037725
transform 1 0 28152 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1676037725
transform 1 0 28888 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input77
timestamp 1676037725
transform 1 0 29716 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1676037725
transform 1 0 30360 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input79
timestamp 1676037725
transform 1 0 31096 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1676037725
transform 1 0 32292 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1676037725
transform 1 0 33212 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input82
timestamp 1676037725
transform 1 0 14904 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1676037725
transform 1 0 15640 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1676037725
transform 1 0 16008 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input85
timestamp 1676037725
transform 1 0 17112 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1676037725
transform 1 0 17848 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1676037725
transform 1 0 18584 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp 1676037725
transform 1 0 19320 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1676037725
transform 1 0 19688 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input90
timestamp 1676037725
transform 1 0 1564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input91
timestamp 1676037725
transform 1 0 1564 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input92
timestamp 1676037725
transform 1 0 1564 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1676037725
transform 1 0 1564 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input94
timestamp 1676037725
transform 1 0 1564 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input95
timestamp 1676037725
transform 1 0 1564 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input96
timestamp 1676037725
transform 1 0 1564 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input97
timestamp 1676037725
transform 1 0 1564 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1676037725
transform 1 0 1564 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1676037725
transform 1 0 1564 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input100
timestamp 1676037725
transform 1 0 1564 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1676037725
transform 1 0 1564 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input102
timestamp 1676037725
transform 1 0 1564 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1676037725
transform 1 0 1564 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input104
timestamp 1676037725
transform 1 0 1564 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input105
timestamp 1676037725
transform 1 0 1564 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input106
timestamp 1676037725
transform 1 0 1564 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input107
timestamp 1676037725
transform 1 0 1564 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input108
timestamp 1676037725
transform 1 0 1564 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input109
timestamp 1676037725
transform 1 0 2760 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1676037725
transform 1 0 1564 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input111
timestamp 1676037725
transform 1 0 1564 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input112
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input113
timestamp 1676037725
transform 1 0 1564 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input114
timestamp 1676037725
transform 1 0 1564 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1676037725
transform 1 0 1564 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1676037725
transform 1 0 1564 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input117
timestamp 1676037725
transform 1 0 1564 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 1676037725
transform 1 0 33948 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1676037725
transform 1 0 41492 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1676037725
transform 1 0 41400 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input121
timestamp 1676037725
transform 1 0 42596 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input122
timestamp 1676037725
transform 1 0 43516 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input123
timestamp 1676037725
transform 1 0 44252 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input124
timestamp 1676037725
transform 1 0 45172 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input125
timestamp 1676037725
transform 1 0 45908 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input126
timestamp 1676037725
transform 1 0 46644 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input127
timestamp 1676037725
transform 1 0 46552 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input128
timestamp 1676037725
transform 1 0 47748 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input129
timestamp 1676037725
transform 1 0 34868 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1676037725
transform 1 0 48484 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input131
timestamp 1676037725
transform 1 0 49220 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input132
timestamp 1676037725
transform 1 0 50324 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input133
timestamp 1676037725
transform 1 0 50232 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input134
timestamp 1676037725
transform 1 0 51244 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input135
timestamp 1676037725
transform 1 0 51980 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input136
timestamp 1676037725
transform 1 0 52900 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input137
timestamp 1676037725
transform 1 0 35604 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input138
timestamp 1676037725
transform 1 0 36340 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input139
timestamp 1676037725
transform 1 0 36248 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input140
timestamp 1676037725
transform 1 0 37444 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input141
timestamp 1676037725
transform 1 0 38180 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input142
timestamp 1676037725
transform 1 0 38916 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input143
timestamp 1676037725
transform 1 0 40020 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input144
timestamp 1676037725
transform 1 0 40756 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input145
timestamp 1676037725
transform 1 0 58052 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input146
timestamp 1676037725
transform 1 0 56120 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input147
timestamp 1676037725
transform 1 0 57224 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input148
timestamp 1676037725
transform 1 0 57868 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input149
timestamp 1676037725
transform 1 0 57868 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input150
timestamp 1676037725
transform 1 0 57868 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input151
timestamp 1676037725
transform 1 0 58052 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input152
timestamp 1676037725
transform 1 0 58052 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1676037725
transform 1 0 58052 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input154
timestamp 1676037725
transform 1 0 57132 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input155
timestamp 1676037725
transform 1 0 56396 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1676037725
transform 1 0 55384 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input157
timestamp 1676037725
transform 1 0 6624 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input158
timestamp 1676037725
transform 1 0 7544 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input159
timestamp 1676037725
transform 1 0 8280 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input160
timestamp 1676037725
transform 1 0 9016 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input161
timestamp 1676037725
transform 1 0 9384 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input162
timestamp 1676037725
transform 1 0 10120 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input163
timestamp 1676037725
transform 1 0 10856 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input164
timestamp 1676037725
transform 1 0 11960 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input165
timestamp 1676037725
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input166
timestamp 1676037725
transform 1 0 1564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input167
timestamp 1676037725
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input168
timestamp 1676037725
transform 1 0 1564 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input169
timestamp 1676037725
transform 1 0 1564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input170
timestamp 1676037725
transform 1 0 1564 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input171
timestamp 1676037725
transform 1 0 1564 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input172
timestamp 1676037725
transform 1 0 1564 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input173
timestamp 1676037725
transform 1 0 1564 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input174
timestamp 1676037725
transform 1 0 1564 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input175
timestamp 1676037725
transform 1 0 2484 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input176
timestamp 1676037725
transform 1 0 2484 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input177
timestamp 1676037725
transform 1 0 3128 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input178
timestamp 1676037725
transform 1 0 3864 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input179
timestamp 1676037725
transform 1 0 4232 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input180
timestamp 1676037725
transform 1 0 4968 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input181
timestamp 1676037725
transform 1 0 5704 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input182
timestamp 1676037725
transform 1 0 36340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input183
timestamp 1676037725
transform 1 0 37168 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input184
timestamp 1676037725
transform 1 0 39836 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input185
timestamp 1676037725
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input186
timestamp 1676037725
transform 1 0 1564 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input187
timestamp 1676037725
transform 1 0 1564 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input188
timestamp 1676037725
transform 1 0 1564 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input189
timestamp 1676037725
transform 1 0 1564 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input190
timestamp 1676037725
transform 1 0 1564 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input191
timestamp 1676037725
transform 1 0 1564 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input192
timestamp 1676037725
transform 1 0 1564 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input193
timestamp 1676037725
transform 1 0 1564 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input194
timestamp 1676037725
transform 1 0 52900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input195
timestamp 1676037725
transform 1 0 52900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input196
timestamp 1676037725
transform 1 0 54004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input197
timestamp 1676037725
transform 1 0 53636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input198
timestamp 1676037725
transform 1 0 53820 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input199
timestamp 1676037725
transform 1 0 54004 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input200
timestamp 1676037725
transform 1 0 54924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input201
timestamp 1676037725
transform 1 0 54556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input202
timestamp 1676037725
transform 1 0 55476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input203
timestamp 1676037725
transform 1 0 55476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input204
timestamp 1676037725
transform 1 0 55844 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input205
timestamp 1676037725
transform 1 0 3128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input206
timestamp 1676037725
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input207
timestamp 1676037725
transform 1 0 4968 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input208
timestamp 1676037725
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input209
timestamp 1676037725
transform 1 0 6532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input210
timestamp 1676037725
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input211
timestamp 1676037725
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input212
timestamp 1676037725
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input213
timestamp 1676037725
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input214
timestamp 1676037725
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input215
timestamp 1676037725
transform 1 0 8280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input216
timestamp 1676037725
transform 1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input217
timestamp 1676037725
transform 1 0 6900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input218
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input219
timestamp 1676037725
transform 1 0 7636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input220
timestamp 1676037725
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input221
timestamp 1676037725
transform 1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input222
timestamp 1676037725
transform 1 0 10856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input223
timestamp 1676037725
transform 1 0 11684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input224
timestamp 1676037725
transform 1 0 12328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input225
timestamp 1676037725
transform 1 0 11684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input226
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input227
timestamp 1676037725
transform 1 0 12420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input228
timestamp 1676037725
transform 1 0 11776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input229
timestamp 1676037725
transform 1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input230
timestamp 1676037725
transform 1 0 14260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input231
timestamp 1676037725
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input232
timestamp 1676037725
transform 1 0 10856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input233
timestamp 1676037725
transform 1 0 12328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input234
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input235
timestamp 1676037725
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input236
timestamp 1676037725
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input237
timestamp 1676037725
transform 1 0 4968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input238
timestamp 1676037725
transform 1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input239
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input240
timestamp 1676037725
transform 1 0 53268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input241
timestamp 1676037725
transform 1 0 12696 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input242
timestamp 1676037725
transform 1 0 1564 0 1 60928
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  input243
timestamp 1676037725
transform 1 0 53176 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input244
timestamp 1676037725
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input245
timestamp 1676037725
transform 1 0 58052 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input246
timestamp 1676037725
transform 1 0 57868 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input247
timestamp 1676037725
transform 1 0 56948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input248
timestamp 1676037725
transform 1 0 57868 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input249
timestamp 1676037725
transform 1 0 58052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input250
timestamp 1676037725
transform 1 0 58052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input251
timestamp 1676037725
transform 1 0 58052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input252
timestamp 1676037725
transform 1 0 58052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input253
timestamp 1676037725
transform 1 0 58052 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input254
timestamp 1676037725
transform 1 0 58052 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input255
timestamp 1676037725
transform 1 0 57868 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input256
timestamp 1676037725
transform 1 0 56948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input257
timestamp 1676037725
transform 1 0 58052 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input258
timestamp 1676037725
transform 1 0 56948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input259
timestamp 1676037725
transform 1 0 58052 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input260
timestamp 1676037725
transform 1 0 57868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input261
timestamp 1676037725
transform 1 0 58052 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input262
timestamp 1676037725
transform 1 0 58052 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input263
timestamp 1676037725
transform 1 0 56948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input264
timestamp 1676037725
transform 1 0 57868 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input265
timestamp 1676037725
transform 1 0 56948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input266
timestamp 1676037725
transform 1 0 57868 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input267
timestamp 1676037725
transform 1 0 58052 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input268
timestamp 1676037725
transform 1 0 58052 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input269
timestamp 1676037725
transform 1 0 57868 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input270
timestamp 1676037725
transform 1 0 56120 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input271
timestamp 1676037725
transform 1 0 56948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input272
timestamp 1676037725
transform 1 0 57040 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input273
timestamp 1676037725
transform 1 0 56948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input274
timestamp 1676037725
transform 1 0 57868 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input275
timestamp 1676037725
transform 1 0 56948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input276
timestamp 1676037725
transform 1 0 57868 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input277
timestamp 1676037725
transform 1 0 57868 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input278
timestamp 1676037725
transform 1 0 58052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input279
timestamp 1676037725
transform 1 0 58052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  max_cap428
timestamp 1676037725
transform 1 0 16836 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  multiplexer_493 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_494
timestamp 1676037725
transform 1 0 26312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_495
timestamp 1676037725
transform 1 0 26312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_496
timestamp 1676037725
transform 1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_497
timestamp 1676037725
transform 1 0 17664 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_498
timestamp 1676037725
transform 1 0 16100 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_499
timestamp 1676037725
transform 1 0 17020 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_500
timestamp 1676037725
transform 1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_501
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_502
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_503
timestamp 1676037725
transform 1 0 58144 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_504
timestamp 1676037725
transform 1 0 58144 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_505
timestamp 1676037725
transform 1 0 58144 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_506
timestamp 1676037725
transform 1 0 58144 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_507
timestamp 1676037725
transform 1 0 26956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_508
timestamp 1676037725
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_509
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_510
timestamp 1676037725
transform 1 0 29072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_511
timestamp 1676037725
transform 1 0 28980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_512
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output280
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output281
timestamp 1676037725
transform 1 0 1564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output282
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output283
timestamp 1676037725
transform 1 0 1564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output284
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output285
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output286
timestamp 1676037725
transform 1 0 1564 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output287
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output288
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output289
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output290
timestamp 1676037725
transform 1 0 1564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output291
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output292
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output293
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output294
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output295
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output296
timestamp 1676037725
transform 1 0 1564 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output297
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output298
timestamp 1676037725
transform 1 0 1564 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output299
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output300
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output301
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output302
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output303
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output304
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output305
timestamp 1676037725
transform 1 0 1564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output306
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output307
timestamp 1676037725
transform 1 0 1564 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output308
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output309
timestamp 1676037725
transform 1 0 25208 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output310
timestamp 1676037725
transform 1 0 26128 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output311
timestamp 1676037725
transform 1 0 26128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output312
timestamp 1676037725
transform 1 0 27508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output313
timestamp 1676037725
transform 1 0 27784 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output314
timestamp 1676037725
transform 1 0 29716 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output315
timestamp 1676037725
transform 1 0 28704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output316
timestamp 1676037725
transform 1 0 30268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output317
timestamp 1676037725
transform 1 0 30176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output318
timestamp 1676037725
transform 1 0 30820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output319
timestamp 1676037725
transform 1 0 31096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output320
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output321
timestamp 1676037725
transform 1 0 32292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output322
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output323
timestamp 1676037725
transform 1 0 34868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output324
timestamp 1676037725
transform 1 0 35788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output325
timestamp 1676037725
transform 1 0 33488 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output326
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output327
timestamp 1676037725
transform 1 0 34868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output328
timestamp 1676037725
transform 1 0 34408 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output329
timestamp 1676037725
transform 1 0 36340 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output330
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output331
timestamp 1676037725
transform 1 0 35328 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output332
timestamp 1676037725
transform 1 0 36248 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output333
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output334
timestamp 1676037725
transform 1 0 38640 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output335
timestamp 1676037725
transform 1 0 40020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output336
timestamp 1676037725
transform 1 0 35788 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output337
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output338
timestamp 1676037725
transform 1 0 17480 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output339
timestamp 1676037725
transform 1 0 17020 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output340
timestamp 1676037725
transform 1 0 18676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output341
timestamp 1676037725
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output342
timestamp 1676037725
transform 1 0 18400 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output343
timestamp 1676037725
transform 1 0 15824 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output344
timestamp 1676037725
transform 1 0 17204 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output345
timestamp 1676037725
transform 1 0 17940 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output346
timestamp 1676037725
transform 1 0 15824 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output347
timestamp 1676037725
transform 1 0 15364 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output348
timestamp 1676037725
transform 1 0 16928 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output349
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output350
timestamp 1676037725
transform 1 0 20976 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output351
timestamp 1676037725
transform 1 0 17848 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output352
timestamp 1676037725
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output353
timestamp 1676037725
transform 1 0 18768 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output354
timestamp 1676037725
transform 1 0 18400 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output355
timestamp 1676037725
transform 1 0 22540 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output356
timestamp 1676037725
transform 1 0 22356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output357
timestamp 1676037725
transform 1 0 21712 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output358
timestamp 1676037725
transform 1 0 13984 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output359
timestamp 1676037725
transform 1 0 22448 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output360
timestamp 1676037725
transform 1 0 23644 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output361
timestamp 1676037725
transform 1 0 25760 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output362
timestamp 1676037725
transform 1 0 22356 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output363
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output364
timestamp 1676037725
transform 1 0 25208 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output365
timestamp 1676037725
transform 1 0 23552 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output366
timestamp 1676037725
transform 1 0 25208 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output367
timestamp 1676037725
transform 1 0 13248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output368
timestamp 1676037725
transform 1 0 14904 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output369
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output370
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output371
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output372
timestamp 1676037725
transform 1 0 1564 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output373
timestamp 1676037725
transform 1 0 1564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output374
timestamp 1676037725
transform 1 0 1564 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output375
timestamp 1676037725
transform 1 0 1564 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output376
timestamp 1676037725
transform 1 0 1564 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output377
timestamp 1676037725
transform 1 0 1564 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output378
timestamp 1676037725
transform 1 0 1564 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output379
timestamp 1676037725
transform 1 0 1564 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output380
timestamp 1676037725
transform 1 0 1564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output381
timestamp 1676037725
transform 1 0 1564 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output382
timestamp 1676037725
transform 1 0 57040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output383
timestamp 1676037725
transform 1 0 56948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output384
timestamp 1676037725
transform 1 0 57868 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output385
timestamp 1676037725
transform 1 0 57868 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output386
timestamp 1676037725
transform 1 0 57868 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output387
timestamp 1676037725
transform 1 0 57868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output388
timestamp 1676037725
transform 1 0 57868 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output389
timestamp 1676037725
transform 1 0 57868 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output390
timestamp 1676037725
transform 1 0 57868 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output391
timestamp 1676037725
transform 1 0 57868 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output392
timestamp 1676037725
transform 1 0 57868 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output393
timestamp 1676037725
transform 1 0 57868 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output394
timestamp 1676037725
transform 1 0 57868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output395
timestamp 1676037725
transform 1 0 57868 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output396
timestamp 1676037725
transform 1 0 57868 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output397
timestamp 1676037725
transform 1 0 56948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output398
timestamp 1676037725
transform 1 0 57868 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output399
timestamp 1676037725
transform 1 0 56948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output400
timestamp 1676037725
transform 1 0 57868 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output401
timestamp 1676037725
transform 1 0 57868 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output402
timestamp 1676037725
transform 1 0 57868 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output403
timestamp 1676037725
transform 1 0 57040 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output404
timestamp 1676037725
transform 1 0 57868 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output405
timestamp 1676037725
transform 1 0 57868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output406
timestamp 1676037725
transform 1 0 57868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output407
timestamp 1676037725
transform 1 0 57868 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output408
timestamp 1676037725
transform 1 0 57040 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output409
timestamp 1676037725
transform 1 0 56948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output410
timestamp 1676037725
transform 1 0 57868 0 1 20672
box -38 -48 590 592
<< labels >>
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 design_clk_o
port 0 nsew signal tristate
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 dsi_all[0]
port 1 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 dsi_all[10]
port 2 nsew signal tristate
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 dsi_all[11]
port 3 nsew signal tristate
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 dsi_all[12]
port 4 nsew signal tristate
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 dsi_all[13]
port 5 nsew signal tristate
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 dsi_all[14]
port 6 nsew signal tristate
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 dsi_all[15]
port 7 nsew signal tristate
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 dsi_all[16]
port 8 nsew signal tristate
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 dsi_all[17]
port 9 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 dsi_all[18]
port 10 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 dsi_all[19]
port 11 nsew signal tristate
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 dsi_all[1]
port 12 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 dsi_all[20]
port 13 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 dsi_all[21]
port 14 nsew signal tristate
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 dsi_all[22]
port 15 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 dsi_all[23]
port 16 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 dsi_all[24]
port 17 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 dsi_all[25]
port 18 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 dsi_all[26]
port 19 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 dsi_all[27]
port 20 nsew signal tristate
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 dsi_all[2]
port 21 nsew signal tristate
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 dsi_all[3]
port 22 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 dsi_all[4]
port 23 nsew signal tristate
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 dsi_all[5]
port 24 nsew signal tristate
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 dsi_all[6]
port 25 nsew signal tristate
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 dsi_all[7]
port 26 nsew signal tristate
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 dsi_all[8]
port 27 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 dsi_all[9]
port 28 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 dso_6502[0]
port 29 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 dso_6502[10]
port 30 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 dso_6502[11]
port 31 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 dso_6502[12]
port 32 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 dso_6502[13]
port 33 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 dso_6502[14]
port 34 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 dso_6502[15]
port 35 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 dso_6502[16]
port 36 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 dso_6502[17]
port 37 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 dso_6502[18]
port 38 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 dso_6502[19]
port 39 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 dso_6502[1]
port 40 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 dso_6502[20]
port 41 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 dso_6502[21]
port 42 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 dso_6502[22]
port 43 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 dso_6502[23]
port 44 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 dso_6502[24]
port 45 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 dso_6502[25]
port 46 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 dso_6502[26]
port 47 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 dso_6502[2]
port 48 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 dso_6502[3]
port 49 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 dso_6502[4]
port 50 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 dso_6502[5]
port 51 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 dso_6502[6]
port 52 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 dso_6502[7]
port 53 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 dso_6502[8]
port 54 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 dso_6502[9]
port 55 nsew signal input
flabel metal2 s 53838 63200 53894 64000 0 FreeSans 224 90 0 0 dso_LCD[0]
port 56 nsew signal input
flabel metal2 s 54574 63200 54630 64000 0 FreeSans 224 90 0 0 dso_LCD[1]
port 57 nsew signal input
flabel metal2 s 55310 63200 55366 64000 0 FreeSans 224 90 0 0 dso_LCD[2]
port 58 nsew signal input
flabel metal2 s 56046 63200 56102 64000 0 FreeSans 224 90 0 0 dso_LCD[3]
port 59 nsew signal input
flabel metal2 s 56782 63200 56838 64000 0 FreeSans 224 90 0 0 dso_LCD[4]
port 60 nsew signal input
flabel metal2 s 57518 63200 57574 64000 0 FreeSans 224 90 0 0 dso_LCD[5]
port 61 nsew signal input
flabel metal2 s 58254 63200 58310 64000 0 FreeSans 224 90 0 0 dso_LCD[6]
port 62 nsew signal input
flabel metal2 s 58990 63200 59046 64000 0 FreeSans 224 90 0 0 dso_LCD[7]
port 63 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 dso_as1802[0]
port 64 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 dso_as1802[10]
port 65 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 dso_as1802[11]
port 66 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 dso_as1802[12]
port 67 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 dso_as1802[13]
port 68 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 dso_as1802[14]
port 69 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 dso_as1802[15]
port 70 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 dso_as1802[16]
port 71 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 dso_as1802[17]
port 72 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 dso_as1802[18]
port 73 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 dso_as1802[19]
port 74 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 dso_as1802[1]
port 75 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 dso_as1802[20]
port 76 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 dso_as1802[21]
port 77 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 dso_as1802[22]
port 78 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 dso_as1802[23]
port 79 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 dso_as1802[24]
port 80 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 dso_as1802[25]
port 81 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 dso_as1802[26]
port 82 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 dso_as1802[2]
port 83 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 dso_as1802[3]
port 84 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 dso_as1802[4]
port 85 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 dso_as1802[5]
port 86 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 dso_as1802[6]
port 87 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 dso_as1802[7]
port 88 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 dso_as1802[8]
port 89 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 dso_as1802[9]
port 90 nsew signal input
flabel metal2 s 13358 63200 13414 64000 0 FreeSans 224 90 0 0 dso_as2650[0]
port 91 nsew signal input
flabel metal2 s 20718 63200 20774 64000 0 FreeSans 224 90 0 0 dso_as2650[10]
port 92 nsew signal input
flabel metal2 s 21454 63200 21510 64000 0 FreeSans 224 90 0 0 dso_as2650[11]
port 93 nsew signal input
flabel metal2 s 22190 63200 22246 64000 0 FreeSans 224 90 0 0 dso_as2650[12]
port 94 nsew signal input
flabel metal2 s 22926 63200 22982 64000 0 FreeSans 224 90 0 0 dso_as2650[13]
port 95 nsew signal input
flabel metal2 s 23662 63200 23718 64000 0 FreeSans 224 90 0 0 dso_as2650[14]
port 96 nsew signal input
flabel metal2 s 24398 63200 24454 64000 0 FreeSans 224 90 0 0 dso_as2650[15]
port 97 nsew signal input
flabel metal2 s 25134 63200 25190 64000 0 FreeSans 224 90 0 0 dso_as2650[16]
port 98 nsew signal input
flabel metal2 s 25870 63200 25926 64000 0 FreeSans 224 90 0 0 dso_as2650[17]
port 99 nsew signal input
flabel metal2 s 26606 63200 26662 64000 0 FreeSans 224 90 0 0 dso_as2650[18]
port 100 nsew signal input
flabel metal2 s 27342 63200 27398 64000 0 FreeSans 224 90 0 0 dso_as2650[19]
port 101 nsew signal input
flabel metal2 s 14094 63200 14150 64000 0 FreeSans 224 90 0 0 dso_as2650[1]
port 102 nsew signal input
flabel metal2 s 28078 63200 28134 64000 0 FreeSans 224 90 0 0 dso_as2650[20]
port 103 nsew signal input
flabel metal2 s 28814 63200 28870 64000 0 FreeSans 224 90 0 0 dso_as2650[21]
port 104 nsew signal input
flabel metal2 s 29550 63200 29606 64000 0 FreeSans 224 90 0 0 dso_as2650[22]
port 105 nsew signal input
flabel metal2 s 30286 63200 30342 64000 0 FreeSans 224 90 0 0 dso_as2650[23]
port 106 nsew signal input
flabel metal2 s 31022 63200 31078 64000 0 FreeSans 224 90 0 0 dso_as2650[24]
port 107 nsew signal input
flabel metal2 s 31758 63200 31814 64000 0 FreeSans 224 90 0 0 dso_as2650[25]
port 108 nsew signal input
flabel metal2 s 32494 63200 32550 64000 0 FreeSans 224 90 0 0 dso_as2650[26]
port 109 nsew signal input
flabel metal2 s 14830 63200 14886 64000 0 FreeSans 224 90 0 0 dso_as2650[2]
port 110 nsew signal input
flabel metal2 s 15566 63200 15622 64000 0 FreeSans 224 90 0 0 dso_as2650[3]
port 111 nsew signal input
flabel metal2 s 16302 63200 16358 64000 0 FreeSans 224 90 0 0 dso_as2650[4]
port 112 nsew signal input
flabel metal2 s 17038 63200 17094 64000 0 FreeSans 224 90 0 0 dso_as2650[5]
port 113 nsew signal input
flabel metal2 s 17774 63200 17830 64000 0 FreeSans 224 90 0 0 dso_as2650[6]
port 114 nsew signal input
flabel metal2 s 18510 63200 18566 64000 0 FreeSans 224 90 0 0 dso_as2650[7]
port 115 nsew signal input
flabel metal2 s 19246 63200 19302 64000 0 FreeSans 224 90 0 0 dso_as2650[8]
port 116 nsew signal input
flabel metal2 s 19982 63200 20038 64000 0 FreeSans 224 90 0 0 dso_as2650[9]
port 117 nsew signal input
flabel metal3 s 0 42712 800 42832 0 FreeSans 480 0 0 0 dso_as512512512[0]
port 118 nsew signal input
flabel metal3 s 0 49512 800 49632 0 FreeSans 480 0 0 0 dso_as512512512[10]
port 119 nsew signal input
flabel metal3 s 0 50192 800 50312 0 FreeSans 480 0 0 0 dso_as512512512[11]
port 120 nsew signal input
flabel metal3 s 0 50872 800 50992 0 FreeSans 480 0 0 0 dso_as512512512[12]
port 121 nsew signal input
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 dso_as512512512[13]
port 122 nsew signal input
flabel metal3 s 0 52232 800 52352 0 FreeSans 480 0 0 0 dso_as512512512[14]
port 123 nsew signal input
flabel metal3 s 0 52912 800 53032 0 FreeSans 480 0 0 0 dso_as512512512[15]
port 124 nsew signal input
flabel metal3 s 0 53592 800 53712 0 FreeSans 480 0 0 0 dso_as512512512[16]
port 125 nsew signal input
flabel metal3 s 0 54272 800 54392 0 FreeSans 480 0 0 0 dso_as512512512[17]
port 126 nsew signal input
flabel metal3 s 0 54952 800 55072 0 FreeSans 480 0 0 0 dso_as512512512[18]
port 127 nsew signal input
flabel metal3 s 0 55632 800 55752 0 FreeSans 480 0 0 0 dso_as512512512[19]
port 128 nsew signal input
flabel metal3 s 0 43392 800 43512 0 FreeSans 480 0 0 0 dso_as512512512[1]
port 129 nsew signal input
flabel metal3 s 0 56312 800 56432 0 FreeSans 480 0 0 0 dso_as512512512[20]
port 130 nsew signal input
flabel metal3 s 0 56992 800 57112 0 FreeSans 480 0 0 0 dso_as512512512[21]
port 131 nsew signal input
flabel metal3 s 0 57672 800 57792 0 FreeSans 480 0 0 0 dso_as512512512[22]
port 132 nsew signal input
flabel metal3 s 0 58352 800 58472 0 FreeSans 480 0 0 0 dso_as512512512[23]
port 133 nsew signal input
flabel metal3 s 0 59032 800 59152 0 FreeSans 480 0 0 0 dso_as512512512[24]
port 134 nsew signal input
flabel metal3 s 0 59712 800 59832 0 FreeSans 480 0 0 0 dso_as512512512[25]
port 135 nsew signal input
flabel metal3 s 0 60392 800 60512 0 FreeSans 480 0 0 0 dso_as512512512[26]
port 136 nsew signal input
flabel metal3 s 0 61072 800 61192 0 FreeSans 480 0 0 0 dso_as512512512[27]
port 137 nsew signal input
flabel metal3 s 0 44072 800 44192 0 FreeSans 480 0 0 0 dso_as512512512[2]
port 138 nsew signal input
flabel metal3 s 0 44752 800 44872 0 FreeSans 480 0 0 0 dso_as512512512[3]
port 139 nsew signal input
flabel metal3 s 0 45432 800 45552 0 FreeSans 480 0 0 0 dso_as512512512[4]
port 140 nsew signal input
flabel metal3 s 0 46112 800 46232 0 FreeSans 480 0 0 0 dso_as512512512[5]
port 141 nsew signal input
flabel metal3 s 0 46792 800 46912 0 FreeSans 480 0 0 0 dso_as512512512[6]
port 142 nsew signal input
flabel metal3 s 0 47472 800 47592 0 FreeSans 480 0 0 0 dso_as512512512[7]
port 143 nsew signal input
flabel metal3 s 0 48152 800 48272 0 FreeSans 480 0 0 0 dso_as512512512[8]
port 144 nsew signal input
flabel metal3 s 0 48832 800 48952 0 FreeSans 480 0 0 0 dso_as512512512[9]
port 145 nsew signal input
flabel metal2 s 33230 63200 33286 64000 0 FreeSans 224 90 0 0 dso_as5401[0]
port 146 nsew signal input
flabel metal2 s 40590 63200 40646 64000 0 FreeSans 224 90 0 0 dso_as5401[10]
port 147 nsew signal input
flabel metal2 s 41326 63200 41382 64000 0 FreeSans 224 90 0 0 dso_as5401[11]
port 148 nsew signal input
flabel metal2 s 42062 63200 42118 64000 0 FreeSans 224 90 0 0 dso_as5401[12]
port 149 nsew signal input
flabel metal2 s 42798 63200 42854 64000 0 FreeSans 224 90 0 0 dso_as5401[13]
port 150 nsew signal input
flabel metal2 s 43534 63200 43590 64000 0 FreeSans 224 90 0 0 dso_as5401[14]
port 151 nsew signal input
flabel metal2 s 44270 63200 44326 64000 0 FreeSans 224 90 0 0 dso_as5401[15]
port 152 nsew signal input
flabel metal2 s 45006 63200 45062 64000 0 FreeSans 224 90 0 0 dso_as5401[16]
port 153 nsew signal input
flabel metal2 s 45742 63200 45798 64000 0 FreeSans 224 90 0 0 dso_as5401[17]
port 154 nsew signal input
flabel metal2 s 46478 63200 46534 64000 0 FreeSans 224 90 0 0 dso_as5401[18]
port 155 nsew signal input
flabel metal2 s 47214 63200 47270 64000 0 FreeSans 224 90 0 0 dso_as5401[19]
port 156 nsew signal input
flabel metal2 s 33966 63200 34022 64000 0 FreeSans 224 90 0 0 dso_as5401[1]
port 157 nsew signal input
flabel metal2 s 47950 63200 48006 64000 0 FreeSans 224 90 0 0 dso_as5401[20]
port 158 nsew signal input
flabel metal2 s 48686 63200 48742 64000 0 FreeSans 224 90 0 0 dso_as5401[21]
port 159 nsew signal input
flabel metal2 s 49422 63200 49478 64000 0 FreeSans 224 90 0 0 dso_as5401[22]
port 160 nsew signal input
flabel metal2 s 50158 63200 50214 64000 0 FreeSans 224 90 0 0 dso_as5401[23]
port 161 nsew signal input
flabel metal2 s 50894 63200 50950 64000 0 FreeSans 224 90 0 0 dso_as5401[24]
port 162 nsew signal input
flabel metal2 s 51630 63200 51686 64000 0 FreeSans 224 90 0 0 dso_as5401[25]
port 163 nsew signal input
flabel metal2 s 52366 63200 52422 64000 0 FreeSans 224 90 0 0 dso_as5401[26]
port 164 nsew signal input
flabel metal2 s 34702 63200 34758 64000 0 FreeSans 224 90 0 0 dso_as5401[2]
port 165 nsew signal input
flabel metal2 s 35438 63200 35494 64000 0 FreeSans 224 90 0 0 dso_as5401[3]
port 166 nsew signal input
flabel metal2 s 36174 63200 36230 64000 0 FreeSans 224 90 0 0 dso_as5401[4]
port 167 nsew signal input
flabel metal2 s 36910 63200 36966 64000 0 FreeSans 224 90 0 0 dso_as5401[5]
port 168 nsew signal input
flabel metal2 s 37646 63200 37702 64000 0 FreeSans 224 90 0 0 dso_as5401[6]
port 169 nsew signal input
flabel metal2 s 38382 63200 38438 64000 0 FreeSans 224 90 0 0 dso_as5401[7]
port 170 nsew signal input
flabel metal2 s 39118 63200 39174 64000 0 FreeSans 224 90 0 0 dso_as5401[8]
port 171 nsew signal input
flabel metal2 s 39854 63200 39910 64000 0 FreeSans 224 90 0 0 dso_as5401[9]
port 172 nsew signal input
flabel metal3 s 59200 56584 60000 56704 0 FreeSans 480 0 0 0 dso_counter[0]
port 173 nsew signal input
flabel metal3 s 59200 62024 60000 62144 0 FreeSans 480 0 0 0 dso_counter[10]
port 174 nsew signal input
flabel metal3 s 59200 62568 60000 62688 0 FreeSans 480 0 0 0 dso_counter[11]
port 175 nsew signal input
flabel metal3 s 59200 57128 60000 57248 0 FreeSans 480 0 0 0 dso_counter[1]
port 176 nsew signal input
flabel metal3 s 59200 57672 60000 57792 0 FreeSans 480 0 0 0 dso_counter[2]
port 177 nsew signal input
flabel metal3 s 59200 58216 60000 58336 0 FreeSans 480 0 0 0 dso_counter[3]
port 178 nsew signal input
flabel metal3 s 59200 58760 60000 58880 0 FreeSans 480 0 0 0 dso_counter[4]
port 179 nsew signal input
flabel metal3 s 59200 59304 60000 59424 0 FreeSans 480 0 0 0 dso_counter[5]
port 180 nsew signal input
flabel metal3 s 59200 59848 60000 59968 0 FreeSans 480 0 0 0 dso_counter[6]
port 181 nsew signal input
flabel metal3 s 59200 60392 60000 60512 0 FreeSans 480 0 0 0 dso_counter[7]
port 182 nsew signal input
flabel metal3 s 59200 60936 60000 61056 0 FreeSans 480 0 0 0 dso_counter[8]
port 183 nsew signal input
flabel metal3 s 59200 61480 60000 61600 0 FreeSans 480 0 0 0 dso_counter[9]
port 184 nsew signal input
flabel metal2 s 6734 63200 6790 64000 0 FreeSans 224 90 0 0 dso_diceroll[0]
port 185 nsew signal input
flabel metal2 s 7470 63200 7526 64000 0 FreeSans 224 90 0 0 dso_diceroll[1]
port 186 nsew signal input
flabel metal2 s 8206 63200 8262 64000 0 FreeSans 224 90 0 0 dso_diceroll[2]
port 187 nsew signal input
flabel metal2 s 8942 63200 8998 64000 0 FreeSans 224 90 0 0 dso_diceroll[3]
port 188 nsew signal input
flabel metal2 s 9678 63200 9734 64000 0 FreeSans 224 90 0 0 dso_diceroll[4]
port 189 nsew signal input
flabel metal2 s 10414 63200 10470 64000 0 FreeSans 224 90 0 0 dso_diceroll[5]
port 190 nsew signal input
flabel metal2 s 11150 63200 11206 64000 0 FreeSans 224 90 0 0 dso_diceroll[6]
port 191 nsew signal input
flabel metal2 s 11886 63200 11942 64000 0 FreeSans 224 90 0 0 dso_diceroll[7]
port 192 nsew signal input
flabel metal3 s 0 30472 800 30592 0 FreeSans 480 0 0 0 dso_mc14500[0]
port 193 nsew signal input
flabel metal3 s 0 31152 800 31272 0 FreeSans 480 0 0 0 dso_mc14500[1]
port 194 nsew signal input
flabel metal3 s 0 31832 800 31952 0 FreeSans 480 0 0 0 dso_mc14500[2]
port 195 nsew signal input
flabel metal3 s 0 32512 800 32632 0 FreeSans 480 0 0 0 dso_mc14500[3]
port 196 nsew signal input
flabel metal3 s 0 33192 800 33312 0 FreeSans 480 0 0 0 dso_mc14500[4]
port 197 nsew signal input
flabel metal3 s 0 33872 800 33992 0 FreeSans 480 0 0 0 dso_mc14500[5]
port 198 nsew signal input
flabel metal3 s 0 34552 800 34672 0 FreeSans 480 0 0 0 dso_mc14500[6]
port 199 nsew signal input
flabel metal3 s 0 35232 800 35352 0 FreeSans 480 0 0 0 dso_mc14500[7]
port 200 nsew signal input
flabel metal3 s 0 35912 800 36032 0 FreeSans 480 0 0 0 dso_mc14500[8]
port 201 nsew signal input
flabel metal2 s 846 63200 902 64000 0 FreeSans 224 90 0 0 dso_multiplier[0]
port 202 nsew signal input
flabel metal2 s 1582 63200 1638 64000 0 FreeSans 224 90 0 0 dso_multiplier[1]
port 203 nsew signal input
flabel metal2 s 2318 63200 2374 64000 0 FreeSans 224 90 0 0 dso_multiplier[2]
port 204 nsew signal input
flabel metal2 s 3054 63200 3110 64000 0 FreeSans 224 90 0 0 dso_multiplier[3]
port 205 nsew signal input
flabel metal2 s 3790 63200 3846 64000 0 FreeSans 224 90 0 0 dso_multiplier[4]
port 206 nsew signal input
flabel metal2 s 4526 63200 4582 64000 0 FreeSans 224 90 0 0 dso_multiplier[5]
port 207 nsew signal input
flabel metal2 s 5262 63200 5318 64000 0 FreeSans 224 90 0 0 dso_multiplier[6]
port 208 nsew signal input
flabel metal2 s 5998 63200 6054 64000 0 FreeSans 224 90 0 0 dso_multiplier[7]
port 209 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 dso_posit[0]
port 210 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 dso_posit[1]
port 211 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 dso_posit[2]
port 212 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 dso_posit[3]
port 213 nsew signal input
flabel metal3 s 0 37272 800 37392 0 FreeSans 480 0 0 0 dso_tbb1143[0]
port 214 nsew signal input
flabel metal3 s 0 37952 800 38072 0 FreeSans 480 0 0 0 dso_tbb1143[1]
port 215 nsew signal input
flabel metal3 s 0 38632 800 38752 0 FreeSans 480 0 0 0 dso_tbb1143[2]
port 216 nsew signal input
flabel metal3 s 0 39312 800 39432 0 FreeSans 480 0 0 0 dso_tbb1143[3]
port 217 nsew signal input
flabel metal3 s 0 39992 800 40112 0 FreeSans 480 0 0 0 dso_tbb1143[4]
port 218 nsew signal input
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 dso_tbb1143[5]
port 219 nsew signal input
flabel metal3 s 0 41352 800 41472 0 FreeSans 480 0 0 0 dso_tbb1143[6]
port 220 nsew signal input
flabel metal3 s 0 42032 800 42152 0 FreeSans 480 0 0 0 dso_tbb1143[7]
port 221 nsew signal input
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 dso_tune
port 222 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 dso_vgatest[0]
port 223 nsew signal input
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 dso_vgatest[1]
port 224 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 dso_vgatest[2]
port 225 nsew signal input
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 dso_vgatest[3]
port 226 nsew signal input
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 dso_vgatest[4]
port 227 nsew signal input
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 dso_vgatest[5]
port 228 nsew signal input
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 dso_vgatest[6]
port 229 nsew signal input
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 dso_vgatest[7]
port 230 nsew signal input
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 dso_vgatest[8]
port 231 nsew signal input
flabel metal2 s 55310 0 55366 800 0 FreeSans 224 90 0 0 dso_vgatest[9]
port 232 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 io_in[0]
port 233 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 io_in[10]
port 234 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 io_in[11]
port 235 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 io_in[12]
port 236 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 io_in[13]
port 237 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 io_in[14]
port 238 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 io_in[15]
port 239 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 io_in[16]
port 240 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 io_in[17]
port 241 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 io_in[18]
port 242 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 io_in[19]
port 243 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 io_in[1]
port 244 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 io_in[20]
port 245 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 io_in[21]
port 246 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 io_in[22]
port 247 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 io_in[23]
port 248 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 io_in[24]
port 249 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 io_in[25]
port 250 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 io_in[26]
port 251 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 io_in[27]
port 252 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 io_in[28]
port 253 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 io_in[29]
port 254 nsew signal input
flabel metal2 s 5078 0 5134 800 0 FreeSans 224 90 0 0 io_in[2]
port 255 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 io_in[30]
port 256 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 io_in[31]
port 257 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 io_in[32]
port 258 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 io_in[33]
port 259 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 io_in[34]
port 260 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 io_in[35]
port 261 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 io_in[36]
port 262 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 io_in[37]
port 263 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 io_in[3]
port 264 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 io_in[4]
port 265 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 io_in[5]
port 266 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 io_in[6]
port 267 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 io_in[7]
port 268 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 io_in[8]
port 269 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 io_in[9]
port 270 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 271 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 272 nsew signal tristate
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 273 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 274 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 275 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 276 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 277 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 278 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 279 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 280 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 281 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 282 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 283 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 284 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 285 nsew signal tristate
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 286 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 287 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 288 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 289 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 290 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 291 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 292 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 293 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 294 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 295 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 296 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 297 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 298 nsew signal tristate
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 299 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 300 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 301 nsew signal tristate
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 302 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 303 nsew signal tristate
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 304 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 305 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 306 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 307 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 308 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 io_out[0]
port 309 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 io_out[10]
port 310 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 io_out[11]
port 311 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 io_out[12]
port 312 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 io_out[13]
port 313 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 io_out[14]
port 314 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 io_out[15]
port 315 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 io_out[16]
port 316 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 io_out[17]
port 317 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 io_out[18]
port 318 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 io_out[19]
port 319 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 io_out[1]
port 320 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 io_out[20]
port 321 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 io_out[21]
port 322 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 io_out[22]
port 323 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 io_out[23]
port 324 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 io_out[24]
port 325 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 io_out[25]
port 326 nsew signal tristate
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 io_out[26]
port 327 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 io_out[27]
port 328 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 io_out[28]
port 329 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 io_out[29]
port 330 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 io_out[2]
port 331 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 io_out[30]
port 332 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 io_out[31]
port 333 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 io_out[32]
port 334 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 io_out[33]
port 335 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 io_out[34]
port 336 nsew signal tristate
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 io_out[35]
port 337 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 io_out[36]
port 338 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 io_out[37]
port 339 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 io_out[3]
port 340 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 io_out[4]
port 341 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 io_out[5]
port 342 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 io_out[6]
port 343 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 io_out[7]
port 344 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 io_out[8]
port 345 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 io_out[9]
port 346 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 oeb_6502
port 347 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 oeb_as1802
port 348 nsew signal input
flabel metal2 s 12622 63200 12678 64000 0 FreeSans 224 90 0 0 oeb_as2650
port 349 nsew signal input
flabel metal3 s 0 61752 800 61872 0 FreeSans 480 0 0 0 oeb_as512512512
port 350 nsew signal input
flabel metal2 s 53102 63200 53158 64000 0 FreeSans 224 90 0 0 oeb_as5401
port 351 nsew signal input
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 oeb_mc14500
port 352 nsew signal input
flabel metal3 s 0 21632 800 21752 0 FreeSans 480 0 0 0 rst_6502
port 353 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 rst_LCD
port 354 nsew signal tristate
flabel metal3 s 0 22992 800 23112 0 FreeSans 480 0 0 0 rst_as1802
port 355 nsew signal tristate
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 rst_as2650
port 356 nsew signal tristate
flabel metal3 s 0 25032 800 25152 0 FreeSans 480 0 0 0 rst_as512512512
port 357 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 rst_as5401
port 358 nsew signal tristate
flabel metal3 s 0 25712 800 25832 0 FreeSans 480 0 0 0 rst_counter
port 359 nsew signal tristate
flabel metal3 s 0 26392 800 26512 0 FreeSans 480 0 0 0 rst_diceroll
port 360 nsew signal tristate
flabel metal3 s 0 27072 800 27192 0 FreeSans 480 0 0 0 rst_mc14500
port 361 nsew signal tristate
flabel metal3 s 0 27752 800 27872 0 FreeSans 480 0 0 0 rst_posit
port 362 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 rst_tbb1143
port 363 nsew signal tristate
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 rst_tune
port 364 nsew signal tristate
flabel metal3 s 0 29792 800 29912 0 FreeSans 480 0 0 0 rst_vgatest
port 365 nsew signal tristate
flabel metal4 s 4208 2128 4528 61520 0 FreeSans 1920 90 0 0 vccd1
port 366 nsew power bidirectional
flabel metal4 s 34928 2128 35248 61520 0 FreeSans 1920 90 0 0 vccd1
port 366 nsew power bidirectional
flabel metal4 s 19568 2128 19888 61520 0 FreeSans 1920 90 0 0 vssd1
port 367 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 61520 0 FreeSans 1920 90 0 0 vssd1
port 367 nsew ground bidirectional
flabel metal3 s 59200 1096 60000 1216 0 FreeSans 480 0 0 0 wb_clk_i
port 368 nsew signal input
flabel metal3 s 59200 1640 60000 1760 0 FreeSans 480 0 0 0 wb_rst_i
port 369 nsew signal input
flabel metal3 s 59200 2184 60000 2304 0 FreeSans 480 0 0 0 wbs_ack_o
port 370 nsew signal tristate
flabel metal3 s 59200 4360 60000 4480 0 FreeSans 480 0 0 0 wbs_adr_i[0]
port 371 nsew signal input
flabel metal3 s 59200 20680 60000 20800 0 FreeSans 480 0 0 0 wbs_adr_i[10]
port 372 nsew signal input
flabel metal3 s 59200 22312 60000 22432 0 FreeSans 480 0 0 0 wbs_adr_i[11]
port 373 nsew signal input
flabel metal3 s 59200 23944 60000 24064 0 FreeSans 480 0 0 0 wbs_adr_i[12]
port 374 nsew signal input
flabel metal3 s 59200 25576 60000 25696 0 FreeSans 480 0 0 0 wbs_adr_i[13]
port 375 nsew signal input
flabel metal3 s 59200 27208 60000 27328 0 FreeSans 480 0 0 0 wbs_adr_i[14]
port 376 nsew signal input
flabel metal3 s 59200 28840 60000 28960 0 FreeSans 480 0 0 0 wbs_adr_i[15]
port 377 nsew signal input
flabel metal3 s 59200 30472 60000 30592 0 FreeSans 480 0 0 0 wbs_adr_i[16]
port 378 nsew signal input
flabel metal3 s 59200 32104 60000 32224 0 FreeSans 480 0 0 0 wbs_adr_i[17]
port 379 nsew signal input
flabel metal3 s 59200 33736 60000 33856 0 FreeSans 480 0 0 0 wbs_adr_i[18]
port 380 nsew signal input
flabel metal3 s 59200 35368 60000 35488 0 FreeSans 480 0 0 0 wbs_adr_i[19]
port 381 nsew signal input
flabel metal3 s 59200 5992 60000 6112 0 FreeSans 480 0 0 0 wbs_adr_i[1]
port 382 nsew signal input
flabel metal3 s 59200 37000 60000 37120 0 FreeSans 480 0 0 0 wbs_adr_i[20]
port 383 nsew signal input
flabel metal3 s 59200 38632 60000 38752 0 FreeSans 480 0 0 0 wbs_adr_i[21]
port 384 nsew signal input
flabel metal3 s 59200 40264 60000 40384 0 FreeSans 480 0 0 0 wbs_adr_i[22]
port 385 nsew signal input
flabel metal3 s 59200 41896 60000 42016 0 FreeSans 480 0 0 0 wbs_adr_i[23]
port 386 nsew signal input
flabel metal3 s 59200 43528 60000 43648 0 FreeSans 480 0 0 0 wbs_adr_i[24]
port 387 nsew signal input
flabel metal3 s 59200 45160 60000 45280 0 FreeSans 480 0 0 0 wbs_adr_i[25]
port 388 nsew signal input
flabel metal3 s 59200 46792 60000 46912 0 FreeSans 480 0 0 0 wbs_adr_i[26]
port 389 nsew signal input
flabel metal3 s 59200 48424 60000 48544 0 FreeSans 480 0 0 0 wbs_adr_i[27]
port 390 nsew signal input
flabel metal3 s 59200 50056 60000 50176 0 FreeSans 480 0 0 0 wbs_adr_i[28]
port 391 nsew signal input
flabel metal3 s 59200 51688 60000 51808 0 FreeSans 480 0 0 0 wbs_adr_i[29]
port 392 nsew signal input
flabel metal3 s 59200 7624 60000 7744 0 FreeSans 480 0 0 0 wbs_adr_i[2]
port 393 nsew signal input
flabel metal3 s 59200 53320 60000 53440 0 FreeSans 480 0 0 0 wbs_adr_i[30]
port 394 nsew signal input
flabel metal3 s 59200 54952 60000 55072 0 FreeSans 480 0 0 0 wbs_adr_i[31]
port 395 nsew signal input
flabel metal3 s 59200 9256 60000 9376 0 FreeSans 480 0 0 0 wbs_adr_i[3]
port 396 nsew signal input
flabel metal3 s 59200 10888 60000 11008 0 FreeSans 480 0 0 0 wbs_adr_i[4]
port 397 nsew signal input
flabel metal3 s 59200 12520 60000 12640 0 FreeSans 480 0 0 0 wbs_adr_i[5]
port 398 nsew signal input
flabel metal3 s 59200 14152 60000 14272 0 FreeSans 480 0 0 0 wbs_adr_i[6]
port 399 nsew signal input
flabel metal3 s 59200 15784 60000 15904 0 FreeSans 480 0 0 0 wbs_adr_i[7]
port 400 nsew signal input
flabel metal3 s 59200 17416 60000 17536 0 FreeSans 480 0 0 0 wbs_adr_i[8]
port 401 nsew signal input
flabel metal3 s 59200 19048 60000 19168 0 FreeSans 480 0 0 0 wbs_adr_i[9]
port 402 nsew signal input
flabel metal3 s 59200 2728 60000 2848 0 FreeSans 480 0 0 0 wbs_cyc_i
port 403 nsew signal input
flabel metal3 s 59200 4904 60000 5024 0 FreeSans 480 0 0 0 wbs_dat_i[0]
port 404 nsew signal input
flabel metal3 s 59200 21224 60000 21344 0 FreeSans 480 0 0 0 wbs_dat_i[10]
port 405 nsew signal input
flabel metal3 s 59200 22856 60000 22976 0 FreeSans 480 0 0 0 wbs_dat_i[11]
port 406 nsew signal input
flabel metal3 s 59200 24488 60000 24608 0 FreeSans 480 0 0 0 wbs_dat_i[12]
port 407 nsew signal input
flabel metal3 s 59200 26120 60000 26240 0 FreeSans 480 0 0 0 wbs_dat_i[13]
port 408 nsew signal input
flabel metal3 s 59200 27752 60000 27872 0 FreeSans 480 0 0 0 wbs_dat_i[14]
port 409 nsew signal input
flabel metal3 s 59200 29384 60000 29504 0 FreeSans 480 0 0 0 wbs_dat_i[15]
port 410 nsew signal input
flabel metal3 s 59200 31016 60000 31136 0 FreeSans 480 0 0 0 wbs_dat_i[16]
port 411 nsew signal input
flabel metal3 s 59200 32648 60000 32768 0 FreeSans 480 0 0 0 wbs_dat_i[17]
port 412 nsew signal input
flabel metal3 s 59200 34280 60000 34400 0 FreeSans 480 0 0 0 wbs_dat_i[18]
port 413 nsew signal input
flabel metal3 s 59200 35912 60000 36032 0 FreeSans 480 0 0 0 wbs_dat_i[19]
port 414 nsew signal input
flabel metal3 s 59200 6536 60000 6656 0 FreeSans 480 0 0 0 wbs_dat_i[1]
port 415 nsew signal input
flabel metal3 s 59200 37544 60000 37664 0 FreeSans 480 0 0 0 wbs_dat_i[20]
port 416 nsew signal input
flabel metal3 s 59200 39176 60000 39296 0 FreeSans 480 0 0 0 wbs_dat_i[21]
port 417 nsew signal input
flabel metal3 s 59200 40808 60000 40928 0 FreeSans 480 0 0 0 wbs_dat_i[22]
port 418 nsew signal input
flabel metal3 s 59200 42440 60000 42560 0 FreeSans 480 0 0 0 wbs_dat_i[23]
port 419 nsew signal input
flabel metal3 s 59200 44072 60000 44192 0 FreeSans 480 0 0 0 wbs_dat_i[24]
port 420 nsew signal input
flabel metal3 s 59200 45704 60000 45824 0 FreeSans 480 0 0 0 wbs_dat_i[25]
port 421 nsew signal input
flabel metal3 s 59200 47336 60000 47456 0 FreeSans 480 0 0 0 wbs_dat_i[26]
port 422 nsew signal input
flabel metal3 s 59200 48968 60000 49088 0 FreeSans 480 0 0 0 wbs_dat_i[27]
port 423 nsew signal input
flabel metal3 s 59200 50600 60000 50720 0 FreeSans 480 0 0 0 wbs_dat_i[28]
port 424 nsew signal input
flabel metal3 s 59200 52232 60000 52352 0 FreeSans 480 0 0 0 wbs_dat_i[29]
port 425 nsew signal input
flabel metal3 s 59200 8168 60000 8288 0 FreeSans 480 0 0 0 wbs_dat_i[2]
port 426 nsew signal input
flabel metal3 s 59200 53864 60000 53984 0 FreeSans 480 0 0 0 wbs_dat_i[30]
port 427 nsew signal input
flabel metal3 s 59200 55496 60000 55616 0 FreeSans 480 0 0 0 wbs_dat_i[31]
port 428 nsew signal input
flabel metal3 s 59200 9800 60000 9920 0 FreeSans 480 0 0 0 wbs_dat_i[3]
port 429 nsew signal input
flabel metal3 s 59200 11432 60000 11552 0 FreeSans 480 0 0 0 wbs_dat_i[4]
port 430 nsew signal input
flabel metal3 s 59200 13064 60000 13184 0 FreeSans 480 0 0 0 wbs_dat_i[5]
port 431 nsew signal input
flabel metal3 s 59200 14696 60000 14816 0 FreeSans 480 0 0 0 wbs_dat_i[6]
port 432 nsew signal input
flabel metal3 s 59200 16328 60000 16448 0 FreeSans 480 0 0 0 wbs_dat_i[7]
port 433 nsew signal input
flabel metal3 s 59200 17960 60000 18080 0 FreeSans 480 0 0 0 wbs_dat_i[8]
port 434 nsew signal input
flabel metal3 s 59200 19592 60000 19712 0 FreeSans 480 0 0 0 wbs_dat_i[9]
port 435 nsew signal input
flabel metal3 s 59200 5448 60000 5568 0 FreeSans 480 0 0 0 wbs_dat_o[0]
port 436 nsew signal tristate
flabel metal3 s 59200 21768 60000 21888 0 FreeSans 480 0 0 0 wbs_dat_o[10]
port 437 nsew signal tristate
flabel metal3 s 59200 23400 60000 23520 0 FreeSans 480 0 0 0 wbs_dat_o[11]
port 438 nsew signal tristate
flabel metal3 s 59200 25032 60000 25152 0 FreeSans 480 0 0 0 wbs_dat_o[12]
port 439 nsew signal tristate
flabel metal3 s 59200 26664 60000 26784 0 FreeSans 480 0 0 0 wbs_dat_o[13]
port 440 nsew signal tristate
flabel metal3 s 59200 28296 60000 28416 0 FreeSans 480 0 0 0 wbs_dat_o[14]
port 441 nsew signal tristate
flabel metal3 s 59200 29928 60000 30048 0 FreeSans 480 0 0 0 wbs_dat_o[15]
port 442 nsew signal tristate
flabel metal3 s 59200 31560 60000 31680 0 FreeSans 480 0 0 0 wbs_dat_o[16]
port 443 nsew signal tristate
flabel metal3 s 59200 33192 60000 33312 0 FreeSans 480 0 0 0 wbs_dat_o[17]
port 444 nsew signal tristate
flabel metal3 s 59200 34824 60000 34944 0 FreeSans 480 0 0 0 wbs_dat_o[18]
port 445 nsew signal tristate
flabel metal3 s 59200 36456 60000 36576 0 FreeSans 480 0 0 0 wbs_dat_o[19]
port 446 nsew signal tristate
flabel metal3 s 59200 7080 60000 7200 0 FreeSans 480 0 0 0 wbs_dat_o[1]
port 447 nsew signal tristate
flabel metal3 s 59200 38088 60000 38208 0 FreeSans 480 0 0 0 wbs_dat_o[20]
port 448 nsew signal tristate
flabel metal3 s 59200 39720 60000 39840 0 FreeSans 480 0 0 0 wbs_dat_o[21]
port 449 nsew signal tristate
flabel metal3 s 59200 41352 60000 41472 0 FreeSans 480 0 0 0 wbs_dat_o[22]
port 450 nsew signal tristate
flabel metal3 s 59200 42984 60000 43104 0 FreeSans 480 0 0 0 wbs_dat_o[23]
port 451 nsew signal tristate
flabel metal3 s 59200 44616 60000 44736 0 FreeSans 480 0 0 0 wbs_dat_o[24]
port 452 nsew signal tristate
flabel metal3 s 59200 46248 60000 46368 0 FreeSans 480 0 0 0 wbs_dat_o[25]
port 453 nsew signal tristate
flabel metal3 s 59200 47880 60000 48000 0 FreeSans 480 0 0 0 wbs_dat_o[26]
port 454 nsew signal tristate
flabel metal3 s 59200 49512 60000 49632 0 FreeSans 480 0 0 0 wbs_dat_o[27]
port 455 nsew signal tristate
flabel metal3 s 59200 51144 60000 51264 0 FreeSans 480 0 0 0 wbs_dat_o[28]
port 456 nsew signal tristate
flabel metal3 s 59200 52776 60000 52896 0 FreeSans 480 0 0 0 wbs_dat_o[29]
port 457 nsew signal tristate
flabel metal3 s 59200 8712 60000 8832 0 FreeSans 480 0 0 0 wbs_dat_o[2]
port 458 nsew signal tristate
flabel metal3 s 59200 54408 60000 54528 0 FreeSans 480 0 0 0 wbs_dat_o[30]
port 459 nsew signal tristate
flabel metal3 s 59200 56040 60000 56160 0 FreeSans 480 0 0 0 wbs_dat_o[31]
port 460 nsew signal tristate
flabel metal3 s 59200 10344 60000 10464 0 FreeSans 480 0 0 0 wbs_dat_o[3]
port 461 nsew signal tristate
flabel metal3 s 59200 11976 60000 12096 0 FreeSans 480 0 0 0 wbs_dat_o[4]
port 462 nsew signal tristate
flabel metal3 s 59200 13608 60000 13728 0 FreeSans 480 0 0 0 wbs_dat_o[5]
port 463 nsew signal tristate
flabel metal3 s 59200 15240 60000 15360 0 FreeSans 480 0 0 0 wbs_dat_o[6]
port 464 nsew signal tristate
flabel metal3 s 59200 16872 60000 16992 0 FreeSans 480 0 0 0 wbs_dat_o[7]
port 465 nsew signal tristate
flabel metal3 s 59200 18504 60000 18624 0 FreeSans 480 0 0 0 wbs_dat_o[8]
port 466 nsew signal tristate
flabel metal3 s 59200 20136 60000 20256 0 FreeSans 480 0 0 0 wbs_dat_o[9]
port 467 nsew signal tristate
flabel metal3 s 59200 3272 60000 3392 0 FreeSans 480 0 0 0 wbs_stb_i
port 468 nsew signal input
flabel metal3 s 59200 3816 60000 3936 0 FreeSans 480 0 0 0 wbs_we_i
port 469 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 64000
<< end >>
