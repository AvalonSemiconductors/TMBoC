// This is the unpowered netlist.
module tholin_avalonsemi_5401 (clk,
    io_oeb,
    rst,
    io_in,
    io_out);
 input clk;
 output io_oeb;
 input rst;
 input [9:0] io_in;
 output [26:0] io_out;

 wire \CIRCUIT_1957.D0 ;
 wire \CIRCUIT_1957.D1 ;
 wire \CIRCUIT_1957.D2 ;
 wire \CIRCUIT_1957.D3 ;
 wire \CIRCUIT_1957.GATES_10.result ;
 wire \CIRCUIT_1957.GATES_27.result ;
 wire \CIRCUIT_1957.GATES_28.result ;
 wire \CIRCUIT_1957.GATES_30.result ;
 wire \CIRCUIT_1957.GATES_33.input2 ;
 wire \CIRCUIT_1957.GATES_35.result ;
 wire \CIRCUIT_1957.GATES_38.result ;
 wire \CIRCUIT_1957.GATES_39.result ;
 wire \CIRCUIT_1957.GATES_40.result ;
 wire \CIRCUIT_1957.GATES_41.result ;
 wire \CIRCUIT_1957.GATES_42.result ;
 wire \CIRCUIT_1957.GATES_53.result ;
 wire \CIRCUIT_1957.GATES_60.result ;
 wire \CIRCUIT_1957.GATES_9.result ;
 wire \CIRCUIT_1957.MEMORY_62.d ;
 wire \CIRCUIT_1957.MEMORY_62.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_63.d ;
 wire \CIRCUIT_1957.MEMORY_63.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_64.d ;
 wire \CIRCUIT_1957.MEMORY_64.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_65.d ;
 wire \CIRCUIT_1957.MEMORY_65.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_66.d ;
 wire \CIRCUIT_1957.MEMORY_66.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_67.d ;
 wire \CIRCUIT_1957.MEMORY_67.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_68.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_69.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_70.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_71.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_72.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_73.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_74.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_75.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_76.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_77.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_78.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_79.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_80.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_81.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_82.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_83.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_84.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_85.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_86.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_87.s_currentState ;
 wire \CIRCUIT_1957.MEMORY_88.s_currentState ;
 wire \CIRCUIT_1957.clock_gen_2_1.CLK1 ;
 wire \CIRCUIT_1957.clock_gen_2_1.GATES_1.input2 ;
 wire \CIRCUIT_1957.clock_gen_2_1.GATES_3.result ;
 wire \CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ;
 wire \CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ;
 wire \CIRCUIT_1957.clock_gen_2_1.MEMORY_5.d ;
 wire \CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ;
 wire \CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ;
 wire \CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1 ;
 wire \CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ;
 wire \CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result ;
 wire \CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState ;
 wire \CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ;
 wire \CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ;
 wire \CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ;
 wire \CIRCUIT_1957.int_memory_1.GATES_1.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_1.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_1.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_1.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_2.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_2.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_2.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_2.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_21.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_22.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_23.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_24.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_25.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_26.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_27.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_28.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_29.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_3.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_3.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_3.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_3.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_30.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_31.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_32.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_33.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_4.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_4.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_4.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_4.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_49.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_49.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_49.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_49.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_5.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_5.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_5.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_5.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_50.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_51.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_51.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_51.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_51.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_53.result ;
 wire \CIRCUIT_1957.int_memory_1.GATES_6.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_6.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_6.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_6.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_7.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_7.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_7.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_7.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_8.input2[0] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_8.input2[1] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_8.input2[2] ;
 wire \CIRCUIT_1957.int_memory_1.GATES_8.input2[3] ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A0 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A1 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A2 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A3 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A4 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A5 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A6 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.A7 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.B0 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.B1 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.B2 ;
 wire \CIRCUIT_1957.int_memory_1.div_1.B3 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.A0 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.A1 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.A2 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.A3 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.B0 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.B1 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.B2 ;
 wire \CIRCUIT_1957.int_memory_1.mul2_1.B3 ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire clknet_0_clk;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire net39;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net40;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ;
 wire clknet_0__0498_;
 wire clknet_1_0__leaf__0498_;
 wire clknet_1_1__leaf__0498_;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ;
 wire clknet_0__0142_;
 wire clknet_1_0__leaf__0142_;
 wire clknet_1_1__leaf__0142_;
 wire clknet_0__0526_;
 wire clknet_1_0__leaf__0526_;
 wire clknet_1_1__leaf__0526_;
 wire clknet_0__0502_;
 wire clknet_1_0__leaf__0502_;
 wire clknet_1_1__leaf__0502_;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ;
 wire \clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result ;
 wire \clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ;
 wire \clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ;
 wire clknet_0__0143_;
 wire clknet_1_0__leaf__0143_;
 wire clknet_1_1__leaf__0143_;

 sky130_fd_sc_hd__clkinv_2 _0534_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState ),
    .Y(_0099_));
 sky130_fd_sc_hd__nor2_1 _0535_ (.A(_0099_),
    .B(\CIRCUIT_1957.MEMORY_64.s_currentState ),
    .Y(_0100_));
 sky130_fd_sc_hd__or4_1 _0536_ (.A(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_65.s_currentState ),
    .C(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .D(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .X(_0101_));
 sky130_fd_sc_hd__buf_2 _0537_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState ),
    .X(_0102_));
 sky130_fd_sc_hd__o22a_1 _0538_ (.A1(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .A2(_0100_),
    .B1(_0101_),
    .B2(_0102_),
    .X(_0103_));
 sky130_fd_sc_hd__nor3b_4 _0539_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .B(_0103_),
    .C_N(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .Y(_0104_));
 sky130_fd_sc_hd__mux2_1 _0540_ (.A0(\CIRCUIT_1957.MEMORY_75.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_83.s_currentState ),
    .S(_0104_),
    .X(_0105_));
 sky130_fd_sc_hd__clkinv_2 _0541_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ),
    .Y(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ));
 sky130_fd_sc_hd__mux2_1 _0542_ (.A0(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .A1(_0105_),
    .S(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .X(_0106_));
 sky130_fd_sc_hd__or4b_1 _0543_ (.A(net22),
    .B(net21),
    .C(net25),
    .D_N(net24),
    .X(_0107_));
 sky130_fd_sc_hd__buf_2 _0544_ (.A(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _0545_ (.A0(_0106_),
    .A1(net20),
    .S(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__clkbuf_1 _0546_ (.A(_0109_),
    .X(_0060_));
 sky130_fd_sc_hd__or3b_1 _0547_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ),
    .B(_0104_),
    .C_N(\CIRCUIT_1957.MEMORY_74.s_currentState ),
    .X(_0110_));
 sky130_fd_sc_hd__o21ai_1 _0548_ (.A1(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_82.s_currentState ),
    .B1(_0104_),
    .Y(_0111_));
 sky130_fd_sc_hd__a21oi_1 _0549_ (.A1(_0110_),
    .A2(_0111_),
    .B1(_0108_),
    .Y(_0112_));
 sky130_fd_sc_hd__a21o_1 _0550_ (.A1(net19),
    .A2(_0108_),
    .B1(_0112_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0551_ (.A0(\CIRCUIT_1957.MEMORY_73.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_81.s_currentState ),
    .S(_0104_),
    .X(_0113_));
 sky130_fd_sc_hd__nand2_1 _0552_ (.A(\CIRCUIT_1957.MEMORY_75.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_74.s_currentState ),
    .Y(_0114_));
 sky130_fd_sc_hd__or4bb_4 _0553_ (.A(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .B(_0114_),
    .C_N(\CIRCUIT_1957.MEMORY_72.s_currentState ),
    .D_N(\CIRCUIT_1957.MEMORY_73.s_currentState ),
    .X(_0115_));
 sky130_fd_sc_hd__nand2_1 _0554_ (.A(\CIRCUIT_1957.MEMORY_70.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_71.s_currentState ),
    .Y(_0116_));
 sky130_fd_sc_hd__nand2_2 _0555_ (.A(\CIRCUIT_1957.MEMORY_68.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_69.s_currentState ),
    .Y(_0117_));
 sky130_fd_sc_hd__nor2_1 _0556_ (.A(_0116_),
    .B(_0117_),
    .Y(_0118_));
 sky130_fd_sc_hd__nor2_4 _0557_ (.A(_0115_),
    .B(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__nor2_1 _0558_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .B(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .Y(_0120_));
 sky130_fd_sc_hd__or3b_1 _0559_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .B(_0099_),
    .C_N(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__nor2_1 _0560_ (.A(_0119_),
    .B(_0121_),
    .Y(_0122_));
 sky130_fd_sc_hd__mux2_1 _0561_ (.A0(_0113_),
    .A1(_0122_),
    .S(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _0562_ (.A0(_0123_),
    .A1(net18),
    .S(_0108_),
    .X(_0124_));
 sky130_fd_sc_hd__clkbuf_1 _0563_ (.A(_0124_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0564_ (.A0(\CIRCUIT_1957.MEMORY_72.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_80.s_currentState ),
    .S(_0104_),
    .X(_0125_));
 sky130_fd_sc_hd__nand2_1 _0565_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .B(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _0566_ (.A(_0126_),
    .Y(_0127_));
 sky130_fd_sc_hd__and2_1 _0567_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .B(_0102_),
    .X(_0128_));
 sky130_fd_sc_hd__o21a_1 _0568_ (.A1(_0120_),
    .A2(_0127_),
    .B1(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _0569_ (.A0(_0125_),
    .A1(_0129_),
    .S(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _0570_ (.A0(_0130_),
    .A1(net17),
    .S(_0108_),
    .X(_0131_));
 sky130_fd_sc_hd__clkbuf_1 _0571_ (.A(_0131_),
    .X(_0057_));
 sky130_fd_sc_hd__mux4_1 _0572_ (.A0(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_71.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_87.s_currentState ),
    .A3(\CIRCUIT_1957.MEMORY_79.s_currentState ),
    .S0(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .S1(_0104_),
    .X(_0132_));
 sky130_fd_sc_hd__clkbuf_1 _0573_ (.A(_0132_),
    .X(net27));
 sky130_fd_sc_hd__mux2_1 _0574_ (.A0(net27),
    .A1(net16),
    .S(_0108_),
    .X(_0133_));
 sky130_fd_sc_hd__clkbuf_1 _0575_ (.A(_0133_),
    .X(_0056_));
 sky130_fd_sc_hd__mux4_1 _0576_ (.A0(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_70.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_86.s_currentState ),
    .A3(\CIRCUIT_1957.MEMORY_78.s_currentState ),
    .S0(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .S1(_0104_),
    .X(_0134_));
 sky130_fd_sc_hd__clkbuf_1 _0577_ (.A(_0134_),
    .X(net26));
 sky130_fd_sc_hd__mux2_1 _0578_ (.A0(net26),
    .A1(net15),
    .S(_0108_),
    .X(_0135_));
 sky130_fd_sc_hd__clkbuf_1 _0579_ (.A(_0135_),
    .X(_0055_));
 sky130_fd_sc_hd__mux4_1 _0580_ (.A0(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_69.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_85.s_currentState ),
    .A3(\CIRCUIT_1957.MEMORY_77.s_currentState ),
    .S0(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .S1(_0104_),
    .X(_0136_));
 sky130_fd_sc_hd__clkbuf_1 _0581_ (.A(_0136_),
    .X(net23));
 sky130_fd_sc_hd__mux2_1 _0582_ (.A0(net23),
    .A1(net14),
    .S(_0108_),
    .X(_0137_));
 sky130_fd_sc_hd__clkbuf_1 _0583_ (.A(_0137_),
    .X(_0054_));
 sky130_fd_sc_hd__mux4_1 _0584_ (.A0(\CIRCUIT_1957.MEMORY_65.s_currentState ),
    .A1(\CIRCUIT_1957.MEMORY_68.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_84.s_currentState ),
    .A3(\CIRCUIT_1957.MEMORY_76.s_currentState ),
    .S0(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .S1(_0104_),
    .X(_0138_));
 sky130_fd_sc_hd__clkbuf_1 _0585_ (.A(_0138_),
    .X(net12));
 sky130_fd_sc_hd__mux2_1 _0586_ (.A0(net12),
    .A1(net13),
    .S(_0108_),
    .X(_0139_));
 sky130_fd_sc_hd__clkbuf_1 _0587_ (.A(_0139_),
    .X(_0053_));
 sky130_fd_sc_hd__clkbuf_4 _0588_ (.A(net11),
    .X(_0140_));
 sky130_fd_sc_hd__buf_4 _0589_ (.A(_0140_),
    .X(_0141_));
 sky130_fd_sc_hd__buf_1 _0590_ (.A(clknet_1_0__leaf_clk),
    .X(_0142_));
 sky130_fd_sc_hd__buf_1 _0591_ (.A(clknet_1_0__leaf__0142_),
    .X(_0143_));
 sky130_fd_sc_hd__nand2_2 _0592_ (.A(_0141_),
    .B(clknet_1_1__leaf__0143_),
    .Y(_0002_));
 sky130_fd_sc_hd__or4b_4 _0593_ (.A(net22),
    .B(net25),
    .C(net24),
    .D_N(net21),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _0594_ (.A0(net5),
    .A1(net1),
    .S(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__clkbuf_1 _0595_ (.A(_0145_),
    .X(\CIRCUIT_1957.D0 ));
 sky130_fd_sc_hd__mux2_1 _0596_ (.A0(net6),
    .A1(net2),
    .S(_0144_),
    .X(_0146_));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(_0146_),
    .X(\CIRCUIT_1957.D1 ));
 sky130_fd_sc_hd__mux2_1 _0598_ (.A0(net7),
    .A1(net3),
    .S(_0144_),
    .X(_0147_));
 sky130_fd_sc_hd__clkbuf_1 _0599_ (.A(_0147_),
    .X(\CIRCUIT_1957.D2 ));
 sky130_fd_sc_hd__mux2_1 _0600_ (.A0(net8),
    .A1(net4),
    .S(_0144_),
    .X(_0148_));
 sky130_fd_sc_hd__clkbuf_1 _0601_ (.A(_0148_),
    .X(\CIRCUIT_1957.D3 ));
 sky130_fd_sc_hd__inv_2 _0602_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ),
    .Y(\CIRCUIT_1957.clock_gen_2_1.GATES_1.input2 ));
 sky130_fd_sc_hd__nand2_2 _0603_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .B(\CIRCUIT_1957.clock_gen_2_1.GATES_1.input2 ),
    .Y(_0149_));
 sky130_fd_sc_hd__and3b_1 _0604_ (.A_N(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .B(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .C(_0128_),
    .X(_0150_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0605_ (.A(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__nand2_1 _0606_ (.A(_0149_),
    .B(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__a21o_1 _0607_ (.A1(\CIRCUIT_1957.GATES_33.input2 ),
    .A2(_0152_),
    .B1(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ),
    .X(_0153_));
 sky130_fd_sc_hd__inv_2 _0608_ (.A(\CIRCUIT_1957.GATES_33.input2 ),
    .Y(_0154_));
 sky130_fd_sc_hd__a31o_1 _0609_ (.A1(_0154_),
    .A2(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ),
    .A3(_0152_),
    .B1(net11),
    .X(_0155_));
 sky130_fd_sc_hd__a21o_1 _0610_ (.A1(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1 ),
    .A2(_0153_),
    .B1(_0155_),
    .X(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ));
 sky130_fd_sc_hd__inv_2 _0611_ (.A(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result ),
    .Y(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1 ));
 sky130_fd_sc_hd__inv_2 _0612_ (.A(_0149_),
    .Y(\CIRCUIT_1957.clock_gen_2_1.CLK1 ));
 sky130_fd_sc_hd__inv_2 _0613_ (.A(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ),
    .Y(_0156_));
 sky130_fd_sc_hd__mux2_1 _0614_ (.A0(_0156_),
    .A1(\CIRCUIT_1957.GATES_33.input2 ),
    .S(_0152_),
    .X(_0157_));
 sky130_fd_sc_hd__and3b_1 _0615_ (.A_N(_0140_),
    .B(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input1 ),
    .C(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__clkbuf_1 _0616_ (.A(_0158_),
    .X(\CIRCUIT_1957.GATES_33.input2 ));
 sky130_fd_sc_hd__a41o_1 _0617_ (.A1(_0154_),
    .A2(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result ),
    .A3(_0149_),
    .A4(_0151_),
    .B1(_0155_),
    .X(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_26.result ));
 sky130_fd_sc_hd__clkinv_2 _0618_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .Y(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.d ));
 sky130_fd_sc_hd__nand2_1 _0619_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .B(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ),
    .Y(_0159_));
 sky130_fd_sc_hd__nor2_1 _0620_ (.A(_0151_),
    .B(_0159_),
    .Y(\CIRCUIT_1957.GATES_53.result ));
 sky130_fd_sc_hd__or4_2 _0621_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .B(_0102_),
    .C(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .D(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .X(_0160_));
 sky130_fd_sc_hd__and2_1 _0622_ (.A(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .B(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__buf_2 _0623_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B1 ),
    .X(_0162_));
 sky130_fd_sc_hd__clkinv_2 _0624_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B0 ),
    .Y(_0163_));
 sky130_fd_sc_hd__nor2_1 _0625_ (.A(_0163_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A0 ),
    .Y(_0164_));
 sky130_fd_sc_hd__and2_1 _0626_ (.A(_0162_),
    .B(_0164_),
    .X(_0165_));
 sky130_fd_sc_hd__buf_2 _0627_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B0 ),
    .X(_0166_));
 sky130_fd_sc_hd__clkbuf_4 _0628_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B3 ),
    .X(_0167_));
 sky130_fd_sc_hd__inv_2 _0629_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B3 ),
    .Y(_0168_));
 sky130_fd_sc_hd__nor2_2 _0630_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B3 ),
    .B(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _0631_ (.A(\CIRCUIT_1957.int_memory_1.div_1.A6 ),
    .Y(_0170_));
 sky130_fd_sc_hd__a211o_1 _0632_ (.A1(_0166_),
    .A2(_0169_),
    .B1(_0170_),
    .C1(\CIRCUIT_1957.int_memory_1.div_1.B1 ),
    .X(_0171_));
 sky130_fd_sc_hd__nor2_1 _0633_ (.A(_0163_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A5 ),
    .Y(_0172_));
 sky130_fd_sc_hd__nand2_1 _0634_ (.A(_0171_),
    .B(_0172_),
    .Y(_0173_));
 sky130_fd_sc_hd__or2b_1 _0635_ (.A(\CIRCUIT_1957.int_memory_1.div_1.A7 ),
    .B_N(\CIRCUIT_1957.int_memory_1.div_1.B1 ),
    .X(_0174_));
 sky130_fd_sc_hd__a31o_1 _0636_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.B0 ),
    .A2(_0169_),
    .A3(_0174_),
    .B1(_0170_),
    .X(_0175_));
 sky130_fd_sc_hd__nand2_1 _0637_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B1 ),
    .B(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _0638_ (.A(\CIRCUIT_1957.int_memory_1.div_1.A7 ),
    .Y(_0177_));
 sky130_fd_sc_hd__nor2_1 _0639_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B0 ),
    .B(\CIRCUIT_1957.int_memory_1.div_1.B1 ),
    .Y(_0178_));
 sky130_fd_sc_hd__and3b_1 _0640_ (.A_N(\CIRCUIT_1957.int_memory_1.div_1.A6 ),
    .B(\CIRCUIT_1957.int_memory_1.div_1.B1 ),
    .C(\CIRCUIT_1957.int_memory_1.div_1.B0 ),
    .X(_0179_));
 sky130_fd_sc_hd__inv_2 _0641_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .Y(_0180_));
 sky130_fd_sc_hd__o311a_1 _0642_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.B3 ),
    .A2(_0178_),
    .A3(_0179_),
    .B1(_0180_),
    .C1(\CIRCUIT_1957.int_memory_1.div_1.A7 ),
    .X(_0181_));
 sky130_fd_sc_hd__a211oi_1 _0643_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .A2(_0177_),
    .B1(_0181_),
    .C1(\CIRCUIT_1957.int_memory_1.div_1.B3 ),
    .Y(_0182_));
 sky130_fd_sc_hd__and2b_1 _0644_ (.A_N(_0178_),
    .B(_0169_),
    .X(_0183_));
 sky130_fd_sc_hd__a311oi_2 _0645_ (.A1(_0173_),
    .A2(_0176_),
    .A3(_0182_),
    .B1(_0183_),
    .C1(_0177_),
    .Y(_0184_));
 sky130_fd_sc_hd__and2_1 _0646_ (.A(_0168_),
    .B(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__a21o_1 _0647_ (.A1(_0171_),
    .A2(_0176_),
    .B1(_0172_),
    .X(_0186_));
 sky130_fd_sc_hd__a32o_1 _0648_ (.A1(_0173_),
    .A2(_0176_),
    .A3(_0182_),
    .B1(_0181_),
    .B2(_0168_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _0649_ (.A0(_0175_),
    .A1(_0186_),
    .S(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__nor2_1 _0650_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .B(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__nor2_1 _0651_ (.A(_0163_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A4 ),
    .Y(_0190_));
 sky130_fd_sc_hd__nor2_1 _0652_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B1 ),
    .B(_0190_),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _0653_ (.A(\CIRCUIT_1957.int_memory_1.div_1.A5 ),
    .Y(_0192_));
 sky130_fd_sc_hd__and3_1 _0654_ (.A(_0166_),
    .B(_0192_),
    .C(_0187_),
    .X(_0193_));
 sky130_fd_sc_hd__a21oi_1 _0655_ (.A1(_0166_),
    .A2(_0187_),
    .B1(_0192_),
    .Y(_0194_));
 sky130_fd_sc_hd__and2_1 _0656_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B1 ),
    .B(_0190_),
    .X(_0195_));
 sky130_fd_sc_hd__o21ba_1 _0657_ (.A1(_0193_),
    .A2(_0194_),
    .B1_N(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__o2bb2a_1 _0658_ (.A1_N(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .A2_N(_0188_),
    .B1(_0191_),
    .B2(_0196_),
    .X(_0197_));
 sky130_fd_sc_hd__nand2_1 _0659_ (.A(_0167_),
    .B(_0177_),
    .Y(_0198_));
 sky130_fd_sc_hd__o311a_1 _0660_ (.A1(_0185_),
    .A2(_0189_),
    .A3(_0197_),
    .B1(_0198_),
    .C1(_0166_),
    .X(_0199_));
 sky130_fd_sc_hd__xor2_2 _0661_ (.A(\CIRCUIT_1957.int_memory_1.div_1.A4 ),
    .B(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__o31ai_2 _0662_ (.A1(_0185_),
    .A2(_0189_),
    .A3(_0197_),
    .B1(_0198_),
    .Y(_0201_));
 sky130_fd_sc_hd__or3_1 _0663_ (.A(_0191_),
    .B(_0196_),
    .C(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__o311a_1 _0664_ (.A1(_0185_),
    .A2(_0189_),
    .A3(_0197_),
    .B1(_0198_),
    .C1(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .X(_0203_));
 sky130_fd_sc_hd__xor2_1 _0665_ (.A(_0188_),
    .B(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__xnor2_1 _0666_ (.A(_0202_),
    .B(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__nor2_1 _0667_ (.A(_0163_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A3 ),
    .Y(_0206_));
 sky130_fd_sc_hd__nand2_1 _0668_ (.A(_0162_),
    .B(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__nor2_1 _0669_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B1 ),
    .B(_0206_),
    .Y(_0208_));
 sky130_fd_sc_hd__a21oi_1 _0670_ (.A1(_0207_),
    .A2(_0200_),
    .B1(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__nor2_1 _0671_ (.A(_0193_),
    .B(_0194_),
    .Y(_0210_));
 sky130_fd_sc_hd__o31a_1 _0672_ (.A1(_0191_),
    .A2(_0195_),
    .A3(_0201_),
    .B1(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__nor4_1 _0673_ (.A(_0210_),
    .B(_0191_),
    .C(_0195_),
    .D(_0201_),
    .Y(_0212_));
 sky130_fd_sc_hd__or3_1 _0674_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .B(_0211_),
    .C(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__o21a_1 _0675_ (.A1(_0211_),
    .A2(_0212_),
    .B1(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .X(_0214_));
 sky130_fd_sc_hd__a221o_1 _0676_ (.A1(_0167_),
    .A2(_0205_),
    .B1(_0209_),
    .B2(_0213_),
    .C1(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__nand2_1 _0677_ (.A(_0168_),
    .B(_0184_),
    .Y(_0216_));
 sky130_fd_sc_hd__or3b_1 _0678_ (.A(_0189_),
    .B(_0197_),
    .C_N(_0184_),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _0679_ (.A0(_0168_),
    .A1(_0216_),
    .S(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__o21a_1 _0680_ (.A1(_0167_),
    .A2(_0205_),
    .B1(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__inv_2 _0681_ (.A(_0207_),
    .Y(_0220_));
 sky130_fd_sc_hd__a211o_1 _0682_ (.A1(_0215_),
    .A2(_0219_),
    .B1(_0220_),
    .C1(_0208_),
    .X(_0221_));
 sky130_fd_sc_hd__xor2_2 _0683_ (.A(_0200_),
    .B(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__nor2_1 _0684_ (.A(_0211_),
    .B(_0212_),
    .Y(_0223_));
 sky130_fd_sc_hd__and2b_1 _0685_ (.A_N(\CIRCUIT_1957.int_memory_1.div_1.A4 ),
    .B(_0199_),
    .X(_0224_));
 sky130_fd_sc_hd__and2b_1 _0686_ (.A_N(_0199_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A4 ),
    .X(_0225_));
 sky130_fd_sc_hd__o311a_1 _0687_ (.A1(_0224_),
    .A2(_0208_),
    .A3(_0225_),
    .B1(_0207_),
    .C1(_0180_),
    .X(_0226_));
 sky130_fd_sc_hd__and2_1 _0688_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .B(_0209_),
    .X(_0227_));
 sky130_fd_sc_hd__a211oi_1 _0689_ (.A1(_0215_),
    .A2(_0219_),
    .B1(_0226_),
    .C1(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__xnor2_1 _0690_ (.A(_0223_),
    .B(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__nand2_1 _0691_ (.A(_0167_),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__clkbuf_4 _0692_ (.A(\CIRCUIT_1957.int_memory_1.div_1.B2 ),
    .X(_0231_));
 sky130_fd_sc_hd__nand2_1 _0693_ (.A(_0231_),
    .B(_0222_),
    .Y(_0232_));
 sky130_fd_sc_hd__nor2_1 _0694_ (.A(_0163_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A2 ),
    .Y(_0233_));
 sky130_fd_sc_hd__and2_1 _0695_ (.A(_0162_),
    .B(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__a21oi_1 _0696_ (.A1(_0215_),
    .A2(_0219_),
    .B1(_0163_),
    .Y(_0235_));
 sky130_fd_sc_hd__xnor2_2 _0697_ (.A(\CIRCUIT_1957.int_memory_1.div_1.A3 ),
    .B(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__or2_1 _0698_ (.A(_0162_),
    .B(_0233_),
    .X(_0237_));
 sky130_fd_sc_hd__o221ai_2 _0699_ (.A1(_0234_),
    .A2(_0236_),
    .B1(_0222_),
    .B2(_0231_),
    .C1(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _0700_ (.A(_0205_),
    .Y(_0239_));
 sky130_fd_sc_hd__nor2_1 _0701_ (.A(_0239_),
    .B(_0218_),
    .Y(_0240_));
 sky130_fd_sc_hd__a211o_1 _0702_ (.A1(_0207_),
    .A2(_0200_),
    .B1(_0208_),
    .C1(_0180_),
    .X(_0241_));
 sky130_fd_sc_hd__a21oi_1 _0703_ (.A1(_0223_),
    .A2(_0241_),
    .B1(_0226_),
    .Y(_0242_));
 sky130_fd_sc_hd__xnor2_1 _0704_ (.A(_0168_),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__mux2_1 _0705_ (.A0(_0239_),
    .A1(_0240_),
    .S(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__o21bai_1 _0706_ (.A1(_0167_),
    .A2(_0229_),
    .B1_N(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__a31o_2 _0707_ (.A1(_0230_),
    .A2(_0232_),
    .A3(_0238_),
    .B1(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__o21ai_1 _0708_ (.A1(_0234_),
    .A2(_0236_),
    .B1(_0237_),
    .Y(_0247_));
 sky130_fd_sc_hd__xnor2_1 _0709_ (.A(_0231_),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__nand2_1 _0710_ (.A(_0246_),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__xnor2_1 _0711_ (.A(_0222_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand2_1 _0712_ (.A(_0167_),
    .B(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__nand3b_1 _0713_ (.A_N(_0234_),
    .B(_0237_),
    .C(_0246_),
    .Y(_0252_));
 sky130_fd_sc_hd__xnor2_2 _0714_ (.A(_0236_),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__nand2_1 _0715_ (.A(_0231_),
    .B(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__nor2_1 _0716_ (.A(_0163_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A1 ),
    .Y(_0255_));
 sky130_fd_sc_hd__and2_1 _0717_ (.A(_0162_),
    .B(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__a21boi_1 _0718_ (.A1(_0166_),
    .A2(_0246_),
    .B1_N(\CIRCUIT_1957.int_memory_1.div_1.A2 ),
    .Y(_0257_));
 sky130_fd_sc_hd__a21oi_2 _0719_ (.A1(_0233_),
    .A2(_0246_),
    .B1(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__or2_1 _0720_ (.A(_0162_),
    .B(_0255_),
    .X(_0259_));
 sky130_fd_sc_hd__o221ai_2 _0721_ (.A1(_0256_),
    .A2(_0258_),
    .B1(_0253_),
    .B2(_0231_),
    .C1(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__nand2_1 _0722_ (.A(_0229_),
    .B(_0244_),
    .Y(_0261_));
 sky130_fd_sc_hd__and3_1 _0723_ (.A(_0168_),
    .B(_0232_),
    .C(_0238_),
    .X(_0262_));
 sky130_fd_sc_hd__a21oi_1 _0724_ (.A1(_0232_),
    .A2(_0238_),
    .B1(_0168_),
    .Y(_0263_));
 sky130_fd_sc_hd__nor2_1 _0725_ (.A(_0262_),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__mux2_1 _0726_ (.A0(_0229_),
    .A1(_0261_),
    .S(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__o21ai_1 _0727_ (.A1(_0167_),
    .A2(_0250_),
    .B1(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__a31o_2 _0728_ (.A1(_0251_),
    .A2(_0254_),
    .A3(_0260_),
    .B1(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__and3_1 _0729_ (.A(_0166_),
    .B(\CIRCUIT_1957.int_memory_1.div_1.A1 ),
    .C(_0267_),
    .X(_0268_));
 sky130_fd_sc_hd__a21oi_1 _0730_ (.A1(_0166_),
    .A2(_0267_),
    .B1(\CIRCUIT_1957.int_memory_1.div_1.A1 ),
    .Y(_0269_));
 sky130_fd_sc_hd__or2_1 _0731_ (.A(_0162_),
    .B(_0164_),
    .X(_0270_));
 sky130_fd_sc_hd__o31a_1 _0732_ (.A1(_0165_),
    .A2(_0268_),
    .A3(_0269_),
    .B1(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__nand2_1 _0733_ (.A(_0162_),
    .B(_0255_),
    .Y(_0272_));
 sky130_fd_sc_hd__a31o_1 _0734_ (.A1(_0272_),
    .A2(_0259_),
    .A3(_0267_),
    .B1(_0258_),
    .X(_0273_));
 sky130_fd_sc_hd__nand4_1 _0735_ (.A(_0272_),
    .B(_0258_),
    .C(_0259_),
    .D(_0267_),
    .Y(_0274_));
 sky130_fd_sc_hd__a21o_1 _0736_ (.A1(_0273_),
    .A2(_0274_),
    .B1(_0231_),
    .X(_0275_));
 sky130_fd_sc_hd__and3_1 _0737_ (.A(_0231_),
    .B(_0273_),
    .C(_0274_),
    .X(_0276_));
 sky130_fd_sc_hd__a21oi_1 _0738_ (.A1(_0271_),
    .A2(_0275_),
    .B1(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__o211ai_1 _0739_ (.A1(_0256_),
    .A2(_0258_),
    .B1(_0259_),
    .C1(_0267_),
    .Y(_0278_));
 sky130_fd_sc_hd__a21o_1 _0740_ (.A1(_0231_),
    .A2(_0267_),
    .B1(_0253_),
    .X(_0279_));
 sky130_fd_sc_hd__nand3_1 _0741_ (.A(_0231_),
    .B(_0253_),
    .C(_0267_),
    .Y(_0280_));
 sky130_fd_sc_hd__nand3_1 _0742_ (.A(_0278_),
    .B(_0279_),
    .C(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__a21o_1 _0743_ (.A1(_0279_),
    .A2(_0280_),
    .B1(_0278_),
    .X(_0282_));
 sky130_fd_sc_hd__inv_2 _0744_ (.A(_0250_),
    .Y(_0283_));
 sky130_fd_sc_hd__nor2_1 _0745_ (.A(_0283_),
    .B(_0265_),
    .Y(_0284_));
 sky130_fd_sc_hd__nand2_1 _0746_ (.A(_0254_),
    .B(_0260_),
    .Y(_0285_));
 sky130_fd_sc_hd__xnor2_1 _0747_ (.A(_0168_),
    .B(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__mux2_1 _0748_ (.A0(_0283_),
    .A1(_0284_),
    .S(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__a31o_1 _0749_ (.A1(_0168_),
    .A2(_0281_),
    .A3(_0282_),
    .B1(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__and2b_1 _0750_ (.A_N(_0277_),
    .B(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__nand2_1 _0751_ (.A(_0281_),
    .B(_0282_),
    .Y(_0290_));
 sky130_fd_sc_hd__a21o_1 _0752_ (.A1(_0281_),
    .A2(_0282_),
    .B1(_0168_),
    .X(_0291_));
 sky130_fd_sc_hd__a21o_2 _0753_ (.A1(_0291_),
    .A2(_0277_),
    .B1(_0288_),
    .X(_0292_));
 sky130_fd_sc_hd__a21oi_1 _0754_ (.A1(_0167_),
    .A2(_0292_),
    .B1(_0290_),
    .Y(_0293_));
 sky130_fd_sc_hd__a31o_1 _0755_ (.A1(_0167_),
    .A2(_0290_),
    .A3(_0287_),
    .B1(_0293_),
    .X(_0294_));
 sky130_fd_sc_hd__or2_1 _0756_ (.A(\CIRCUIT_1957.MEMORY_68.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_69.s_currentState ),
    .X(_0295_));
 sky130_fd_sc_hd__or2_2 _0757_ (.A(_0116_),
    .B(_0295_),
    .X(_0296_));
 sky130_fd_sc_hd__a21oi_1 _0758_ (.A1(_0289_),
    .A2(_0294_),
    .B1(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__o21a_1 _0759_ (.A1(_0289_),
    .A2(_0294_),
    .B1(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__nand2_1 _0760_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .Y(_0299_));
 sky130_fd_sc_hd__nand2_1 _0761_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .Y(_0300_));
 sky130_fd_sc_hd__a22oi_1 _0762_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .B1(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .B2(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .Y(_0301_));
 sky130_fd_sc_hd__o21ba_1 _0763_ (.A1(_0299_),
    .A2(_0300_),
    .B1_N(_0301_),
    .X(_0302_));
 sky130_fd_sc_hd__and2_1 _0764_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .X(_0303_));
 sky130_fd_sc_hd__and4_1 _0765_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .C(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .D(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .X(_0304_));
 sky130_fd_sc_hd__a31o_1 _0766_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .A3(_0303_),
    .B1(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__and3_1 _0767_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .C(_0303_),
    .X(_0306_));
 sky130_fd_sc_hd__a21oi_1 _0768_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .B1(_0303_),
    .Y(_0307_));
 sky130_fd_sc_hd__nor2_1 _0769_ (.A(_0306_),
    .B(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__and2_1 _0770_ (.A(_0305_),
    .B(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__nor2_1 _0771_ (.A(_0305_),
    .B(_0308_),
    .Y(_0310_));
 sky130_fd_sc_hd__or2_1 _0772_ (.A(_0309_),
    .B(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__xor2_1 _0773_ (.A(_0302_),
    .B(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_1 _0774_ (.A(_0303_),
    .B(_0304_),
    .Y(_0313_));
 sky130_fd_sc_hd__a22oi_1 _0775_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .B1(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .B2(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .Y(_0314_));
 sky130_fd_sc_hd__or2_1 _0776_ (.A(_0305_),
    .B(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__a21o_1 _0777_ (.A1(_0313_),
    .A2(_0315_),
    .B1(_0300_),
    .X(_0316_));
 sky130_fd_sc_hd__or2_1 _0778_ (.A(_0312_),
    .B(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__nand2_1 _0779_ (.A(_0312_),
    .B(_0316_),
    .Y(_0318_));
 sky130_fd_sc_hd__nand2b_1 _0780_ (.A_N(\CIRCUIT_1957.MEMORY_70.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_71.s_currentState ),
    .Y(_0319_));
 sky130_fd_sc_hd__nand2b_2 _0781_ (.A_N(\CIRCUIT_1957.MEMORY_68.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_69.s_currentState ),
    .Y(_0320_));
 sky130_fd_sc_hd__nor2_2 _0782_ (.A(_0319_),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__or2_2 _0783_ (.A(\CIRCUIT_1957.MEMORY_70.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_71.s_currentState ),
    .X(_0322_));
 sky130_fd_sc_hd__nor2_1 _0784_ (.A(_0295_),
    .B(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__nand2b_2 _0785_ (.A_N(\CIRCUIT_1957.MEMORY_69.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_68.s_currentState ),
    .Y(_0324_));
 sky130_fd_sc_hd__nor2_1 _0786_ (.A(_0324_),
    .B(_0322_),
    .Y(_0325_));
 sky130_fd_sc_hd__nand2b_2 _0787_ (.A_N(\CIRCUIT_1957.MEMORY_71.s_currentState ),
    .B(\CIRCUIT_1957.MEMORY_70.s_currentState ),
    .Y(_0326_));
 sky130_fd_sc_hd__nor2_2 _0788_ (.A(_0324_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__nor2_2 _0789_ (.A(_0117_),
    .B(_0322_),
    .Y(_0328_));
 sky130_fd_sc_hd__a22o_1 _0790_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[3] ),
    .A2(_0327_),
    .B1(_0328_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_6.input2[3] ),
    .X(_0329_));
 sky130_fd_sc_hd__a221o_1 _0791_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[3] ),
    .A2(_0323_),
    .B1(_0325_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_4.input2[3] ),
    .C1(_0329_),
    .X(_0330_));
 sky130_fd_sc_hd__nor2_2 _0792_ (.A(_0295_),
    .B(_0326_),
    .Y(_0331_));
 sky130_fd_sc_hd__nor2_2 _0793_ (.A(_0320_),
    .B(_0322_),
    .Y(_0332_));
 sky130_fd_sc_hd__nor2_2 _0794_ (.A(_0117_),
    .B(_0326_),
    .Y(_0333_));
 sky130_fd_sc_hd__nor2_2 _0795_ (.A(_0320_),
    .B(_0326_),
    .Y(_0334_));
 sky130_fd_sc_hd__a22o_1 _0796_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[3] ),
    .A2(_0333_),
    .B1(_0334_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_1.input2[3] ),
    .X(_0335_));
 sky130_fd_sc_hd__a221o_1 _0797_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[3] ),
    .A2(_0331_),
    .B1(_0332_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_5.input2[3] ),
    .C1(_0335_),
    .X(_0336_));
 sky130_fd_sc_hd__inv_2 _0798_ (.A(_0162_),
    .Y(_0337_));
 sky130_fd_sc_hd__or2_1 _0799_ (.A(_0116_),
    .B(_0320_),
    .X(_0338_));
 sky130_fd_sc_hd__inv_2 _0800_ (.A(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand2_1 _0801_ (.A(_0166_),
    .B(_0177_),
    .Y(_0340_));
 sky130_fd_sc_hd__nor2_1 _0802_ (.A(_0324_),
    .B(_0319_),
    .Y(_0341_));
 sky130_fd_sc_hd__nor2_1 _0803_ (.A(_0295_),
    .B(_0319_),
    .Y(_0342_));
 sky130_fd_sc_hd__a22o_1 _0804_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[3] ),
    .A2(_0341_),
    .B1(_0342_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_49.input2[3] ),
    .X(_0343_));
 sky130_fd_sc_hd__a41o_1 _0805_ (.A1(_0337_),
    .A2(_0169_),
    .A3(_0339_),
    .A4(_0340_),
    .B1(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__or3_1 _0806_ (.A(_0330_),
    .B(_0336_),
    .C(_0344_),
    .X(_0345_));
 sky130_fd_sc_hd__a31o_1 _0807_ (.A1(_0317_),
    .A2(_0318_),
    .A3(_0321_),
    .B1(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__or2_1 _0808_ (.A(_0117_),
    .B(_0319_),
    .X(_0347_));
 sky130_fd_sc_hd__a21oi_1 _0809_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .A2(_0305_),
    .B1(_0306_),
    .Y(_0348_));
 sky130_fd_sc_hd__a22oi_1 _0810_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .B1(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .B2(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .Y(_0349_));
 sky130_fd_sc_hd__and4_1 _0811_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .C(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .D(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .X(_0350_));
 sky130_fd_sc_hd__or3_1 _0812_ (.A(_0348_),
    .B(_0349_),
    .C(_0350_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_1 _0813_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_1 _0814_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .Y(_0353_));
 sky130_fd_sc_hd__a21oi_1 _0815_ (.A1(_0353_),
    .A2(_0351_),
    .B1(_0352_),
    .Y(_0354_));
 sky130_fd_sc_hd__a21oi_1 _0816_ (.A1(_0351_),
    .A2(_0352_),
    .B1(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__nor2_1 _0817_ (.A(_0349_),
    .B(_0350_),
    .Y(_0356_));
 sky130_fd_sc_hd__or2b_1 _0818_ (.A(_0356_),
    .B_N(_0348_),
    .X(_0357_));
 sky130_fd_sc_hd__xor2_1 _0819_ (.A(_0353_),
    .B(_0299_),
    .X(_0358_));
 sky130_fd_sc_hd__and2_1 _0820_ (.A(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .B(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .X(_0359_));
 sky130_fd_sc_hd__o21a_1 _0821_ (.A1(_0359_),
    .A2(_0309_),
    .B1(_0348_),
    .X(_0360_));
 sky130_fd_sc_hd__a2bb2o_1 _0822_ (.A1_N(_0353_),
    .A2_N(_0299_),
    .B1(_0358_),
    .B2(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_1 _0823_ (.A(_0351_),
    .B(_0357_),
    .Y(_0362_));
 sky130_fd_sc_hd__xnor2_1 _0824_ (.A(_0362_),
    .B(_0361_),
    .Y(_0363_));
 sky130_fd_sc_hd__and2_1 _0825_ (.A(_0358_),
    .B(_0360_),
    .X(_0364_));
 sky130_fd_sc_hd__nor2_1 _0826_ (.A(_0358_),
    .B(_0360_),
    .Y(_0365_));
 sky130_fd_sc_hd__or2_1 _0827_ (.A(_0364_),
    .B(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__o22a_1 _0828_ (.A1(_0299_),
    .A2(_0300_),
    .B1(_0301_),
    .B2(_0311_),
    .X(_0367_));
 sky130_fd_sc_hd__xnor2_1 _0829_ (.A(_0366_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__nor2_1 _0830_ (.A(_0317_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__o21bai_1 _0831_ (.A1(_0366_),
    .A2(_0367_),
    .B1_N(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__and2_1 _0832_ (.A(_0363_),
    .B(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__a31o_1 _0833_ (.A1(_0351_),
    .A2(_0357_),
    .A3(_0361_),
    .B1(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__a21oi_1 _0834_ (.A1(_0355_),
    .A2(_0372_),
    .B1(_0354_),
    .Y(_0373_));
 sky130_fd_sc_hd__nand2_1 _0835_ (.A(_0215_),
    .B(_0219_),
    .Y(_0374_));
 sky130_fd_sc_hd__nor2_2 _0836_ (.A(_0116_),
    .B(_0324_),
    .Y(_0375_));
 sky130_fd_sc_hd__a2bb2o_1 _0837_ (.A1_N(_0347_),
    .A2_N(_0373_),
    .B1(_0374_),
    .B2(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__or3_1 _0838_ (.A(_0298_),
    .B(_0346_),
    .C(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__a22o_2 _0839_ (.A1(_0115_),
    .A2(\CIRCUIT_1957.D3 ),
    .B1(_0377_),
    .B2(_0119_),
    .X(_0378_));
 sky130_fd_sc_hd__xnor2_1 _0840_ (.A(_0099_),
    .B(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _0841_ (.A(_0161_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__xnor2_1 _0842_ (.A(_0180_),
    .B(_0271_),
    .Y(_0381_));
 sky130_fd_sc_hd__and4_1 _0843_ (.A(_0273_),
    .B(_0274_),
    .C(_0292_),
    .D(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__a22oi_1 _0844_ (.A1(_0273_),
    .A2(_0274_),
    .B1(_0292_),
    .B2(_0381_),
    .Y(_0383_));
 sky130_fd_sc_hd__o21ba_1 _0845_ (.A1(_0382_),
    .A2(_0383_),
    .B1_N(_0296_),
    .X(_0384_));
 sky130_fd_sc_hd__xnor2_1 _0846_ (.A(_0355_),
    .B(_0372_),
    .Y(_0385_));
 sky130_fd_sc_hd__nor2_1 _0847_ (.A(_0347_),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a22o_1 _0848_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[2] ),
    .A2(_0327_),
    .B1(_0323_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_3.input2[2] ),
    .X(_0387_));
 sky130_fd_sc_hd__a221o_1 _0849_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[2] ),
    .A2(_0328_),
    .B1(_0325_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_4.input2[2] ),
    .C1(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__nand3_1 _0850_ (.A(_0300_),
    .B(_0313_),
    .C(_0315_),
    .Y(_0389_));
 sky130_fd_sc_hd__o21a_1 _0851_ (.A1(_0163_),
    .A2(\CIRCUIT_1957.int_memory_1.div_1.A6 ),
    .B1(_0174_),
    .X(_0390_));
 sky130_fd_sc_hd__a22o_1 _0852_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[2] ),
    .A2(_0331_),
    .B1(_0332_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_5.input2[2] ),
    .X(_0391_));
 sky130_fd_sc_hd__a221o_1 _0853_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[2] ),
    .A2(_0341_),
    .B1(_0342_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_49.input2[2] ),
    .C1(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__a31o_1 _0854_ (.A1(_0169_),
    .A2(_0390_),
    .A3(_0339_),
    .B1(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__a221o_1 _0855_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[2] ),
    .A2(_0333_),
    .B1(_0334_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_1.input2[2] ),
    .C1(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__a31o_1 _0856_ (.A1(_0316_),
    .A2(_0321_),
    .A3(_0389_),
    .B1(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__or3_1 _0857_ (.A(_0386_),
    .B(_0388_),
    .C(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__a211o_1 _0858_ (.A1(_0246_),
    .A2(_0375_),
    .B1(_0384_),
    .C1(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _0859_ (.A1(_0115_),
    .A2(\CIRCUIT_1957.D2 ),
    .B1(_0397_),
    .B2(_0119_),
    .X(_0398_));
 sky130_fd_sc_hd__xnor2_1 _0860_ (.A(_0099_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__and3_1 _0861_ (.A(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .B(_0160_),
    .C(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__inv_2 _0862_ (.A(net10),
    .Y(_0401_));
 sky130_fd_sc_hd__inv_2 _0863_ (.A(_0118_),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _0864_ (.A(_0165_),
    .Y(_0403_));
 sky130_fd_sc_hd__nor2_1 _0865_ (.A(_0268_),
    .B(_0269_),
    .Y(_0404_));
 sky130_fd_sc_hd__a41o_1 _0866_ (.A1(_0403_),
    .A2(_0270_),
    .A3(_0404_),
    .A4(_0292_),
    .B1(_0296_),
    .X(_0405_));
 sky130_fd_sc_hd__a31o_1 _0867_ (.A1(_0403_),
    .A2(_0270_),
    .A3(_0292_),
    .B1(_0404_),
    .X(_0406_));
 sky130_fd_sc_hd__and2b_1 _0868_ (.A_N(_0405_),
    .B(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__a22o_1 _0869_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[1] ),
    .A2(_0323_),
    .B1(_0334_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_1.input2[1] ),
    .X(_0408_));
 sky130_fd_sc_hd__a221o_1 _0870_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_4.input2[1] ),
    .A2(_0325_),
    .B1(_0342_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_49.input2[1] ),
    .C1(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__inv_2 _0871_ (.A(_0304_),
    .Y(_0410_));
 sky130_fd_sc_hd__a22o_1 _0872_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .B1(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .B2(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .X(_0411_));
 sky130_fd_sc_hd__a22o_1 _0873_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[1] ),
    .A2(_0331_),
    .B1(_0332_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_5.input2[1] ),
    .X(_0412_));
 sky130_fd_sc_hd__a221o_1 _0874_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[1] ),
    .A2(_0328_),
    .B1(_0333_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_2.input2[1] ),
    .C1(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__a31o_1 _0875_ (.A1(_0410_),
    .A2(_0321_),
    .A3(_0411_),
    .B1(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__a221o_1 _0876_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[1] ),
    .A2(_0327_),
    .B1(_0341_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_51.input2[1] ),
    .C1(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__xnor2_1 _0877_ (.A(_0363_),
    .B(_0370_),
    .Y(_0416_));
 sky130_fd_sc_hd__a2bb2o_1 _0878_ (.A1_N(_0347_),
    .A2_N(_0416_),
    .B1(_0339_),
    .B2(_0187_),
    .X(_0417_));
 sky130_fd_sc_hd__or3_1 _0879_ (.A(_0409_),
    .B(_0415_),
    .C(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__a21o_1 _0880_ (.A1(_0267_),
    .A2(_0375_),
    .B1(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__o21ai_1 _0881_ (.A1(_0407_),
    .A2(_0419_),
    .B1(_0119_),
    .Y(_0420_));
 sky130_fd_sc_hd__nand2_1 _0882_ (.A(_0115_),
    .B(\CIRCUIT_1957.D1 ),
    .Y(_0421_));
 sky130_fd_sc_hd__o311a_1 _0883_ (.A1(_0401_),
    .A2(_0115_),
    .A3(_0402_),
    .B1(_0420_),
    .C1(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__xnor2_1 _0884_ (.A(_0102_),
    .B(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__and2_1 _0885_ (.A(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .B(_0160_),
    .X(_0424_));
 sky130_fd_sc_hd__nand2_1 _0886_ (.A(_0423_),
    .B(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__nand2_1 _0887_ (.A(_0164_),
    .B(_0292_),
    .Y(_0426_));
 sky130_fd_sc_hd__a21bo_1 _0888_ (.A1(_0166_),
    .A2(_0292_),
    .B1_N(\CIRCUIT_1957.int_memory_1.div_1.A0 ),
    .X(_0427_));
 sky130_fd_sc_hd__a21oi_1 _0889_ (.A1(_0426_),
    .A2(_0427_),
    .B1(_0296_),
    .Y(_0428_));
 sky130_fd_sc_hd__or2_1 _0890_ (.A(_0347_),
    .B(_0369_),
    .X(_0429_));
 sky130_fd_sc_hd__a21oi_1 _0891_ (.A1(_0317_),
    .A2(_0368_),
    .B1(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__nor2_1 _0892_ (.A(_0201_),
    .B(_0338_),
    .Y(_0431_));
 sky130_fd_sc_hd__a32o_1 _0893_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .A2(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .A3(_0321_),
    .B1(_0331_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_7.input2[0] ),
    .X(_0432_));
 sky130_fd_sc_hd__a221o_1 _0894_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[0] ),
    .A2(_0327_),
    .B1(_0325_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_4.input2[0] ),
    .C1(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__a22o_1 _0895_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[0] ),
    .A2(_0323_),
    .B1(_0332_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_5.input2[0] ),
    .X(_0434_));
 sky130_fd_sc_hd__a221o_1 _0896_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[0] ),
    .A2(_0328_),
    .B1(_0342_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_49.input2[0] ),
    .C1(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__a211o_1 _0897_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_1.input2[0] ),
    .A2(_0334_),
    .B1(_0433_),
    .C1(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__a221o_1 _0898_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[0] ),
    .A2(_0333_),
    .B1(_0341_),
    .B2(\CIRCUIT_1957.int_memory_1.GATES_51.input2[0] ),
    .C1(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__a211o_1 _0899_ (.A1(_0292_),
    .A2(_0375_),
    .B1(_0431_),
    .C1(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__o31ai_2 _0900_ (.A1(_0428_),
    .A2(_0430_),
    .A3(_0438_),
    .B1(_0119_),
    .Y(_0439_));
 sky130_fd_sc_hd__inv_2 _0901_ (.A(net9),
    .Y(_0440_));
 sky130_fd_sc_hd__nand2_1 _0902_ (.A(_0115_),
    .B(\CIRCUIT_1957.D0 ),
    .Y(_0441_));
 sky130_fd_sc_hd__o31a_1 _0903_ (.A1(_0440_),
    .A2(_0115_),
    .A3(_0402_),
    .B1(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__a21o_1 _0904_ (.A1(_0439_),
    .A2(_0442_),
    .B1(_0102_),
    .X(_0443_));
 sky130_fd_sc_hd__nand3_1 _0905_ (.A(_0102_),
    .B(_0439_),
    .C(_0442_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand2_1 _0906_ (.A(\CIRCUIT_1957.MEMORY_65.s_currentState ),
    .B(_0160_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand3_1 _0907_ (.A(_0443_),
    .B(_0444_),
    .C(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__and2b_1 _0908_ (.A_N(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ),
    .B(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ),
    .X(_0447_));
 sky130_fd_sc_hd__nand2_1 _0909_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__mux2_1 _0910_ (.A0(\CIRCUIT_1957.MEMORY_64.s_currentState ),
    .A1(_0102_),
    .S(_0448_),
    .X(_0449_));
 sky130_fd_sc_hd__a21oi_1 _0911_ (.A1(_0443_),
    .A2(_0444_),
    .B1(_0445_),
    .Y(_0450_));
 sky130_fd_sc_hd__a21o_1 _0912_ (.A1(_0446_),
    .A2(_0449_),
    .B1(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__xor2_1 _0913_ (.A(_0423_),
    .B(_0424_),
    .X(_0452_));
 sky130_fd_sc_hd__nand2_1 _0914_ (.A(_0451_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand2_1 _0915_ (.A(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .B(_0160_),
    .Y(_0454_));
 sky130_fd_sc_hd__xor2_1 _0916_ (.A(_0399_),
    .B(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__a21oi_1 _0917_ (.A1(_0425_),
    .A2(_0453_),
    .B1(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__xor2_1 _0918_ (.A(_0161_),
    .B(_0379_),
    .X(_0457_));
 sky130_fd_sc_hd__o21ai_1 _0919_ (.A1(_0400_),
    .A2(_0456_),
    .B1(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__a21o_2 _0920_ (.A1(_0126_),
    .A2(_0160_),
    .B1(_0128_),
    .X(_0459_));
 sky130_fd_sc_hd__inv_2 _0921_ (.A(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__a21oi_1 _0922_ (.A1(_0380_),
    .A2(_0458_),
    .B1(_0460_),
    .Y(\CIRCUIT_1957.MEMORY_64.d ));
 sky130_fd_sc_hd__nand2_1 _0923_ (.A(_0443_),
    .B(_0445_),
    .Y(_0461_));
 sky130_fd_sc_hd__and2_1 _0924_ (.A(_0439_),
    .B(_0442_),
    .X(_0462_));
 sky130_fd_sc_hd__inv_2 _0925_ (.A(\CIRCUIT_1957.MEMORY_65.s_currentState ),
    .Y(_0463_));
 sky130_fd_sc_hd__or3b_1 _0926_ (.A(_0462_),
    .B(_0463_),
    .C_N(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .X(_0464_));
 sky130_fd_sc_hd__and2b_1 _0927_ (.A_N(_0450_),
    .B(_0446_),
    .X(_0465_));
 sky130_fd_sc_hd__o21ai_1 _0928_ (.A1(_0465_),
    .A2(_0449_),
    .B1(_0459_),
    .Y(_0466_));
 sky130_fd_sc_hd__a21oi_1 _0929_ (.A1(_0465_),
    .A2(_0449_),
    .B1(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__a41o_1 _0930_ (.A1(_0444_),
    .A2(_0460_),
    .A3(_0461_),
    .A4(_0464_),
    .B1(_0467_),
    .X(\CIRCUIT_1957.MEMORY_65.d ));
 sky130_fd_sc_hd__or2_1 _0931_ (.A(_0451_),
    .B(_0452_),
    .X(_0468_));
 sky130_fd_sc_hd__inv_2 _0932_ (.A(_0422_),
    .Y(_0469_));
 sky130_fd_sc_hd__a31o_1 _0933_ (.A1(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .A3(_0469_),
    .B1(_0459_),
    .X(_0470_));
 sky130_fd_sc_hd__a21oi_1 _0934_ (.A1(_0102_),
    .A2(_0422_),
    .B1(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__a21o_1 _0935_ (.A1(_0099_),
    .A2(_0469_),
    .B1(_0424_),
    .X(_0472_));
 sky130_fd_sc_hd__a32o_1 _0936_ (.A1(_0453_),
    .A2(_0459_),
    .A3(_0468_),
    .B1(_0471_),
    .B2(_0472_),
    .X(\CIRCUIT_1957.MEMORY_66.d ));
 sky130_fd_sc_hd__a31o_1 _0937_ (.A1(_0425_),
    .A2(_0453_),
    .A3(_0455_),
    .B1(_0460_),
    .X(_0473_));
 sky130_fd_sc_hd__inv_2 _0938_ (.A(_0398_),
    .Y(_0474_));
 sky130_fd_sc_hd__o21ai_1 _0939_ (.A1(_0102_),
    .A2(_0474_),
    .B1(_0454_),
    .Y(_0475_));
 sky130_fd_sc_hd__a31o_1 _0940_ (.A1(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .A3(_0398_),
    .B1(_0459_),
    .X(_0476_));
 sky130_fd_sc_hd__a21oi_1 _0941_ (.A1(_0102_),
    .A2(_0474_),
    .B1(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__a2bb2o_1 _0942_ (.A1_N(_0456_),
    .A2_N(_0473_),
    .B1(_0475_),
    .B2(_0477_),
    .X(\CIRCUIT_1957.MEMORY_67.d ));
 sky130_fd_sc_hd__nor2_1 _0943_ (.A(_0099_),
    .B(_0378_),
    .Y(_0478_));
 sky130_fd_sc_hd__a21oi_1 _0944_ (.A1(_0099_),
    .A2(_0378_),
    .B1(_0161_),
    .Y(_0479_));
 sky130_fd_sc_hd__a311o_1 _0945_ (.A1(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .A2(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .A3(_0378_),
    .B1(_0459_),
    .C1(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__o31a_1 _0946_ (.A1(_0400_),
    .A2(_0456_),
    .A3(_0457_),
    .B1(_0459_),
    .X(_0481_));
 sky130_fd_sc_hd__a2bb2o_1 _0947_ (.A1_N(_0478_),
    .A2_N(_0480_),
    .B1(_0481_),
    .B2(_0458_),
    .X(\CIRCUIT_1957.MEMORY_63.d ));
 sky130_fd_sc_hd__clkbuf_1 _0948_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .X(_0482_));
 sky130_fd_sc_hd__clkbuf_1 _0949_ (.A(_0482_),
    .X(\CIRCUIT_1957.clock_gen_2_1.GATES_3.result ));
 sky130_fd_sc_hd__and3_1 _0950_ (.A(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ),
    .B(_0099_),
    .C(_0120_),
    .X(_0483_));
 sky130_fd_sc_hd__clkbuf_1 _0951_ (.A(_0483_),
    .X(\CIRCUIT_1957.MEMORY_62.d ));
 sky130_fd_sc_hd__o21a_1 _0952_ (.A1(_0151_),
    .A2(_0159_),
    .B1(\CIRCUIT_1957.MEMORY_88.s_currentState ),
    .X(\CIRCUIT_1957.GATES_60.result ));
 sky130_fd_sc_hd__and3_1 _0953_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .B(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ),
    .C(_0151_),
    .X(_0484_));
 sky130_fd_sc_hd__and3_1 _0954_ (.A(_0154_),
    .B(\CIRCUIT_1957.dest_reg_sel_new_1.GATES_14.input2 ),
    .C(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__clkbuf_1 _0955_ (.A(_0485_),
    .X(\CIRCUIT_1957.GATES_42.result ));
 sky130_fd_sc_hd__and3_1 _0956_ (.A(_0128_),
    .B(_0127_),
    .C(_0149_),
    .X(_0486_));
 sky130_fd_sc_hd__clkbuf_1 _0957_ (.A(_0486_),
    .X(\CIRCUIT_1957.GATES_41.result ));
 sky130_fd_sc_hd__and2_1 _0958_ (.A(\CIRCUIT_1957.GATES_33.input2 ),
    .B(_0484_),
    .X(_0487_));
 sky130_fd_sc_hd__clkbuf_1 _0959_ (.A(_0487_),
    .X(\CIRCUIT_1957.GATES_40.result ));
 sky130_fd_sc_hd__and3_1 _0960_ (.A(_0154_),
    .B(_0156_),
    .C(_0484_),
    .X(_0488_));
 sky130_fd_sc_hd__clkbuf_1 _0961_ (.A(_0488_),
    .X(\CIRCUIT_1957.GATES_39.result ));
 sky130_fd_sc_hd__and3_1 _0962_ (.A(_0128_),
    .B(_0120_),
    .C(_0149_),
    .X(_0489_));
 sky130_fd_sc_hd__clkbuf_1 _0963_ (.A(_0489_),
    .X(\CIRCUIT_1957.GATES_38.result ));
 sky130_fd_sc_hd__mux2_1 _0964_ (.A0(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .A1(_0378_),
    .S(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .X(_0490_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0965_ (.A(_0490_),
    .X(\CIRCUIT_1957.GATES_35.result ));
 sky130_fd_sc_hd__mux2_1 _0966_ (.A0(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .A1(_0398_),
    .S(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .X(_0491_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0967_ (.A(_0491_),
    .X(\CIRCUIT_1957.GATES_30.result ));
 sky130_fd_sc_hd__mux2_1 _0968_ (.A0(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .A1(_0469_),
    .S(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .X(_0492_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0969_ (.A(_0492_),
    .X(\CIRCUIT_1957.GATES_28.result ));
 sky130_fd_sc_hd__inv_2 _0970_ (.A(_0462_),
    .Y(_0493_));
 sky130_fd_sc_hd__mux2_1 _0971_ (.A0(\CIRCUIT_1957.MEMORY_65.s_currentState ),
    .A1(_0493_),
    .S(\CIRCUIT_1957.MEMORY_62.s_currentState ),
    .X(_0494_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _0972_ (.A(_0494_),
    .X(\CIRCUIT_1957.GATES_27.result ));
 sky130_fd_sc_hd__and3_1 _0973_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .B(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ),
    .C(_0447_),
    .X(_0495_));
 sky130_fd_sc_hd__clkbuf_1 _0974_ (.A(_0495_),
    .X(\CIRCUIT_1957.GATES_10.result ));
 sky130_fd_sc_hd__a31o_1 _0975_ (.A1(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .A2(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ),
    .A3(_0460_),
    .B1(\CIRCUIT_1957.GATES_10.result ),
    .X(\CIRCUIT_1957.GATES_9.result ));
 sky130_fd_sc_hd__buf_2 _0976_ (.A(_0119_),
    .X(_0496_));
 sky130_fd_sc_hd__and3_2 _0977_ (.A(clknet_1_1__leaf__0142_),
    .B(_0496_),
    .C(_0327_),
    .X(_0497_));
 sky130_fd_sc_hd__buf_1 _0978_ (.A(_0497_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_21.result ));
 sky130_fd_sc_hd__buf_1 _0979_ (.A(clknet_1_0__leaf_clk),
    .X(_0498_));
 sky130_fd_sc_hd__and3_2 _0980_ (.A(clknet_1_0__leaf__0498_),
    .B(_0496_),
    .C(_0334_),
    .X(_0499_));
 sky130_fd_sc_hd__buf_1 _0981_ (.A(_0499_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_22.result ));
 sky130_fd_sc_hd__and3_2 _0982_ (.A(clknet_1_1__leaf__0498_),
    .B(_0496_),
    .C(_0333_),
    .X(_0500_));
 sky130_fd_sc_hd__buf_1 _0983_ (.A(_0500_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_23.result ));
 sky130_fd_sc_hd__and3_2 _0984_ (.A(clknet_1_1__leaf__0498_),
    .B(_0496_),
    .C(_0321_),
    .X(_0501_));
 sky130_fd_sc_hd__buf_1 _0985_ (.A(_0501_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_24.result ));
 sky130_fd_sc_hd__nand2_2 _0986_ (.A(clknet_1_1__leaf__0142_),
    .B(_0496_),
    .Y(_0502_));
 sky130_fd_sc_hd__nor2_2 _0987_ (.A(_0347_),
    .B(clknet_1_0__leaf__0502_),
    .Y(\CIRCUIT_1957.int_memory_1.GATES_25.result ));
 sky130_fd_sc_hd__nor2_2 _0988_ (.A(_0296_),
    .B(clknet_1_0__leaf__0502_),
    .Y(\CIRCUIT_1957.int_memory_1.GATES_26.result ));
 sky130_fd_sc_hd__and3_2 _0989_ (.A(clknet_1_1__leaf__0498_),
    .B(_0496_),
    .C(_0375_),
    .X(_0503_));
 sky130_fd_sc_hd__buf_1 _0990_ (.A(_0503_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_27.result ));
 sky130_fd_sc_hd__nor2_2 _0991_ (.A(_0338_),
    .B(clknet_1_1__leaf__0502_),
    .Y(\CIRCUIT_1957.int_memory_1.GATES_28.result ));
 sky130_fd_sc_hd__and3_2 _0992_ (.A(clknet_1_0__leaf__0498_),
    .B(_0496_),
    .C(_0323_),
    .X(_0504_));
 sky130_fd_sc_hd__buf_1 _0993_ (.A(_0504_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_29.result ));
 sky130_fd_sc_hd__and3_2 _0994_ (.A(clknet_1_0__leaf__0498_),
    .B(_0496_),
    .C(_0325_),
    .X(_0505_));
 sky130_fd_sc_hd__buf_1 _0995_ (.A(_0505_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_30.result ));
 sky130_fd_sc_hd__and3_2 _0996_ (.A(clknet_1_0__leaf__0498_),
    .B(_0496_),
    .C(_0332_),
    .X(_0506_));
 sky130_fd_sc_hd__buf_1 _0997_ (.A(_0506_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_31.result ));
 sky130_fd_sc_hd__and3_2 _0998_ (.A(clknet_1_0__leaf__0498_),
    .B(_0496_),
    .C(_0328_),
    .X(_0507_));
 sky130_fd_sc_hd__buf_1 _0999_ (.A(_0507_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_32.result ));
 sky130_fd_sc_hd__and3_2 _1000_ (.A(clknet_1_0__leaf__0498_),
    .B(_0119_),
    .C(_0331_),
    .X(_0508_));
 sky130_fd_sc_hd__buf_1 _1001_ (.A(_0508_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_33.result ));
 sky130_fd_sc_hd__and3_2 _1002_ (.A(clknet_1_1__leaf__0498_),
    .B(_0119_),
    .C(_0342_),
    .X(_0509_));
 sky130_fd_sc_hd__buf_1 _1003_ (.A(_0509_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_50.result ));
 sky130_fd_sc_hd__and3_2 _1004_ (.A(clknet_1_0__leaf_clk),
    .B(_0119_),
    .C(_0341_),
    .X(_0510_));
 sky130_fd_sc_hd__buf_1 _1005_ (.A(_0510_),
    .X(\CIRCUIT_1957.int_memory_1.GATES_53.result ));
 sky130_fd_sc_hd__clkbuf_4 _1006_ (.A(_0121_),
    .X(_0511_));
 sky130_fd_sc_hd__buf_2 _1007_ (.A(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__inv_2 _1008_ (.A(\CIRCUIT_1957.MEMORY_67.s_currentState ),
    .Y(_0513_));
 sky130_fd_sc_hd__nor2_2 _1009_ (.A(_0513_),
    .B(_0511_),
    .Y(_0514_));
 sky130_fd_sc_hd__clkbuf_4 _1010_ (.A(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__a21o_1 _1011_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[2] ),
    .A2(_0512_),
    .B1(_0515_),
    .X(_0027_));
 sky130_fd_sc_hd__inv_2 _1012_ (.A(\CIRCUIT_1957.MEMORY_63.s_currentState ),
    .Y(_0516_));
 sky130_fd_sc_hd__nor2_2 _1013_ (.A(_0516_),
    .B(_0511_),
    .Y(_0517_));
 sky130_fd_sc_hd__clkbuf_4 _1014_ (.A(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__a21o_1 _1015_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[3] ),
    .A2(_0512_),
    .B1(_0518_),
    .X(_0028_));
 sky130_fd_sc_hd__nor2_2 _1016_ (.A(_0463_),
    .B(_0511_),
    .Y(_0519_));
 sky130_fd_sc_hd__clkbuf_4 _1017_ (.A(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__a21o_1 _1018_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_4.input2[0] ),
    .A2(_0512_),
    .B1(_0520_),
    .X(_0029_));
 sky130_fd_sc_hd__inv_2 _1019_ (.A(\CIRCUIT_1957.MEMORY_66.s_currentState ),
    .Y(_0521_));
 sky130_fd_sc_hd__nor2_2 _1020_ (.A(_0521_),
    .B(_0511_),
    .Y(_0522_));
 sky130_fd_sc_hd__clkbuf_4 _1021_ (.A(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__a21o_1 _1022_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_4.input2[1] ),
    .A2(_0512_),
    .B1(_0523_),
    .X(_0030_));
 sky130_fd_sc_hd__a21o_1 _1023_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_4.input2[2] ),
    .A2(_0512_),
    .B1(_0515_),
    .X(_0031_));
 sky130_fd_sc_hd__a21o_1 _1024_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_4.input2[3] ),
    .A2(_0512_),
    .B1(_0518_),
    .X(_0032_));
 sky130_fd_sc_hd__a21o_1 _1025_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_5.input2[0] ),
    .A2(_0512_),
    .B1(_0520_),
    .X(_0033_));
 sky130_fd_sc_hd__a21o_1 _1026_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_5.input2[1] ),
    .A2(_0512_),
    .B1(_0523_),
    .X(_0034_));
 sky130_fd_sc_hd__a21o_1 _1027_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_5.input2[2] ),
    .A2(_0512_),
    .B1(_0515_),
    .X(_0035_));
 sky130_fd_sc_hd__a21o_1 _1028_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_5.input2[3] ),
    .A2(_0512_),
    .B1(_0518_),
    .X(_0036_));
 sky130_fd_sc_hd__buf_2 _1029_ (.A(_0511_),
    .X(_0524_));
 sky130_fd_sc_hd__a21o_1 _1030_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[0] ),
    .A2(_0524_),
    .B1(_0520_),
    .X(_0037_));
 sky130_fd_sc_hd__a21o_1 _1031_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[1] ),
    .A2(_0524_),
    .B1(_0523_),
    .X(_0038_));
 sky130_fd_sc_hd__a21o_1 _1032_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[2] ),
    .A2(_0524_),
    .B1(_0515_),
    .X(_0039_));
 sky130_fd_sc_hd__a21o_1 _1033_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_6.input2[3] ),
    .A2(_0524_),
    .B1(_0518_),
    .X(_0040_));
 sky130_fd_sc_hd__a21o_1 _1034_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[0] ),
    .A2(_0524_),
    .B1(_0520_),
    .X(_0041_));
 sky130_fd_sc_hd__a21o_1 _1035_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[1] ),
    .A2(_0524_),
    .B1(_0523_),
    .X(_0042_));
 sky130_fd_sc_hd__a21o_1 _1036_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[2] ),
    .A2(_0524_),
    .B1(_0515_),
    .X(_0043_));
 sky130_fd_sc_hd__a21o_1 _1037_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_7.input2[3] ),
    .A2(_0524_),
    .B1(_0518_),
    .X(_0044_));
 sky130_fd_sc_hd__a21o_1 _1038_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[0] ),
    .A2(_0524_),
    .B1(_0520_),
    .X(_0045_));
 sky130_fd_sc_hd__a21o_1 _1039_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[1] ),
    .A2(_0524_),
    .B1(_0523_),
    .X(_0046_));
 sky130_fd_sc_hd__buf_2 _1040_ (.A(_0511_),
    .X(_0525_));
 sky130_fd_sc_hd__a21o_1 _1041_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[2] ),
    .A2(_0525_),
    .B1(_0515_),
    .X(_0047_));
 sky130_fd_sc_hd__a21o_1 _1042_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_8.input2[3] ),
    .A2(_0525_),
    .B1(_0518_),
    .X(_0048_));
 sky130_fd_sc_hd__a21o_1 _1043_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_49.input2[0] ),
    .A2(_0525_),
    .B1(_0520_),
    .X(_0049_));
 sky130_fd_sc_hd__a21o_1 _1044_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_49.input2[1] ),
    .A2(_0525_),
    .B1(_0523_),
    .X(_0050_));
 sky130_fd_sc_hd__a21o_1 _1045_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_49.input2[2] ),
    .A2(_0525_),
    .B1(_0515_),
    .X(_0051_));
 sky130_fd_sc_hd__a21o_1 _1046_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_49.input2[3] ),
    .A2(_0525_),
    .B1(_0518_),
    .X(_0052_));
 sky130_fd_sc_hd__nand2_2 _1047_ (.A(_0141_),
    .B(clknet_1_1__leaf__0143_),
    .Y(_0000_));
 sky130_fd_sc_hd__buf_1 _1048_ (.A(clknet_1_1__leaf__0142_),
    .X(_0526_));
 sky130_fd_sc_hd__nand2_2 _1049_ (.A(_0141_),
    .B(clknet_1_1__leaf__0526_),
    .Y(_0001_));
 sky130_fd_sc_hd__clkinv_2 _1050_ (.A(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ),
    .Y(_0003_));
 sky130_fd_sc_hd__nand2_2 _1051_ (.A(_0141_),
    .B(clknet_1_1__leaf__0526_),
    .Y(_0004_));
 sky130_fd_sc_hd__nand2_2 _1052_ (.A(_0141_),
    .B(clknet_1_1__leaf__0526_),
    .Y(_0005_));
 sky130_fd_sc_hd__nand2_2 _1053_ (.A(_0141_),
    .B(clknet_1_1__leaf__0526_),
    .Y(_0006_));
 sky130_fd_sc_hd__nand2_2 _1054_ (.A(_0141_),
    .B(clknet_1_1__leaf__0526_),
    .Y(_0007_));
 sky130_fd_sc_hd__nand2_2 _1055_ (.A(_0141_),
    .B(clknet_1_1__leaf__0526_),
    .Y(_0008_));
 sky130_fd_sc_hd__nand2_2 _1056_ (.A(_0141_),
    .B(clknet_1_0__leaf__0526_),
    .Y(_0009_));
 sky130_fd_sc_hd__nand2_2 _1057_ (.A(_0141_),
    .B(clknet_1_0__leaf__0526_),
    .Y(_0010_));
 sky130_fd_sc_hd__nand2_2 _1058_ (.A(_0140_),
    .B(clknet_1_0__leaf__0526_),
    .Y(_0011_));
 sky130_fd_sc_hd__nand2_2 _1059_ (.A(_0140_),
    .B(clknet_1_0__leaf__0526_),
    .Y(_0012_));
 sky130_fd_sc_hd__nand2_2 _1060_ (.A(_0140_),
    .B(clknet_1_0__leaf__0142_),
    .Y(_0013_));
 sky130_fd_sc_hd__nand2_2 _1061_ (.A(_0140_),
    .B(clknet_1_0__leaf__0142_),
    .Y(_0014_));
 sky130_fd_sc_hd__nand2_2 _1062_ (.A(_0140_),
    .B(clknet_1_0__leaf__0142_),
    .Y(_0015_));
 sky130_fd_sc_hd__nand2_2 _1063_ (.A(_0140_),
    .B(clknet_1_1__leaf__0142_),
    .Y(_0016_));
 sky130_fd_sc_hd__nand2_2 _1064_ (.A(_0140_),
    .B(clknet_1_0__leaf__0142_),
    .Y(_0017_));
 sky130_fd_sc_hd__nand2_2 _1065_ (.A(_0140_),
    .B(clknet_1_0__leaf__0142_),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1067__2 (.A(clknet_1_0__leaf__0143_),
    .Y(net41));
 sky130_fd_sc_hd__inv_2 _1068__3 (.A(clknet_1_0__leaf__0143_),
    .Y(net42));
 sky130_fd_sc_hd__inv_2 _1069__4 (.A(clknet_1_0__leaf__0143_),
    .Y(net43));
 sky130_fd_sc_hd__inv_2 _1070__5 (.A(clknet_1_0__leaf__0143_),
    .Y(net44));
 sky130_fd_sc_hd__inv_2 _1071__6 (.A(clknet_1_1__leaf__0143_),
    .Y(net45));
 sky130_fd_sc_hd__inv_2 _1072__7 (.A(clknet_1_1__leaf__0143_),
    .Y(net46));
 sky130_fd_sc_hd__inv_2 _1073__8 (.A(clknet_1_1__leaf__0143_),
    .Y(net47));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__a21o_1 _1074_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[0] ),
    .A2(_0525_),
    .B1(_0520_),
    .X(_0061_));
 sky130_fd_sc_hd__a21o_1 _1075_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[1] ),
    .A2(_0525_),
    .B1(_0523_),
    .X(_0062_));
 sky130_fd_sc_hd__a21o_1 _1076_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[2] ),
    .A2(_0525_),
    .B1(_0515_),
    .X(_0063_));
 sky130_fd_sc_hd__a21o_1 _1077_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_51.input2[3] ),
    .A2(_0525_),
    .B1(_0518_),
    .X(_0064_));
 sky130_fd_sc_hd__or2_1 _1078_ (.A(net25),
    .B(net11),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_1 _1079_ (.A(_0527_),
    .X(_0065_));
 sky130_fd_sc_hd__and2b_1 _1080_ (.A_N(net11),
    .B(net21),
    .X(_0528_));
 sky130_fd_sc_hd__clkbuf_1 _1081_ (.A(_0528_),
    .X(_0066_));
 sky130_fd_sc_hd__and2b_1 _1082_ (.A_N(net11),
    .B(net22),
    .X(_0529_));
 sky130_fd_sc_hd__clkbuf_1 _1083_ (.A(_0529_),
    .X(_0067_));
 sky130_fd_sc_hd__and2b_1 _1084_ (.A_N(net11),
    .B(net24),
    .X(_0530_));
 sky130_fd_sc_hd__clkbuf_1 _1085_ (.A(_0530_),
    .X(_0068_));
 sky130_fd_sc_hd__buf_2 _1086_ (.A(_0511_),
    .X(_0531_));
 sky130_fd_sc_hd__a21o_1 _1087_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_1.input2[0] ),
    .A2(_0531_),
    .B1(_0520_),
    .X(_0069_));
 sky130_fd_sc_hd__a21o_1 _1088_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_1.input2[1] ),
    .A2(_0531_),
    .B1(_0523_),
    .X(_0070_));
 sky130_fd_sc_hd__a21o_1 _1089_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_1.input2[2] ),
    .A2(_0531_),
    .B1(_0515_),
    .X(_0071_));
 sky130_fd_sc_hd__a21o_1 _1090_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_1.input2[3] ),
    .A2(_0531_),
    .B1(_0518_),
    .X(_0072_));
 sky130_fd_sc_hd__a21o_1 _1091_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[0] ),
    .A2(_0531_),
    .B1(_0520_),
    .X(_0073_));
 sky130_fd_sc_hd__a21o_1 _1092_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[1] ),
    .A2(_0531_),
    .B1(_0523_),
    .X(_0074_));
 sky130_fd_sc_hd__a21o_1 _1093_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[2] ),
    .A2(_0531_),
    .B1(_0515_),
    .X(_0075_));
 sky130_fd_sc_hd__a21o_1 _1094_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_2.input2[3] ),
    .A2(_0531_),
    .B1(_0518_),
    .X(_0076_));
 sky130_fd_sc_hd__a21o_1 _1095_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ),
    .A2(_0531_),
    .B1(_0520_),
    .X(_0077_));
 sky130_fd_sc_hd__a21o_1 _1096_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ),
    .A2(_0531_),
    .B1(_0523_),
    .X(_0078_));
 sky130_fd_sc_hd__buf_2 _1097_ (.A(_0511_),
    .X(_0532_));
 sky130_fd_sc_hd__a21o_1 _1098_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ),
    .A2(_0532_),
    .B1(_0514_),
    .X(_0079_));
 sky130_fd_sc_hd__a21o_1 _1099_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ),
    .A2(_0532_),
    .B1(_0517_),
    .X(_0080_));
 sky130_fd_sc_hd__a21o_1 _1100_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ),
    .A2(_0532_),
    .B1(_0519_),
    .X(_0081_));
 sky130_fd_sc_hd__a21o_1 _1101_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ),
    .A2(_0532_),
    .B1(_0522_),
    .X(_0082_));
 sky130_fd_sc_hd__a21o_1 _1102_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ),
    .A2(_0532_),
    .B1(_0514_),
    .X(_0083_));
 sky130_fd_sc_hd__a21o_1 _1103_ (.A1(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ),
    .A2(_0532_),
    .B1(_0517_),
    .X(_0084_));
 sky130_fd_sc_hd__a21o_1 _1104_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A0 ),
    .A2(_0532_),
    .B1(_0519_),
    .X(_0085_));
 sky130_fd_sc_hd__a21o_1 _1105_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A1 ),
    .A2(_0532_),
    .B1(_0522_),
    .X(_0086_));
 sky130_fd_sc_hd__a21o_1 _1106_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A2 ),
    .A2(_0532_),
    .B1(_0514_),
    .X(_0087_));
 sky130_fd_sc_hd__a21o_1 _1107_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A3 ),
    .A2(_0532_),
    .B1(_0517_),
    .X(_0088_));
 sky130_fd_sc_hd__buf_2 _1108_ (.A(_0511_),
    .X(_0533_));
 sky130_fd_sc_hd__a21o_1 _1109_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A4 ),
    .A2(_0533_),
    .B1(_0519_),
    .X(_0089_));
 sky130_fd_sc_hd__a21o_1 _1110_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A5 ),
    .A2(_0533_),
    .B1(_0522_),
    .X(_0090_));
 sky130_fd_sc_hd__a21o_1 _1111_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A6 ),
    .A2(_0533_),
    .B1(_0514_),
    .X(_0091_));
 sky130_fd_sc_hd__a21o_1 _1112_ (.A1(\CIRCUIT_1957.int_memory_1.div_1.A7 ),
    .A2(_0533_),
    .B1(_0517_),
    .X(_0092_));
 sky130_fd_sc_hd__a21o_1 _1113_ (.A1(_0166_),
    .A2(_0533_),
    .B1(_0519_),
    .X(_0093_));
 sky130_fd_sc_hd__a21o_1 _1114_ (.A1(_0162_),
    .A2(_0533_),
    .B1(_0522_),
    .X(_0094_));
 sky130_fd_sc_hd__a21o_1 _1115_ (.A1(_0231_),
    .A2(_0533_),
    .B1(_0514_),
    .X(_0095_));
 sky130_fd_sc_hd__a21o_1 _1116_ (.A1(_0167_),
    .A2(_0533_),
    .B1(_0517_),
    .X(_0096_));
 sky130_fd_sc_hd__a21o_1 _1117_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[0] ),
    .A2(_0533_),
    .B1(_0519_),
    .X(_0097_));
 sky130_fd_sc_hd__a21o_1 _1118_ (.A1(\CIRCUIT_1957.int_memory_1.GATES_3.input2[1] ),
    .A2(_0533_),
    .B1(_0522_),
    .X(_0098_));
 sky130_fd_sc_hd__dfxtp_1 _1119_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .D(_0027_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_3.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1120_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .D(_0028_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_3.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1121_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .D(_0029_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_4.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1122_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .D(_0030_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_4.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1123_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .D(_0031_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_4.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1124_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .D(_0032_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_4.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1125_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .D(_0033_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_5.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1126_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .D(_0034_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_5.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1127_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .D(_0035_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_5.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1128_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .D(_0036_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_5.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1129_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .D(_0037_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_6.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1130_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .D(_0038_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_6.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1131_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .D(_0039_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_6.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1132_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .D(_0040_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_6.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1133_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .D(_0041_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_7.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1134_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .D(_0042_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_7.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1135_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .D(_0043_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_7.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1136_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .D(_0044_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_7.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1137_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .D(_0045_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_8.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1138_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .D(_0046_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_8.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1139_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .D(_0047_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_8.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1140_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .D(_0048_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_8.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1141_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .D(_0049_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_49.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1142_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .D(_0050_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_49.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1143_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .D(_0051_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_49.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1144_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .D(_0052_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_49.input2[3] ));
 sky130_fd_sc_hd__dfstp_1 _1145_ (.CLK(\CIRCUIT_1957.clock_gen_2_1.GATES_3.result ),
    .D(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.d ),
    .SET_B(_0000_),
    .Q(\CIRCUIT_1957.clock_gen_2_1.MEMORY_4.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _1146_ (.CLK(clknet_1_0__leaf_clk),
    .D(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.d ),
    .RESET_B(_0001_),
    .Q(\CIRCUIT_1957.clock_gen_2_1.MEMORY_5.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1147_ (.CLK(_0003_),
    .D(\CIRCUIT_1957.clock_gen_2_1.GATES_1.input2 ),
    .RESET_B(_0002_),
    .Q(\CIRCUIT_1957.clock_gen_2_1.MEMORY_6.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1148_ (.CLK(\CIRCUIT_1957.clock_gen_2_1.CLK1 ),
    .D(\CIRCUIT_1957.D0 ),
    .RESET_B(_0004_),
    .Q(\CIRCUIT_1957.inst_dec_1.MEMORY_21.s_currentState ));
 sky130_fd_sc_hd__dfrtp_4 _1149_ (.CLK(\CIRCUIT_1957.clock_gen_2_1.CLK1 ),
    .D(\CIRCUIT_1957.D1 ),
    .RESET_B(_0005_),
    .Q(\CIRCUIT_1957.inst_dec_1.MEMORY_22.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1150_ (.CLK(\CIRCUIT_1957.clock_gen_2_1.CLK1 ),
    .D(\CIRCUIT_1957.D2 ),
    .RESET_B(_0006_),
    .Q(\CIRCUIT_1957.inst_dec_1.MEMORY_23.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1151_ (.CLK(\CIRCUIT_1957.clock_gen_2_1.CLK1 ),
    .D(\CIRCUIT_1957.D3 ),
    .RESET_B(_0007_),
    .Q(\CIRCUIT_1957.inst_dec_1.MEMORY_24.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1152_ (.CLK(clknet_1_1__leaf_clk),
    .D(\CIRCUIT_1957.GATES_53.result ),
    .RESET_B(_0008_),
    .Q(\CIRCUIT_1957.MEMORY_88.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1153_ (.CLK(\CIRCUIT_1957.GATES_42.result ),
    .D(\CIRCUIT_1957.GATES_35.result ),
    .Q(\CIRCUIT_1957.MEMORY_87.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1154_ (.CLK(\CIRCUIT_1957.GATES_42.result ),
    .D(\CIRCUIT_1957.GATES_30.result ),
    .Q(\CIRCUIT_1957.MEMORY_86.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1155_ (.CLK(\CIRCUIT_1957.GATES_42.result ),
    .D(\CIRCUIT_1957.GATES_28.result ),
    .Q(\CIRCUIT_1957.MEMORY_85.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1156_ (.CLK(\CIRCUIT_1957.GATES_42.result ),
    .D(\CIRCUIT_1957.GATES_27.result ),
    .Q(\CIRCUIT_1957.MEMORY_84.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1157_ (.CLK(\CIRCUIT_1957.GATES_40.result ),
    .D(\CIRCUIT_1957.GATES_35.result ),
    .Q(\CIRCUIT_1957.MEMORY_83.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1158_ (.CLK(\CIRCUIT_1957.GATES_40.result ),
    .D(\CIRCUIT_1957.GATES_30.result ),
    .Q(\CIRCUIT_1957.MEMORY_82.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1159_ (.CLK(\CIRCUIT_1957.GATES_40.result ),
    .D(\CIRCUIT_1957.GATES_28.result ),
    .Q(\CIRCUIT_1957.MEMORY_81.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1160_ (.CLK(\CIRCUIT_1957.GATES_40.result ),
    .D(\CIRCUIT_1957.GATES_27.result ),
    .Q(\CIRCUIT_1957.MEMORY_80.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1161_ (.CLK(\CIRCUIT_1957.GATES_39.result ),
    .D(\CIRCUIT_1957.GATES_35.result ),
    .Q(\CIRCUIT_1957.MEMORY_79.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1162_ (.CLK(\CIRCUIT_1957.GATES_39.result ),
    .D(\CIRCUIT_1957.GATES_30.result ),
    .Q(\CIRCUIT_1957.MEMORY_78.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1163_ (.CLK(\CIRCUIT_1957.GATES_39.result ),
    .D(\CIRCUIT_1957.GATES_28.result ),
    .Q(\CIRCUIT_1957.MEMORY_77.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1164_ (.CLK(\CIRCUIT_1957.GATES_39.result ),
    .D(\CIRCUIT_1957.GATES_27.result ),
    .Q(\CIRCUIT_1957.MEMORY_76.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1165_ (.CLK(\CIRCUIT_1957.GATES_41.result ),
    .D(\CIRCUIT_1957.GATES_35.result ),
    .RESET_B(_0009_),
    .Q(\CIRCUIT_1957.MEMORY_75.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1166_ (.CLK(\CIRCUIT_1957.GATES_41.result ),
    .D(\CIRCUIT_1957.GATES_30.result ),
    .RESET_B(_0010_),
    .Q(\CIRCUIT_1957.MEMORY_74.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1167_ (.CLK(\CIRCUIT_1957.GATES_41.result ),
    .D(\CIRCUIT_1957.GATES_28.result ),
    .RESET_B(_0011_),
    .Q(\CIRCUIT_1957.MEMORY_73.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1168_ (.CLK(\CIRCUIT_1957.GATES_41.result ),
    .D(\CIRCUIT_1957.GATES_27.result ),
    .RESET_B(_0012_),
    .Q(\CIRCUIT_1957.MEMORY_72.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1169_ (.CLK(\CIRCUIT_1957.GATES_38.result ),
    .D(\CIRCUIT_1957.GATES_35.result ),
    .RESET_B(_0013_),
    .Q(\CIRCUIT_1957.MEMORY_71.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1170_ (.CLK(\CIRCUIT_1957.GATES_38.result ),
    .D(\CIRCUIT_1957.GATES_30.result ),
    .RESET_B(_0014_),
    .Q(\CIRCUIT_1957.MEMORY_70.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1171_ (.CLK(\CIRCUIT_1957.GATES_38.result ),
    .D(\CIRCUIT_1957.GATES_28.result ),
    .RESET_B(_0015_),
    .Q(\CIRCUIT_1957.MEMORY_69.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1172_ (.CLK(\CIRCUIT_1957.GATES_38.result ),
    .D(\CIRCUIT_1957.GATES_27.result ),
    .RESET_B(_0016_),
    .Q(\CIRCUIT_1957.MEMORY_68.s_currentState ));
 sky130_fd_sc_hd__dfxtp_2 _1173_ (.CLK(\CIRCUIT_1957.GATES_9.result ),
    .D(\CIRCUIT_1957.MEMORY_67.d ),
    .Q(\CIRCUIT_1957.MEMORY_67.s_currentState ));
 sky130_fd_sc_hd__dfxtp_2 _1174_ (.CLK(\CIRCUIT_1957.GATES_9.result ),
    .D(\CIRCUIT_1957.MEMORY_66.d ),
    .Q(\CIRCUIT_1957.MEMORY_66.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1175_ (.CLK(\CIRCUIT_1957.GATES_9.result ),
    .D(\CIRCUIT_1957.MEMORY_65.d ),
    .Q(\CIRCUIT_1957.MEMORY_65.s_currentState ));
 sky130_fd_sc_hd__dfrtp_1 _1176_ (.CLK(\CIRCUIT_1957.GATES_10.result ),
    .D(\CIRCUIT_1957.MEMORY_64.d ),
    .RESET_B(_0017_),
    .Q(\CIRCUIT_1957.MEMORY_64.s_currentState ));
 sky130_fd_sc_hd__dfxtp_2 _1177_ (.CLK(\CIRCUIT_1957.GATES_9.result ),
    .D(\CIRCUIT_1957.MEMORY_63.d ),
    .Q(\CIRCUIT_1957.MEMORY_63.s_currentState ));
 sky130_fd_sc_hd__dfrtp_2 _1178_ (.CLK(\CIRCUIT_1957.GATES_60.result ),
    .D(\CIRCUIT_1957.MEMORY_62.d ),
    .RESET_B(_0018_),
    .Q(\CIRCUIT_1957.MEMORY_62.s_currentState ));
 sky130_fd_sc_hd__dfxtp_1 _1179_ (.CLK(net40),
    .D(_0053_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _1180_ (.CLK(net41),
    .D(_0054_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _1181_ (.CLK(net42),
    .D(_0055_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _1182_ (.CLK(net43),
    .D(_0056_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _1183_ (.CLK(net44),
    .D(_0057_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _1184_ (.CLK(net45),
    .D(_0058_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _1185_ (.CLK(net46),
    .D(_0059_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _1186_ (.CLK(net47),
    .D(_0060_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _1187_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .D(_0061_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_51.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1188_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .D(_0062_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_51.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1189_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .D(_0063_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_51.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1190_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .D(_0064_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_51.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1191_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0065_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _1192_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0066_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _1193_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0067_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _1194_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0068_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _1195_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .D(_0069_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_1.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1196_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .D(_0070_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_1.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1197_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .D(_0071_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_1.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1198_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .D(_0072_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_1.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1199_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .D(_0073_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_2.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1200_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .D(_0074_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_2.input2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _1201_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .D(_0075_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_2.input2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _1202_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .D(_0076_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_2.input2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _1203_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .D(_0077_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.A0 ));
 sky130_fd_sc_hd__dfxtp_1 _1204_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .D(_0078_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.A1 ));
 sky130_fd_sc_hd__dfxtp_1 _1205_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .D(_0079_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.A2 ));
 sky130_fd_sc_hd__dfxtp_1 _1206_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .D(_0080_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.A3 ));
 sky130_fd_sc_hd__dfxtp_1 _1207_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .D(_0081_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.B0 ));
 sky130_fd_sc_hd__dfxtp_1 _1208_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .D(_0082_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.B1 ));
 sky130_fd_sc_hd__dfxtp_1 _1209_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .D(_0083_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.B2 ));
 sky130_fd_sc_hd__dfxtp_1 _1210_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .D(_0084_),
    .Q(\CIRCUIT_1957.int_memory_1.mul2_1.B3 ));
 sky130_fd_sc_hd__dfxtp_1 _1211_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .D(_0085_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A0 ));
 sky130_fd_sc_hd__dfxtp_1 _1212_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .D(_0086_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A1 ));
 sky130_fd_sc_hd__dfxtp_1 _1213_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .D(_0087_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A2 ));
 sky130_fd_sc_hd__dfxtp_1 _1214_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .D(_0088_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A3 ));
 sky130_fd_sc_hd__dfxtp_1 _1215_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .D(_0089_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A4 ));
 sky130_fd_sc_hd__dfxtp_1 _1216_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .D(_0090_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A5 ));
 sky130_fd_sc_hd__dfxtp_1 _1217_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .D(_0091_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A6 ));
 sky130_fd_sc_hd__dfxtp_1 _1218_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .D(_0092_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.A7 ));
 sky130_fd_sc_hd__dfxtp_1 _1219_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .D(_0093_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.B0 ));
 sky130_fd_sc_hd__dfxtp_2 _1220_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .D(_0094_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.B1 ));
 sky130_fd_sc_hd__dfxtp_2 _1221_ (.CLK(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .D(_0095_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.B2 ));
 sky130_fd_sc_hd__dfxtp_1 _1222_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .D(_0096_),
    .Q(\CIRCUIT_1957.int_memory_1.div_1.B3 ));
 sky130_fd_sc_hd__dfxtp_1 _1223_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .D(_0097_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_3.input2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _1224_ (.CLK(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .D(_0098_),
    .Q(\CIRCUIT_1957.int_memory_1.GATES_3.input2[1] ));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_39 (.HI(net39));
 sky130_fd_sc_hd__inv_2 _1066__1 (.A(clknet_1_0__leaf__0143_),
    .Y(net40));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_38 (.HI(net38));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(io_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(io_in[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(io_in[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(io_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(io_in[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(io_in[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(io_in[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(io_in[8]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(io_in[9]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(rst),
    .X(net11));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_2 output18 (.A(net18),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(io_out[3]));
 sky130_fd_sc_hd__conb_1 tholin_avalonsemi_5401_28 (.LO(net28));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_53.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_53.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_53.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_53.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_53.result ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0498_ (.A(_0498_),
    .X(clknet_0__0498_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0498_ (.A(clknet_0__0498_),
    .X(clknet_1_0__leaf__0498_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0498_ (.A(clknet_0__0498_),
    .X(clknet_1_1__leaf__0498_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_50.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_50.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_50.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_50.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_50.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_33.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_33.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_33.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_33.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_33.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_32.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_32.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_32.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_32.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_32.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_31.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_31.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_31.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_31.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_31.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_30.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_30.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_30.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_30.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_30.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_29.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_29.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_29.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_29.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_29.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_27.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_27.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_27.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_27.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_27.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_24.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_24.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_24.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_24.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_24.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_23.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_23.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_23.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_23.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_23.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_22.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_22.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_22.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_22.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_22.result ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0142_ (.A(_0142_),
    .X(clknet_0__0142_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0142_ (.A(clknet_0__0142_),
    .X(clknet_1_0__leaf__0142_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0142_ (.A(clknet_0__0142_),
    .X(clknet_1_1__leaf__0142_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0526_ (.A(_0526_),
    .X(clknet_0__0526_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0526_ (.A(clknet_0__0526_),
    .X(clknet_1_0__leaf__0526_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0526_ (.A(clknet_0__0526_),
    .X(clknet_1_1__leaf__0526_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0502_ (.A(_0502_),
    .X(clknet_0__0502_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0502_ (.A(clknet_0__0502_),
    .X(clknet_1_0__leaf__0502_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0502_ (.A(clknet_0__0502_),
    .X(clknet_1_1__leaf__0502_));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_28.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_28.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_28.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_28.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_28.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_26.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_26.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_26.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_26.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_26.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_25.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_25.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_25.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_25.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_25.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_CIRCUIT_1957.int_memory_1.GATES_21.result  (.A(\CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .X(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_CIRCUIT_1957.int_memory_1.GATES_21.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .X(\clknet_1_0__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_CIRCUIT_1957.int_memory_1.GATES_21.result  (.A(\clknet_0_CIRCUIT_1957.int_memory_1.GATES_21.result ),
    .X(\clknet_1_1__leaf_CIRCUIT_1957.int_memory_1.GATES_21.result ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__0143_ (.A(_0143_),
    .X(clknet_0__0143_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__0143_ (.A(clknet_0__0143_),
    .X(clknet_1_0__leaf__0143_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__0143_ (.A(clknet_0__0143_),
    .X(clknet_1_1__leaf__0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1012__A (.DIODE(\CIRCUIT_1957.MEMORY_63.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0964__A0 (.DIODE(\CIRCUIT_1957.MEMORY_63.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0945__A2 (.DIODE(\CIRCUIT_1957.MEMORY_63.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0622__A (.DIODE(\CIRCUIT_1957.MEMORY_63.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0572__A0 (.DIODE(\CIRCUIT_1957.MEMORY_63.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0536__C (.DIODE(\CIRCUIT_1957.MEMORY_63.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1019__A (.DIODE(\CIRCUIT_1957.MEMORY_66.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0968__A0 (.DIODE(\CIRCUIT_1957.MEMORY_66.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0933__A2 (.DIODE(\CIRCUIT_1957.MEMORY_66.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0885__A (.DIODE(\CIRCUIT_1957.MEMORY_66.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0580__A0 (.DIODE(\CIRCUIT_1957.MEMORY_66.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0536__A (.DIODE(\CIRCUIT_1957.MEMORY_66.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__A (.DIODE(\CIRCUIT_1957.MEMORY_67.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0966__A0 (.DIODE(\CIRCUIT_1957.MEMORY_67.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0940__A2 (.DIODE(\CIRCUIT_1957.MEMORY_67.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__A (.DIODE(\CIRCUIT_1957.MEMORY_67.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__A (.DIODE(\CIRCUIT_1957.MEMORY_67.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0576__A0 (.DIODE(\CIRCUIT_1957.MEMORY_67.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0536__D (.DIODE(\CIRCUIT_1957.MEMORY_67.s_currentState ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1002__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0976__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0900__B1 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0881__B1 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__B2 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__B2 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0560__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0600__S (.DIODE(_0144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0598__S (.DIODE(_0144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0596__S (.DIODE(_0144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0594__S (.DIODE(_0144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0962__C (.DIODE(_0149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__C (.DIODE(_0149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0617__A3 (.DIODE(_0149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0612__A (.DIODE(_0149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0606__A (.DIODE(_0149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0803__A (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__A (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__A (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__B (.DIODE(_0295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0793__B (.DIODE(_0322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__B (.DIODE(_0322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__B (.DIODE(_0322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0784__B (.DIODE(_0322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0795__B (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__B (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0792__B (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0788__B (.DIODE(_0326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__C (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0893__B1 (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0873__A2 (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__A2 (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__A2 (.DIODE(_0331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__C (.DIODE(_0333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__A2 (.DIODE(_0333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0874__B1 (.DIODE(_0333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__A2 (.DIODE(_0333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0796__A2 (.DIODE(_0333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__B (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__B (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__B (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__B (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0989__B (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__B (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__B (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0982__B (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__B (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0977__B (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__A (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__A (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__A (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1040__A (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1029__A (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1020__B (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1016__B (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__B (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__B (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1007__A (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__B1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__B1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__B1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__B1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__B1 (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__A (.DIODE(_0514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1089__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1076__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1041__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1027__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1011__B1 (.DIODE(_0515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1116__B1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__B1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1107__B1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1103__B1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1099__B1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1014__A (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1042__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1024__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1015__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1095__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1074__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1043__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1034__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1025__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1018__B1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__B1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__B1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__B1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__B1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__B1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__A (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1096__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1092__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1075__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1044__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1026__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1022__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__A2 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__A2 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__A2 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__A2 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__A2 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1034__A2 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__A2 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__A2 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__A2 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__A2 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1116__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1109__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(io_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(io_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(io_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA__1084__A_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__A_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1080__A_N (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1078__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__0609__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__0588__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__0590__A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1004__A (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__CLK (.DIODE(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__A (.DIODE(clknet_1_0__leaf__0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__A (.DIODE(clknet_1_0__leaf__0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__A (.DIODE(clknet_1_0__leaf__0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__A (.DIODE(clknet_1_0__leaf__0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__A (.DIODE(clknet_1_0__leaf__0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__A (.DIODE(clknet_1_0__leaf__0498_));
 sky130_fd_sc_hd__decap_4 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_297 ();
 assign io_oeb = net38;
 assign io_out[22] = net34;
 assign io_out[23] = net35;
 assign io_out[24] = net36;
 assign io_out[25] = net37;
 assign io_out[26] = net39;
 assign io_out[4] = net28;
 assign io_out[5] = net29;
 assign io_out[6] = net30;
 assign io_out[7] = net31;
 assign io_out[8] = net32;
 assign io_out[9] = net33;
endmodule

