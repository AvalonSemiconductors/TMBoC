VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as512512512
  CLASS BLOCK ;
  FOREIGN wrapped_as512512512 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1800.000 BY 3100.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1470.200 1800.000 1470.800 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 38.120 1800.000 38.720 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 568.520 1800.000 569.120 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 621.560 1800.000 622.160 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 674.600 1800.000 675.200 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 727.640 1800.000 728.240 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 780.680 1800.000 781.280 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 833.720 1800.000 834.320 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 886.760 1800.000 887.360 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 939.800 1800.000 940.400 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 992.840 1800.000 993.440 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1045.880 1800.000 1046.480 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 91.160 1800.000 91.760 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1098.920 1800.000 1099.520 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1151.960 1800.000 1152.560 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1205.000 1800.000 1205.600 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1258.040 1800.000 1258.640 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1311.080 1800.000 1311.680 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1364.120 1800.000 1364.720 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1417.160 1800.000 1417.760 ;
    END
  END io_in[26]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 144.200 1800.000 144.800 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 197.240 1800.000 197.840 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 250.280 1800.000 250.880 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 303.320 1800.000 303.920 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 356.360 1800.000 356.960 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 409.400 1800.000 410.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 462.440 1800.000 463.040 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 515.480 1800.000 516.080 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 3061.400 1800.000 3062.000 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1576.280 1800.000 1576.880 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2106.680 1800.000 2107.280 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2159.720 1800.000 2160.320 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2212.760 1800.000 2213.360 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2265.800 1800.000 2266.400 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2318.840 1800.000 2319.440 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2371.880 1800.000 2372.480 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2424.920 1800.000 2425.520 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2477.960 1800.000 2478.560 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2531.000 1800.000 2531.600 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2584.040 1800.000 2584.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1629.320 1800.000 1629.920 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2637.080 1800.000 2637.680 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2690.120 1800.000 2690.720 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2743.160 1800.000 2743.760 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2796.200 1800.000 2796.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2849.240 1800.000 2849.840 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2902.280 1800.000 2902.880 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2955.320 1800.000 2955.920 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 3008.360 1800.000 3008.960 ;
    END
  END io_out[27]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1682.360 1800.000 1682.960 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1735.400 1800.000 1736.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1788.440 1800.000 1789.040 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1841.480 1800.000 1842.080 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1894.520 1800.000 1895.120 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1947.560 1800.000 1948.160 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2000.600 1800.000 2001.200 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 2053.640 1800.000 2054.240 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1796.000 1523.240 1800.000 1523.840 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 3087.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 3087.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 3087.440 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 3085.785 1794.650 3087.390 ;
        RECT 5.330 3080.345 1794.650 3083.175 ;
        RECT 5.330 3074.905 1794.650 3077.735 ;
        RECT 5.330 3069.465 1794.650 3072.295 ;
        RECT 5.330 3064.025 1794.650 3066.855 ;
        RECT 5.330 3058.585 1794.650 3061.415 ;
        RECT 5.330 3053.145 1794.650 3055.975 ;
        RECT 5.330 3047.705 1794.650 3050.535 ;
        RECT 5.330 3042.265 1794.650 3045.095 ;
        RECT 5.330 3036.825 1794.650 3039.655 ;
        RECT 5.330 3031.385 1794.650 3034.215 ;
        RECT 5.330 3025.945 1794.650 3028.775 ;
        RECT 5.330 3020.505 1794.650 3023.335 ;
        RECT 5.330 3015.065 1794.650 3017.895 ;
        RECT 5.330 3009.625 1794.650 3012.455 ;
        RECT 5.330 3004.185 1794.650 3007.015 ;
        RECT 5.330 2998.745 1794.650 3001.575 ;
        RECT 5.330 2993.305 1794.650 2996.135 ;
        RECT 5.330 2987.865 1794.650 2990.695 ;
        RECT 5.330 2982.425 1794.650 2985.255 ;
        RECT 5.330 2976.985 1794.650 2979.815 ;
        RECT 5.330 2971.545 1794.650 2974.375 ;
        RECT 5.330 2966.105 1794.650 2968.935 ;
        RECT 5.330 2960.665 1794.650 2963.495 ;
        RECT 5.330 2955.225 1794.650 2958.055 ;
        RECT 5.330 2949.785 1794.650 2952.615 ;
        RECT 5.330 2944.345 1794.650 2947.175 ;
        RECT 5.330 2938.905 1794.650 2941.735 ;
        RECT 5.330 2933.465 1794.650 2936.295 ;
        RECT 5.330 2928.025 1794.650 2930.855 ;
        RECT 5.330 2922.585 1794.650 2925.415 ;
        RECT 5.330 2917.145 1794.650 2919.975 ;
        RECT 5.330 2911.705 1794.650 2914.535 ;
        RECT 5.330 2906.265 1794.650 2909.095 ;
        RECT 5.330 2900.825 1794.650 2903.655 ;
        RECT 5.330 2895.385 1794.650 2898.215 ;
        RECT 5.330 2889.945 1794.650 2892.775 ;
        RECT 5.330 2884.505 1794.650 2887.335 ;
        RECT 5.330 2879.065 1794.650 2881.895 ;
        RECT 5.330 2873.625 1794.650 2876.455 ;
        RECT 5.330 2868.185 1794.650 2871.015 ;
        RECT 5.330 2862.745 1794.650 2865.575 ;
        RECT 5.330 2857.305 1794.650 2860.135 ;
        RECT 5.330 2851.865 1794.650 2854.695 ;
        RECT 5.330 2846.425 1794.650 2849.255 ;
        RECT 5.330 2840.985 1794.650 2843.815 ;
        RECT 5.330 2835.545 1794.650 2838.375 ;
        RECT 5.330 2830.105 1794.650 2832.935 ;
        RECT 5.330 2824.665 1794.650 2827.495 ;
        RECT 5.330 2819.225 1794.650 2822.055 ;
        RECT 5.330 2813.785 1794.650 2816.615 ;
        RECT 5.330 2808.345 1794.650 2811.175 ;
        RECT 5.330 2802.905 1794.650 2805.735 ;
        RECT 5.330 2797.465 1794.650 2800.295 ;
        RECT 5.330 2792.025 1794.650 2794.855 ;
        RECT 5.330 2786.585 1794.650 2789.415 ;
        RECT 5.330 2781.145 1794.650 2783.975 ;
        RECT 5.330 2775.705 1794.650 2778.535 ;
        RECT 5.330 2770.265 1794.650 2773.095 ;
        RECT 5.330 2764.825 1794.650 2767.655 ;
        RECT 5.330 2759.385 1794.650 2762.215 ;
        RECT 5.330 2753.945 1794.650 2756.775 ;
        RECT 5.330 2748.505 1794.650 2751.335 ;
        RECT 5.330 2743.065 1794.650 2745.895 ;
        RECT 5.330 2737.625 1794.650 2740.455 ;
        RECT 5.330 2732.185 1794.650 2735.015 ;
        RECT 5.330 2726.745 1794.650 2729.575 ;
        RECT 5.330 2721.305 1794.650 2724.135 ;
        RECT 5.330 2715.865 1794.650 2718.695 ;
        RECT 5.330 2710.425 1794.650 2713.255 ;
        RECT 5.330 2704.985 1794.650 2707.815 ;
        RECT 5.330 2699.545 1794.650 2702.375 ;
        RECT 5.330 2694.105 1794.650 2696.935 ;
        RECT 5.330 2688.665 1794.650 2691.495 ;
        RECT 5.330 2683.225 1794.650 2686.055 ;
        RECT 5.330 2677.785 1794.650 2680.615 ;
        RECT 5.330 2672.345 1794.650 2675.175 ;
        RECT 5.330 2666.905 1794.650 2669.735 ;
        RECT 5.330 2661.465 1794.650 2664.295 ;
        RECT 5.330 2656.025 1794.650 2658.855 ;
        RECT 5.330 2650.585 1794.650 2653.415 ;
        RECT 5.330 2645.145 1794.650 2647.975 ;
        RECT 5.330 2639.705 1794.650 2642.535 ;
        RECT 5.330 2634.265 1794.650 2637.095 ;
        RECT 5.330 2628.825 1794.650 2631.655 ;
        RECT 5.330 2623.385 1794.650 2626.215 ;
        RECT 5.330 2617.945 1794.650 2620.775 ;
        RECT 5.330 2612.505 1794.650 2615.335 ;
        RECT 5.330 2607.065 1794.650 2609.895 ;
        RECT 5.330 2601.625 1794.650 2604.455 ;
        RECT 5.330 2596.185 1794.650 2599.015 ;
        RECT 5.330 2590.745 1794.650 2593.575 ;
        RECT 5.330 2585.305 1794.650 2588.135 ;
        RECT 5.330 2579.865 1794.650 2582.695 ;
        RECT 5.330 2574.425 1794.650 2577.255 ;
        RECT 5.330 2568.985 1794.650 2571.815 ;
        RECT 5.330 2563.545 1794.650 2566.375 ;
        RECT 5.330 2558.105 1794.650 2560.935 ;
        RECT 5.330 2552.665 1794.650 2555.495 ;
        RECT 5.330 2547.225 1794.650 2550.055 ;
        RECT 5.330 2541.785 1794.650 2544.615 ;
        RECT 5.330 2536.345 1794.650 2539.175 ;
        RECT 5.330 2530.905 1794.650 2533.735 ;
        RECT 5.330 2525.465 1794.650 2528.295 ;
        RECT 5.330 2520.025 1794.650 2522.855 ;
        RECT 5.330 2514.585 1794.650 2517.415 ;
        RECT 5.330 2509.145 1794.650 2511.975 ;
        RECT 5.330 2503.705 1794.650 2506.535 ;
        RECT 5.330 2498.265 1794.650 2501.095 ;
        RECT 5.330 2492.825 1794.650 2495.655 ;
        RECT 5.330 2487.385 1794.650 2490.215 ;
        RECT 5.330 2481.945 1794.650 2484.775 ;
        RECT 5.330 2476.505 1794.650 2479.335 ;
        RECT 5.330 2471.065 1794.650 2473.895 ;
        RECT 5.330 2465.625 1794.650 2468.455 ;
        RECT 5.330 2460.185 1794.650 2463.015 ;
        RECT 5.330 2454.745 1794.650 2457.575 ;
        RECT 5.330 2449.305 1794.650 2452.135 ;
        RECT 5.330 2443.865 1794.650 2446.695 ;
        RECT 5.330 2438.425 1794.650 2441.255 ;
        RECT 5.330 2432.985 1794.650 2435.815 ;
        RECT 5.330 2427.545 1794.650 2430.375 ;
        RECT 5.330 2422.105 1794.650 2424.935 ;
        RECT 5.330 2416.665 1794.650 2419.495 ;
        RECT 5.330 2411.225 1794.650 2414.055 ;
        RECT 5.330 2405.785 1794.650 2408.615 ;
        RECT 5.330 2400.345 1794.650 2403.175 ;
        RECT 5.330 2394.905 1794.650 2397.735 ;
        RECT 5.330 2389.465 1794.650 2392.295 ;
        RECT 5.330 2384.025 1794.650 2386.855 ;
        RECT 5.330 2378.585 1794.650 2381.415 ;
        RECT 5.330 2373.145 1794.650 2375.975 ;
        RECT 5.330 2367.705 1794.650 2370.535 ;
        RECT 5.330 2362.265 1794.650 2365.095 ;
        RECT 5.330 2356.825 1794.650 2359.655 ;
        RECT 5.330 2351.385 1794.650 2354.215 ;
        RECT 5.330 2345.945 1794.650 2348.775 ;
        RECT 5.330 2340.505 1794.650 2343.335 ;
        RECT 5.330 2335.065 1794.650 2337.895 ;
        RECT 5.330 2329.625 1794.650 2332.455 ;
        RECT 5.330 2324.185 1794.650 2327.015 ;
        RECT 5.330 2318.745 1794.650 2321.575 ;
        RECT 5.330 2313.305 1794.650 2316.135 ;
        RECT 5.330 2307.865 1794.650 2310.695 ;
        RECT 5.330 2302.425 1794.650 2305.255 ;
        RECT 5.330 2296.985 1794.650 2299.815 ;
        RECT 5.330 2291.545 1794.650 2294.375 ;
        RECT 5.330 2286.105 1794.650 2288.935 ;
        RECT 5.330 2280.665 1794.650 2283.495 ;
        RECT 5.330 2275.225 1794.650 2278.055 ;
        RECT 5.330 2269.785 1794.650 2272.615 ;
        RECT 5.330 2264.345 1794.650 2267.175 ;
        RECT 5.330 2258.905 1794.650 2261.735 ;
        RECT 5.330 2253.465 1794.650 2256.295 ;
        RECT 5.330 2248.025 1794.650 2250.855 ;
        RECT 5.330 2242.585 1794.650 2245.415 ;
        RECT 5.330 2237.145 1794.650 2239.975 ;
        RECT 5.330 2231.705 1794.650 2234.535 ;
        RECT 5.330 2226.265 1794.650 2229.095 ;
        RECT 5.330 2220.825 1794.650 2223.655 ;
        RECT 5.330 2215.385 1794.650 2218.215 ;
        RECT 5.330 2209.945 1794.650 2212.775 ;
        RECT 5.330 2204.505 1794.650 2207.335 ;
        RECT 5.330 2199.065 1794.650 2201.895 ;
        RECT 5.330 2193.625 1794.650 2196.455 ;
        RECT 5.330 2188.185 1794.650 2191.015 ;
        RECT 5.330 2182.745 1794.650 2185.575 ;
        RECT 5.330 2177.305 1794.650 2180.135 ;
        RECT 5.330 2171.865 1794.650 2174.695 ;
        RECT 5.330 2166.425 1794.650 2169.255 ;
        RECT 5.330 2160.985 1794.650 2163.815 ;
        RECT 5.330 2155.545 1794.650 2158.375 ;
        RECT 5.330 2150.105 1794.650 2152.935 ;
        RECT 5.330 2144.665 1794.650 2147.495 ;
        RECT 5.330 2139.225 1794.650 2142.055 ;
        RECT 5.330 2133.785 1794.650 2136.615 ;
        RECT 5.330 2128.345 1794.650 2131.175 ;
        RECT 5.330 2122.905 1794.650 2125.735 ;
        RECT 5.330 2117.465 1794.650 2120.295 ;
        RECT 5.330 2112.025 1794.650 2114.855 ;
        RECT 5.330 2106.585 1794.650 2109.415 ;
        RECT 5.330 2101.145 1794.650 2103.975 ;
        RECT 5.330 2095.705 1794.650 2098.535 ;
        RECT 5.330 2090.265 1794.650 2093.095 ;
        RECT 5.330 2084.825 1794.650 2087.655 ;
        RECT 5.330 2079.385 1794.650 2082.215 ;
        RECT 5.330 2073.945 1794.650 2076.775 ;
        RECT 5.330 2068.505 1794.650 2071.335 ;
        RECT 5.330 2063.065 1794.650 2065.895 ;
        RECT 5.330 2057.625 1794.650 2060.455 ;
        RECT 5.330 2052.185 1794.650 2055.015 ;
        RECT 5.330 2046.745 1794.650 2049.575 ;
        RECT 5.330 2041.305 1794.650 2044.135 ;
        RECT 5.330 2035.865 1794.650 2038.695 ;
        RECT 5.330 2030.425 1794.650 2033.255 ;
        RECT 5.330 2024.985 1794.650 2027.815 ;
        RECT 5.330 2019.545 1794.650 2022.375 ;
        RECT 5.330 2014.105 1794.650 2016.935 ;
        RECT 5.330 2008.665 1794.650 2011.495 ;
        RECT 5.330 2003.225 1794.650 2006.055 ;
        RECT 5.330 1997.785 1794.650 2000.615 ;
        RECT 5.330 1992.345 1794.650 1995.175 ;
        RECT 5.330 1986.905 1794.650 1989.735 ;
        RECT 5.330 1981.465 1794.650 1984.295 ;
        RECT 5.330 1976.025 1794.650 1978.855 ;
        RECT 5.330 1970.585 1794.650 1973.415 ;
        RECT 5.330 1965.145 1794.650 1967.975 ;
        RECT 5.330 1959.705 1794.650 1962.535 ;
        RECT 5.330 1954.265 1794.650 1957.095 ;
        RECT 5.330 1948.825 1794.650 1951.655 ;
        RECT 5.330 1943.385 1794.650 1946.215 ;
        RECT 5.330 1937.945 1794.650 1940.775 ;
        RECT 5.330 1932.505 1794.650 1935.335 ;
        RECT 5.330 1927.065 1794.650 1929.895 ;
        RECT 5.330 1921.625 1794.650 1924.455 ;
        RECT 5.330 1916.185 1794.650 1919.015 ;
        RECT 5.330 1910.745 1794.650 1913.575 ;
        RECT 5.330 1905.305 1794.650 1908.135 ;
        RECT 5.330 1899.865 1794.650 1902.695 ;
        RECT 5.330 1894.425 1794.650 1897.255 ;
        RECT 5.330 1888.985 1794.650 1891.815 ;
        RECT 5.330 1883.545 1794.650 1886.375 ;
        RECT 5.330 1878.105 1794.650 1880.935 ;
        RECT 5.330 1872.665 1794.650 1875.495 ;
        RECT 5.330 1867.225 1794.650 1870.055 ;
        RECT 5.330 1861.785 1794.650 1864.615 ;
        RECT 5.330 1856.345 1794.650 1859.175 ;
        RECT 5.330 1850.905 1794.650 1853.735 ;
        RECT 5.330 1845.465 1794.650 1848.295 ;
        RECT 5.330 1840.025 1794.650 1842.855 ;
        RECT 5.330 1834.585 1794.650 1837.415 ;
        RECT 5.330 1829.145 1794.650 1831.975 ;
        RECT 5.330 1823.705 1794.650 1826.535 ;
        RECT 5.330 1818.265 1794.650 1821.095 ;
        RECT 5.330 1812.825 1794.650 1815.655 ;
        RECT 5.330 1807.385 1794.650 1810.215 ;
        RECT 5.330 1801.945 1794.650 1804.775 ;
        RECT 5.330 1796.505 1794.650 1799.335 ;
        RECT 5.330 1791.065 1794.650 1793.895 ;
        RECT 5.330 1785.625 1794.650 1788.455 ;
        RECT 5.330 1780.185 1794.650 1783.015 ;
        RECT 5.330 1774.745 1794.650 1777.575 ;
        RECT 5.330 1769.305 1794.650 1772.135 ;
        RECT 5.330 1763.865 1794.650 1766.695 ;
        RECT 5.330 1758.425 1794.650 1761.255 ;
        RECT 5.330 1752.985 1794.650 1755.815 ;
        RECT 5.330 1747.545 1794.650 1750.375 ;
        RECT 5.330 1742.105 1794.650 1744.935 ;
        RECT 5.330 1736.665 1794.650 1739.495 ;
        RECT 5.330 1731.225 1794.650 1734.055 ;
        RECT 5.330 1725.785 1794.650 1728.615 ;
        RECT 5.330 1720.345 1794.650 1723.175 ;
        RECT 5.330 1714.905 1794.650 1717.735 ;
        RECT 5.330 1709.465 1794.650 1712.295 ;
        RECT 5.330 1704.025 1794.650 1706.855 ;
        RECT 5.330 1698.585 1794.650 1701.415 ;
        RECT 5.330 1693.145 1794.650 1695.975 ;
        RECT 5.330 1687.705 1794.650 1690.535 ;
        RECT 5.330 1682.265 1794.650 1685.095 ;
        RECT 5.330 1676.825 1794.650 1679.655 ;
        RECT 5.330 1671.385 1794.650 1674.215 ;
        RECT 5.330 1665.945 1794.650 1668.775 ;
        RECT 5.330 1660.505 1794.650 1663.335 ;
        RECT 5.330 1655.065 1794.650 1657.895 ;
        RECT 5.330 1649.625 1794.650 1652.455 ;
        RECT 5.330 1644.185 1794.650 1647.015 ;
        RECT 5.330 1638.745 1794.650 1641.575 ;
        RECT 5.330 1633.305 1794.650 1636.135 ;
        RECT 5.330 1627.865 1794.650 1630.695 ;
        RECT 5.330 1622.425 1794.650 1625.255 ;
        RECT 5.330 1616.985 1794.650 1619.815 ;
        RECT 5.330 1611.545 1794.650 1614.375 ;
        RECT 5.330 1606.105 1794.650 1608.935 ;
        RECT 5.330 1600.665 1794.650 1603.495 ;
        RECT 5.330 1595.225 1794.650 1598.055 ;
        RECT 5.330 1589.785 1794.650 1592.615 ;
        RECT 5.330 1584.345 1794.650 1587.175 ;
        RECT 5.330 1578.905 1794.650 1581.735 ;
        RECT 5.330 1573.465 1794.650 1576.295 ;
        RECT 5.330 1568.025 1794.650 1570.855 ;
        RECT 5.330 1562.585 1794.650 1565.415 ;
        RECT 5.330 1557.145 1794.650 1559.975 ;
        RECT 5.330 1551.705 1794.650 1554.535 ;
        RECT 5.330 1546.265 1794.650 1549.095 ;
        RECT 5.330 1540.825 1794.650 1543.655 ;
        RECT 5.330 1535.385 1794.650 1538.215 ;
        RECT 5.330 1529.945 1794.650 1532.775 ;
        RECT 5.330 1524.505 1794.650 1527.335 ;
        RECT 5.330 1519.065 1794.650 1521.895 ;
        RECT 5.330 1513.625 1794.650 1516.455 ;
        RECT 5.330 1508.185 1794.650 1511.015 ;
        RECT 5.330 1502.745 1794.650 1505.575 ;
        RECT 5.330 1497.305 1794.650 1500.135 ;
        RECT 5.330 1491.865 1794.650 1494.695 ;
        RECT 5.330 1486.425 1794.650 1489.255 ;
        RECT 5.330 1480.985 1794.650 1483.815 ;
        RECT 5.330 1475.545 1794.650 1478.375 ;
        RECT 5.330 1470.105 1794.650 1472.935 ;
        RECT 5.330 1464.665 1794.650 1467.495 ;
        RECT 5.330 1459.225 1794.650 1462.055 ;
        RECT 5.330 1453.785 1794.650 1456.615 ;
        RECT 5.330 1448.345 1794.650 1451.175 ;
        RECT 5.330 1442.905 1794.650 1445.735 ;
        RECT 5.330 1437.465 1794.650 1440.295 ;
        RECT 5.330 1432.025 1794.650 1434.855 ;
        RECT 5.330 1426.585 1794.650 1429.415 ;
        RECT 5.330 1421.145 1794.650 1423.975 ;
        RECT 5.330 1415.705 1794.650 1418.535 ;
        RECT 5.330 1410.265 1794.650 1413.095 ;
        RECT 5.330 1404.825 1794.650 1407.655 ;
        RECT 5.330 1399.385 1794.650 1402.215 ;
        RECT 5.330 1393.945 1794.650 1396.775 ;
        RECT 5.330 1388.505 1794.650 1391.335 ;
        RECT 5.330 1383.065 1794.650 1385.895 ;
        RECT 5.330 1377.625 1794.650 1380.455 ;
        RECT 5.330 1372.185 1794.650 1375.015 ;
        RECT 5.330 1366.745 1794.650 1369.575 ;
        RECT 5.330 1361.305 1794.650 1364.135 ;
        RECT 5.330 1355.865 1794.650 1358.695 ;
        RECT 5.330 1350.425 1794.650 1353.255 ;
        RECT 5.330 1344.985 1794.650 1347.815 ;
        RECT 5.330 1339.545 1794.650 1342.375 ;
        RECT 5.330 1334.105 1794.650 1336.935 ;
        RECT 5.330 1328.665 1794.650 1331.495 ;
        RECT 5.330 1323.225 1794.650 1326.055 ;
        RECT 5.330 1317.785 1794.650 1320.615 ;
        RECT 5.330 1312.345 1794.650 1315.175 ;
        RECT 5.330 1306.905 1794.650 1309.735 ;
        RECT 5.330 1301.465 1794.650 1304.295 ;
        RECT 5.330 1296.025 1794.650 1298.855 ;
        RECT 5.330 1290.585 1794.650 1293.415 ;
        RECT 5.330 1285.145 1794.650 1287.975 ;
        RECT 5.330 1279.705 1794.650 1282.535 ;
        RECT 5.330 1274.265 1794.650 1277.095 ;
        RECT 5.330 1268.825 1794.650 1271.655 ;
        RECT 5.330 1263.385 1794.650 1266.215 ;
        RECT 5.330 1257.945 1794.650 1260.775 ;
        RECT 5.330 1252.505 1794.650 1255.335 ;
        RECT 5.330 1247.065 1794.650 1249.895 ;
        RECT 5.330 1241.625 1794.650 1244.455 ;
        RECT 5.330 1236.185 1794.650 1239.015 ;
        RECT 5.330 1230.745 1794.650 1233.575 ;
        RECT 5.330 1225.305 1794.650 1228.135 ;
        RECT 5.330 1219.865 1794.650 1222.695 ;
        RECT 5.330 1214.425 1794.650 1217.255 ;
        RECT 5.330 1208.985 1794.650 1211.815 ;
        RECT 5.330 1203.545 1794.650 1206.375 ;
        RECT 5.330 1198.105 1794.650 1200.935 ;
        RECT 5.330 1192.665 1794.650 1195.495 ;
        RECT 5.330 1187.225 1794.650 1190.055 ;
        RECT 5.330 1181.785 1794.650 1184.615 ;
        RECT 5.330 1176.345 1794.650 1179.175 ;
        RECT 5.330 1170.905 1794.650 1173.735 ;
        RECT 5.330 1165.465 1794.650 1168.295 ;
        RECT 5.330 1160.025 1794.650 1162.855 ;
        RECT 5.330 1154.585 1794.650 1157.415 ;
        RECT 5.330 1149.145 1794.650 1151.975 ;
        RECT 5.330 1143.705 1794.650 1146.535 ;
        RECT 5.330 1138.265 1794.650 1141.095 ;
        RECT 5.330 1132.825 1794.650 1135.655 ;
        RECT 5.330 1127.385 1794.650 1130.215 ;
        RECT 5.330 1121.945 1794.650 1124.775 ;
        RECT 5.330 1116.505 1794.650 1119.335 ;
        RECT 5.330 1111.065 1794.650 1113.895 ;
        RECT 5.330 1105.625 1794.650 1108.455 ;
        RECT 5.330 1100.185 1794.650 1103.015 ;
        RECT 5.330 1094.745 1794.650 1097.575 ;
        RECT 5.330 1089.305 1794.650 1092.135 ;
        RECT 5.330 1083.865 1794.650 1086.695 ;
        RECT 5.330 1078.425 1794.650 1081.255 ;
        RECT 5.330 1072.985 1794.650 1075.815 ;
        RECT 5.330 1067.545 1794.650 1070.375 ;
        RECT 5.330 1062.105 1794.650 1064.935 ;
        RECT 5.330 1056.665 1794.650 1059.495 ;
        RECT 5.330 1051.225 1794.650 1054.055 ;
        RECT 5.330 1045.785 1794.650 1048.615 ;
        RECT 5.330 1040.345 1794.650 1043.175 ;
        RECT 5.330 1034.905 1794.650 1037.735 ;
        RECT 5.330 1029.465 1794.650 1032.295 ;
        RECT 5.330 1024.025 1794.650 1026.855 ;
        RECT 5.330 1018.585 1794.650 1021.415 ;
        RECT 5.330 1013.145 1794.650 1015.975 ;
        RECT 5.330 1007.705 1794.650 1010.535 ;
        RECT 5.330 1002.265 1794.650 1005.095 ;
        RECT 5.330 996.825 1794.650 999.655 ;
        RECT 5.330 991.385 1794.650 994.215 ;
        RECT 5.330 985.945 1794.650 988.775 ;
        RECT 5.330 980.505 1794.650 983.335 ;
        RECT 5.330 975.065 1794.650 977.895 ;
        RECT 5.330 969.625 1794.650 972.455 ;
        RECT 5.330 964.185 1794.650 967.015 ;
        RECT 5.330 958.745 1794.650 961.575 ;
        RECT 5.330 953.305 1794.650 956.135 ;
        RECT 5.330 947.865 1794.650 950.695 ;
        RECT 5.330 942.425 1794.650 945.255 ;
        RECT 5.330 936.985 1794.650 939.815 ;
        RECT 5.330 931.545 1794.650 934.375 ;
        RECT 5.330 926.105 1794.650 928.935 ;
        RECT 5.330 920.665 1794.650 923.495 ;
        RECT 5.330 915.225 1794.650 918.055 ;
        RECT 5.330 909.785 1794.650 912.615 ;
        RECT 5.330 904.345 1794.650 907.175 ;
        RECT 5.330 898.905 1794.650 901.735 ;
        RECT 5.330 893.465 1794.650 896.295 ;
        RECT 5.330 888.025 1794.650 890.855 ;
        RECT 5.330 882.585 1794.650 885.415 ;
        RECT 5.330 877.145 1794.650 879.975 ;
        RECT 5.330 871.705 1794.650 874.535 ;
        RECT 5.330 866.265 1794.650 869.095 ;
        RECT 5.330 860.825 1794.650 863.655 ;
        RECT 5.330 855.385 1794.650 858.215 ;
        RECT 5.330 849.945 1794.650 852.775 ;
        RECT 5.330 844.505 1794.650 847.335 ;
        RECT 5.330 839.065 1794.650 841.895 ;
        RECT 5.330 833.625 1794.650 836.455 ;
        RECT 5.330 828.185 1794.650 831.015 ;
        RECT 5.330 822.745 1794.650 825.575 ;
        RECT 5.330 817.305 1794.650 820.135 ;
        RECT 5.330 811.865 1794.650 814.695 ;
        RECT 5.330 806.425 1794.650 809.255 ;
        RECT 5.330 800.985 1794.650 803.815 ;
        RECT 5.330 795.545 1794.650 798.375 ;
        RECT 5.330 790.105 1794.650 792.935 ;
        RECT 5.330 784.665 1794.650 787.495 ;
        RECT 5.330 779.225 1794.650 782.055 ;
        RECT 5.330 773.785 1794.650 776.615 ;
        RECT 5.330 768.345 1794.650 771.175 ;
        RECT 5.330 762.905 1794.650 765.735 ;
        RECT 5.330 757.465 1794.650 760.295 ;
        RECT 5.330 752.025 1794.650 754.855 ;
        RECT 5.330 746.585 1794.650 749.415 ;
        RECT 5.330 741.145 1794.650 743.975 ;
        RECT 5.330 735.705 1794.650 738.535 ;
        RECT 5.330 730.265 1794.650 733.095 ;
        RECT 5.330 724.825 1794.650 727.655 ;
        RECT 5.330 719.385 1794.650 722.215 ;
        RECT 5.330 713.945 1794.650 716.775 ;
        RECT 5.330 708.505 1794.650 711.335 ;
        RECT 5.330 703.065 1794.650 705.895 ;
        RECT 5.330 697.625 1794.650 700.455 ;
        RECT 5.330 692.185 1794.650 695.015 ;
        RECT 5.330 686.745 1794.650 689.575 ;
        RECT 5.330 681.305 1794.650 684.135 ;
        RECT 5.330 675.865 1794.650 678.695 ;
        RECT 5.330 670.425 1794.650 673.255 ;
        RECT 5.330 664.985 1794.650 667.815 ;
        RECT 5.330 659.545 1794.650 662.375 ;
        RECT 5.330 654.105 1794.650 656.935 ;
        RECT 5.330 648.665 1794.650 651.495 ;
        RECT 5.330 643.225 1794.650 646.055 ;
        RECT 5.330 637.785 1794.650 640.615 ;
        RECT 5.330 632.345 1794.650 635.175 ;
        RECT 5.330 626.905 1794.650 629.735 ;
        RECT 5.330 621.465 1794.650 624.295 ;
        RECT 5.330 616.025 1794.650 618.855 ;
        RECT 5.330 610.585 1794.650 613.415 ;
        RECT 5.330 605.145 1794.650 607.975 ;
        RECT 5.330 599.705 1794.650 602.535 ;
        RECT 5.330 594.265 1794.650 597.095 ;
        RECT 5.330 588.825 1794.650 591.655 ;
        RECT 5.330 583.385 1794.650 586.215 ;
        RECT 5.330 577.945 1794.650 580.775 ;
        RECT 5.330 572.505 1794.650 575.335 ;
        RECT 5.330 567.065 1794.650 569.895 ;
        RECT 5.330 561.625 1794.650 564.455 ;
        RECT 5.330 556.185 1794.650 559.015 ;
        RECT 5.330 550.745 1794.650 553.575 ;
        RECT 5.330 545.305 1794.650 548.135 ;
        RECT 5.330 539.865 1794.650 542.695 ;
        RECT 5.330 534.425 1794.650 537.255 ;
        RECT 5.330 528.985 1794.650 531.815 ;
        RECT 5.330 523.545 1794.650 526.375 ;
        RECT 5.330 518.105 1794.650 520.935 ;
        RECT 5.330 512.665 1794.650 515.495 ;
        RECT 5.330 507.225 1794.650 510.055 ;
        RECT 5.330 501.785 1794.650 504.615 ;
        RECT 5.330 496.345 1794.650 499.175 ;
        RECT 5.330 490.905 1794.650 493.735 ;
        RECT 5.330 485.465 1794.650 488.295 ;
        RECT 5.330 480.025 1794.650 482.855 ;
        RECT 5.330 474.585 1794.650 477.415 ;
        RECT 5.330 469.145 1794.650 471.975 ;
        RECT 5.330 463.705 1794.650 466.535 ;
        RECT 5.330 458.265 1794.650 461.095 ;
        RECT 5.330 452.825 1794.650 455.655 ;
        RECT 5.330 447.385 1794.650 450.215 ;
        RECT 5.330 441.945 1794.650 444.775 ;
        RECT 5.330 436.505 1794.650 439.335 ;
        RECT 5.330 431.065 1794.650 433.895 ;
        RECT 5.330 425.625 1794.650 428.455 ;
        RECT 5.330 420.185 1794.650 423.015 ;
        RECT 5.330 414.745 1794.650 417.575 ;
        RECT 5.330 409.305 1794.650 412.135 ;
        RECT 5.330 403.865 1794.650 406.695 ;
        RECT 5.330 398.425 1794.650 401.255 ;
        RECT 5.330 392.985 1794.650 395.815 ;
        RECT 5.330 387.545 1794.650 390.375 ;
        RECT 5.330 382.105 1794.650 384.935 ;
        RECT 5.330 376.665 1794.650 379.495 ;
        RECT 5.330 371.225 1794.650 374.055 ;
        RECT 5.330 365.785 1794.650 368.615 ;
        RECT 5.330 360.345 1794.650 363.175 ;
        RECT 5.330 354.905 1794.650 357.735 ;
        RECT 5.330 349.465 1794.650 352.295 ;
        RECT 5.330 344.025 1794.650 346.855 ;
        RECT 5.330 338.585 1794.650 341.415 ;
        RECT 5.330 333.145 1794.650 335.975 ;
        RECT 5.330 327.705 1794.650 330.535 ;
        RECT 5.330 322.265 1794.650 325.095 ;
        RECT 5.330 316.825 1794.650 319.655 ;
        RECT 5.330 311.385 1794.650 314.215 ;
        RECT 5.330 305.945 1794.650 308.775 ;
        RECT 5.330 300.505 1794.650 303.335 ;
        RECT 5.330 295.065 1794.650 297.895 ;
        RECT 5.330 289.625 1794.650 292.455 ;
        RECT 5.330 284.185 1794.650 287.015 ;
        RECT 5.330 278.745 1794.650 281.575 ;
        RECT 5.330 273.305 1794.650 276.135 ;
        RECT 5.330 267.865 1794.650 270.695 ;
        RECT 5.330 262.425 1794.650 265.255 ;
        RECT 5.330 256.985 1794.650 259.815 ;
        RECT 5.330 251.545 1794.650 254.375 ;
        RECT 5.330 246.105 1794.650 248.935 ;
        RECT 5.330 240.665 1794.650 243.495 ;
        RECT 5.330 235.225 1794.650 238.055 ;
        RECT 5.330 229.785 1794.650 232.615 ;
        RECT 5.330 224.345 1794.650 227.175 ;
        RECT 5.330 218.905 1794.650 221.735 ;
        RECT 5.330 213.465 1794.650 216.295 ;
        RECT 5.330 208.025 1794.650 210.855 ;
        RECT 5.330 202.585 1794.650 205.415 ;
        RECT 5.330 197.145 1794.650 199.975 ;
        RECT 5.330 191.705 1794.650 194.535 ;
        RECT 5.330 186.265 1794.650 189.095 ;
        RECT 5.330 180.825 1794.650 183.655 ;
        RECT 5.330 175.385 1794.650 178.215 ;
        RECT 5.330 169.945 1794.650 172.775 ;
        RECT 5.330 164.505 1794.650 167.335 ;
        RECT 5.330 159.065 1794.650 161.895 ;
        RECT 5.330 153.625 1794.650 156.455 ;
        RECT 5.330 148.185 1794.650 151.015 ;
        RECT 5.330 142.745 1794.650 145.575 ;
        RECT 5.330 137.305 1794.650 140.135 ;
        RECT 5.330 131.865 1794.650 134.695 ;
        RECT 5.330 126.425 1794.650 129.255 ;
        RECT 5.330 120.985 1794.650 123.815 ;
        RECT 5.330 115.545 1794.650 118.375 ;
        RECT 5.330 110.105 1794.650 112.935 ;
        RECT 5.330 104.665 1794.650 107.495 ;
        RECT 5.330 99.225 1794.650 102.055 ;
        RECT 5.330 93.785 1794.650 96.615 ;
        RECT 5.330 88.345 1794.650 91.175 ;
        RECT 5.330 82.905 1794.650 85.735 ;
        RECT 5.330 77.465 1794.650 80.295 ;
        RECT 5.330 72.025 1794.650 74.855 ;
        RECT 5.330 66.585 1794.650 69.415 ;
        RECT 5.330 61.145 1794.650 63.975 ;
        RECT 5.330 55.705 1794.650 58.535 ;
        RECT 5.330 50.265 1794.650 53.095 ;
        RECT 5.330 44.825 1794.650 47.655 ;
        RECT 5.330 39.385 1794.650 42.215 ;
        RECT 5.330 33.945 1794.650 36.775 ;
        RECT 5.330 28.505 1794.650 31.335 ;
        RECT 5.330 23.065 1794.650 25.895 ;
        RECT 5.330 17.625 1794.650 20.455 ;
        RECT 5.330 12.185 1794.650 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 1794.460 3087.285 ;
      LAYER met1 ;
        RECT 5.520 10.640 1797.150 3087.440 ;
      LAYER met2 ;
        RECT 21.070 10.695 1797.120 3087.385 ;
      LAYER met3 ;
        RECT 21.050 3062.400 1796.235 3087.365 ;
        RECT 21.050 3061.000 1795.600 3062.400 ;
        RECT 21.050 3009.360 1796.235 3061.000 ;
        RECT 21.050 3007.960 1795.600 3009.360 ;
        RECT 21.050 2956.320 1796.235 3007.960 ;
        RECT 21.050 2954.920 1795.600 2956.320 ;
        RECT 21.050 2903.280 1796.235 2954.920 ;
        RECT 21.050 2901.880 1795.600 2903.280 ;
        RECT 21.050 2850.240 1796.235 2901.880 ;
        RECT 21.050 2848.840 1795.600 2850.240 ;
        RECT 21.050 2797.200 1796.235 2848.840 ;
        RECT 21.050 2795.800 1795.600 2797.200 ;
        RECT 21.050 2744.160 1796.235 2795.800 ;
        RECT 21.050 2742.760 1795.600 2744.160 ;
        RECT 21.050 2691.120 1796.235 2742.760 ;
        RECT 21.050 2689.720 1795.600 2691.120 ;
        RECT 21.050 2638.080 1796.235 2689.720 ;
        RECT 21.050 2636.680 1795.600 2638.080 ;
        RECT 21.050 2585.040 1796.235 2636.680 ;
        RECT 21.050 2583.640 1795.600 2585.040 ;
        RECT 21.050 2532.000 1796.235 2583.640 ;
        RECT 21.050 2530.600 1795.600 2532.000 ;
        RECT 21.050 2478.960 1796.235 2530.600 ;
        RECT 21.050 2477.560 1795.600 2478.960 ;
        RECT 21.050 2425.920 1796.235 2477.560 ;
        RECT 21.050 2424.520 1795.600 2425.920 ;
        RECT 21.050 2372.880 1796.235 2424.520 ;
        RECT 21.050 2371.480 1795.600 2372.880 ;
        RECT 21.050 2319.840 1796.235 2371.480 ;
        RECT 21.050 2318.440 1795.600 2319.840 ;
        RECT 21.050 2266.800 1796.235 2318.440 ;
        RECT 21.050 2265.400 1795.600 2266.800 ;
        RECT 21.050 2213.760 1796.235 2265.400 ;
        RECT 21.050 2212.360 1795.600 2213.760 ;
        RECT 21.050 2160.720 1796.235 2212.360 ;
        RECT 21.050 2159.320 1795.600 2160.720 ;
        RECT 21.050 2107.680 1796.235 2159.320 ;
        RECT 21.050 2106.280 1795.600 2107.680 ;
        RECT 21.050 2054.640 1796.235 2106.280 ;
        RECT 21.050 2053.240 1795.600 2054.640 ;
        RECT 21.050 2001.600 1796.235 2053.240 ;
        RECT 21.050 2000.200 1795.600 2001.600 ;
        RECT 21.050 1948.560 1796.235 2000.200 ;
        RECT 21.050 1947.160 1795.600 1948.560 ;
        RECT 21.050 1895.520 1796.235 1947.160 ;
        RECT 21.050 1894.120 1795.600 1895.520 ;
        RECT 21.050 1842.480 1796.235 1894.120 ;
        RECT 21.050 1841.080 1795.600 1842.480 ;
        RECT 21.050 1789.440 1796.235 1841.080 ;
        RECT 21.050 1788.040 1795.600 1789.440 ;
        RECT 21.050 1736.400 1796.235 1788.040 ;
        RECT 21.050 1735.000 1795.600 1736.400 ;
        RECT 21.050 1683.360 1796.235 1735.000 ;
        RECT 21.050 1681.960 1795.600 1683.360 ;
        RECT 21.050 1630.320 1796.235 1681.960 ;
        RECT 21.050 1628.920 1795.600 1630.320 ;
        RECT 21.050 1577.280 1796.235 1628.920 ;
        RECT 21.050 1575.880 1795.600 1577.280 ;
        RECT 21.050 1524.240 1796.235 1575.880 ;
        RECT 21.050 1522.840 1795.600 1524.240 ;
        RECT 21.050 1471.200 1796.235 1522.840 ;
        RECT 21.050 1469.800 1795.600 1471.200 ;
        RECT 21.050 1418.160 1796.235 1469.800 ;
        RECT 21.050 1416.760 1795.600 1418.160 ;
        RECT 21.050 1365.120 1796.235 1416.760 ;
        RECT 21.050 1363.720 1795.600 1365.120 ;
        RECT 21.050 1312.080 1796.235 1363.720 ;
        RECT 21.050 1310.680 1795.600 1312.080 ;
        RECT 21.050 1259.040 1796.235 1310.680 ;
        RECT 21.050 1257.640 1795.600 1259.040 ;
        RECT 21.050 1206.000 1796.235 1257.640 ;
        RECT 21.050 1204.600 1795.600 1206.000 ;
        RECT 21.050 1152.960 1796.235 1204.600 ;
        RECT 21.050 1151.560 1795.600 1152.960 ;
        RECT 21.050 1099.920 1796.235 1151.560 ;
        RECT 21.050 1098.520 1795.600 1099.920 ;
        RECT 21.050 1046.880 1796.235 1098.520 ;
        RECT 21.050 1045.480 1795.600 1046.880 ;
        RECT 21.050 993.840 1796.235 1045.480 ;
        RECT 21.050 992.440 1795.600 993.840 ;
        RECT 21.050 940.800 1796.235 992.440 ;
        RECT 21.050 939.400 1795.600 940.800 ;
        RECT 21.050 887.760 1796.235 939.400 ;
        RECT 21.050 886.360 1795.600 887.760 ;
        RECT 21.050 834.720 1796.235 886.360 ;
        RECT 21.050 833.320 1795.600 834.720 ;
        RECT 21.050 781.680 1796.235 833.320 ;
        RECT 21.050 780.280 1795.600 781.680 ;
        RECT 21.050 728.640 1796.235 780.280 ;
        RECT 21.050 727.240 1795.600 728.640 ;
        RECT 21.050 675.600 1796.235 727.240 ;
        RECT 21.050 674.200 1795.600 675.600 ;
        RECT 21.050 622.560 1796.235 674.200 ;
        RECT 21.050 621.160 1795.600 622.560 ;
        RECT 21.050 569.520 1796.235 621.160 ;
        RECT 21.050 568.120 1795.600 569.520 ;
        RECT 21.050 516.480 1796.235 568.120 ;
        RECT 21.050 515.080 1795.600 516.480 ;
        RECT 21.050 463.440 1796.235 515.080 ;
        RECT 21.050 462.040 1795.600 463.440 ;
        RECT 21.050 410.400 1796.235 462.040 ;
        RECT 21.050 409.000 1795.600 410.400 ;
        RECT 21.050 357.360 1796.235 409.000 ;
        RECT 21.050 355.960 1795.600 357.360 ;
        RECT 21.050 304.320 1796.235 355.960 ;
        RECT 21.050 302.920 1795.600 304.320 ;
        RECT 21.050 251.280 1796.235 302.920 ;
        RECT 21.050 249.880 1795.600 251.280 ;
        RECT 21.050 198.240 1796.235 249.880 ;
        RECT 21.050 196.840 1795.600 198.240 ;
        RECT 21.050 145.200 1796.235 196.840 ;
        RECT 21.050 143.800 1795.600 145.200 ;
        RECT 21.050 92.160 1796.235 143.800 ;
        RECT 21.050 90.760 1795.600 92.160 ;
        RECT 21.050 39.120 1796.235 90.760 ;
        RECT 21.050 37.720 1795.600 39.120 ;
        RECT 21.050 10.715 1796.235 37.720 ;
      LAYER met4 ;
        RECT 254.215 54.575 327.840 3074.785 ;
        RECT 330.240 54.575 404.640 3074.785 ;
        RECT 407.040 54.575 481.440 3074.785 ;
        RECT 483.840 54.575 558.240 3074.785 ;
        RECT 560.640 54.575 635.040 3074.785 ;
        RECT 637.440 54.575 711.840 3074.785 ;
        RECT 714.240 54.575 788.640 3074.785 ;
        RECT 791.040 54.575 865.440 3074.785 ;
        RECT 867.840 54.575 942.240 3074.785 ;
        RECT 944.640 54.575 1019.040 3074.785 ;
        RECT 1021.440 54.575 1095.840 3074.785 ;
        RECT 1098.240 54.575 1172.640 3074.785 ;
        RECT 1175.040 54.575 1249.440 3074.785 ;
        RECT 1251.840 54.575 1326.240 3074.785 ;
        RECT 1328.640 54.575 1403.040 3074.785 ;
        RECT 1405.440 54.575 1479.840 3074.785 ;
        RECT 1482.240 54.575 1556.640 3074.785 ;
        RECT 1559.040 54.575 1633.440 3074.785 ;
        RECT 1635.840 54.575 1710.240 3074.785 ;
        RECT 1712.640 54.575 1765.185 3074.785 ;
  END
END wrapped_as512512512
END LIBRARY

