magic
tech sky130B
magscale 1 2
timestamp 1680008680
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 934 76 59786 59152
<< metal2 >>
rect 2226 59200 2282 60000
rect 3514 59200 3570 60000
rect 4802 59200 4858 60000
rect 6090 59200 6146 60000
rect 7378 59200 7434 60000
rect 8666 59200 8722 60000
rect 9954 59200 10010 60000
rect 11242 59200 11298 60000
rect 12530 59200 12586 60000
rect 13818 59200 13874 60000
rect 15106 59200 15162 60000
rect 16394 59200 16450 60000
rect 17682 59200 17738 60000
rect 18970 59200 19026 60000
rect 20258 59200 20314 60000
rect 21546 59200 21602 60000
rect 22834 59200 22890 60000
rect 24122 59200 24178 60000
rect 25410 59200 25466 60000
rect 26698 59200 26754 60000
rect 27986 59200 28042 60000
rect 29274 59200 29330 60000
rect 30562 59200 30618 60000
rect 31850 59200 31906 60000
rect 33138 59200 33194 60000
rect 34426 59200 34482 60000
rect 35714 59200 35770 60000
rect 37002 59200 37058 60000
rect 38290 59200 38346 60000
rect 39578 59200 39634 60000
rect 40866 59200 40922 60000
rect 42154 59200 42210 60000
rect 43442 59200 43498 60000
rect 44730 59200 44786 60000
rect 46018 59200 46074 60000
rect 47306 59200 47362 60000
rect 48594 59200 48650 60000
rect 49882 59200 49938 60000
rect 51170 59200 51226 60000
rect 52458 59200 52514 60000
rect 53746 59200 53802 60000
rect 55034 59200 55090 60000
rect 56322 59200 56378 60000
rect 57610 59200 57666 60000
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 53930 0 53986 800
<< obsm2 >>
rect 938 59144 2170 59200
rect 2338 59144 3458 59200
rect 3626 59144 4746 59200
rect 4914 59144 6034 59200
rect 6202 59144 7322 59200
rect 7490 59144 8610 59200
rect 8778 59144 9898 59200
rect 10066 59144 11186 59200
rect 11354 59144 12474 59200
rect 12642 59144 13762 59200
rect 13930 59144 15050 59200
rect 15218 59144 16338 59200
rect 16506 59144 17626 59200
rect 17794 59144 18914 59200
rect 19082 59144 20202 59200
rect 20370 59144 21490 59200
rect 21658 59144 22778 59200
rect 22946 59144 24066 59200
rect 24234 59144 25354 59200
rect 25522 59144 26642 59200
rect 26810 59144 27930 59200
rect 28098 59144 29218 59200
rect 29386 59144 30506 59200
rect 30674 59144 31794 59200
rect 31962 59144 33082 59200
rect 33250 59144 34370 59200
rect 34538 59144 35658 59200
rect 35826 59144 36946 59200
rect 37114 59144 38234 59200
rect 38402 59144 39522 59200
rect 39690 59144 40810 59200
rect 40978 59144 42098 59200
rect 42266 59144 43386 59200
rect 43554 59144 44674 59200
rect 44842 59144 45962 59200
rect 46130 59144 47250 59200
rect 47418 59144 48538 59200
rect 48706 59144 49826 59200
rect 49994 59144 51114 59200
rect 51282 59144 52402 59200
rect 52570 59144 53690 59200
rect 53858 59144 54978 59200
rect 55146 59144 56266 59200
rect 56434 59144 57554 59200
rect 57722 59144 59780 59200
rect 938 856 59780 59144
rect 938 70 5850 856
rect 6018 70 6126 856
rect 6294 70 6402 856
rect 6570 70 6678 856
rect 6846 70 6954 856
rect 7122 70 7230 856
rect 7398 70 7506 856
rect 7674 70 7782 856
rect 7950 70 8058 856
rect 8226 70 8334 856
rect 8502 70 8610 856
rect 8778 70 8886 856
rect 9054 70 9162 856
rect 9330 70 9438 856
rect 9606 70 9714 856
rect 9882 70 9990 856
rect 10158 70 10266 856
rect 10434 70 10542 856
rect 10710 70 10818 856
rect 10986 70 11094 856
rect 11262 70 11370 856
rect 11538 70 11646 856
rect 11814 70 11922 856
rect 12090 70 12198 856
rect 12366 70 12474 856
rect 12642 70 12750 856
rect 12918 70 13026 856
rect 13194 70 13302 856
rect 13470 70 13578 856
rect 13746 70 13854 856
rect 14022 70 14130 856
rect 14298 70 14406 856
rect 14574 70 14682 856
rect 14850 70 14958 856
rect 15126 70 15234 856
rect 15402 70 15510 856
rect 15678 70 15786 856
rect 15954 70 16062 856
rect 16230 70 16338 856
rect 16506 70 16614 856
rect 16782 70 16890 856
rect 17058 70 17166 856
rect 17334 70 17442 856
rect 17610 70 17718 856
rect 17886 70 17994 856
rect 18162 70 18270 856
rect 18438 70 18546 856
rect 18714 70 18822 856
rect 18990 70 19098 856
rect 19266 70 19374 856
rect 19542 70 19650 856
rect 19818 70 19926 856
rect 20094 70 20202 856
rect 20370 70 20478 856
rect 20646 70 20754 856
rect 20922 70 21030 856
rect 21198 70 21306 856
rect 21474 70 21582 856
rect 21750 70 21858 856
rect 22026 70 22134 856
rect 22302 70 22410 856
rect 22578 70 22686 856
rect 22854 70 22962 856
rect 23130 70 23238 856
rect 23406 70 23514 856
rect 23682 70 23790 856
rect 23958 70 24066 856
rect 24234 70 24342 856
rect 24510 70 24618 856
rect 24786 70 24894 856
rect 25062 70 25170 856
rect 25338 70 25446 856
rect 25614 70 25722 856
rect 25890 70 25998 856
rect 26166 70 26274 856
rect 26442 70 26550 856
rect 26718 70 26826 856
rect 26994 70 27102 856
rect 27270 70 27378 856
rect 27546 70 27654 856
rect 27822 70 27930 856
rect 28098 70 28206 856
rect 28374 70 28482 856
rect 28650 70 28758 856
rect 28926 70 29034 856
rect 29202 70 29310 856
rect 29478 70 29586 856
rect 29754 70 29862 856
rect 30030 70 30138 856
rect 30306 70 30414 856
rect 30582 70 30690 856
rect 30858 70 30966 856
rect 31134 70 31242 856
rect 31410 70 31518 856
rect 31686 70 31794 856
rect 31962 70 32070 856
rect 32238 70 32346 856
rect 32514 70 32622 856
rect 32790 70 32898 856
rect 33066 70 33174 856
rect 33342 70 33450 856
rect 33618 70 33726 856
rect 33894 70 34002 856
rect 34170 70 34278 856
rect 34446 70 34554 856
rect 34722 70 34830 856
rect 34998 70 35106 856
rect 35274 70 35382 856
rect 35550 70 35658 856
rect 35826 70 35934 856
rect 36102 70 36210 856
rect 36378 70 36486 856
rect 36654 70 36762 856
rect 36930 70 37038 856
rect 37206 70 37314 856
rect 37482 70 37590 856
rect 37758 70 37866 856
rect 38034 70 38142 856
rect 38310 70 38418 856
rect 38586 70 38694 856
rect 38862 70 38970 856
rect 39138 70 39246 856
rect 39414 70 39522 856
rect 39690 70 39798 856
rect 39966 70 40074 856
rect 40242 70 40350 856
rect 40518 70 40626 856
rect 40794 70 40902 856
rect 41070 70 41178 856
rect 41346 70 41454 856
rect 41622 70 41730 856
rect 41898 70 42006 856
rect 42174 70 42282 856
rect 42450 70 42558 856
rect 42726 70 42834 856
rect 43002 70 43110 856
rect 43278 70 43386 856
rect 43554 70 43662 856
rect 43830 70 43938 856
rect 44106 70 44214 856
rect 44382 70 44490 856
rect 44658 70 44766 856
rect 44934 70 45042 856
rect 45210 70 45318 856
rect 45486 70 45594 856
rect 45762 70 45870 856
rect 46038 70 46146 856
rect 46314 70 46422 856
rect 46590 70 46698 856
rect 46866 70 46974 856
rect 47142 70 47250 856
rect 47418 70 47526 856
rect 47694 70 47802 856
rect 47970 70 48078 856
rect 48246 70 48354 856
rect 48522 70 48630 856
rect 48798 70 48906 856
rect 49074 70 49182 856
rect 49350 70 49458 856
rect 49626 70 49734 856
rect 49902 70 50010 856
rect 50178 70 50286 856
rect 50454 70 50562 856
rect 50730 70 50838 856
rect 51006 70 51114 856
rect 51282 70 51390 856
rect 51558 70 51666 856
rect 51834 70 51942 856
rect 52110 70 52218 856
rect 52386 70 52494 856
rect 52662 70 52770 856
rect 52938 70 53046 856
rect 53214 70 53322 856
rect 53490 70 53598 856
rect 53766 70 53874 856
rect 54042 70 59780 856
<< metal3 >>
rect 59200 58624 60000 58744
rect 59200 58216 60000 58336
rect 59200 57808 60000 57928
rect 59200 57400 60000 57520
rect 59200 56992 60000 57112
rect 59200 56584 60000 56704
rect 59200 56176 60000 56296
rect 0 55768 800 55888
rect 59200 55768 60000 55888
rect 0 55224 800 55344
rect 59200 55360 60000 55480
rect 59200 54952 60000 55072
rect 0 54680 800 54800
rect 59200 54544 60000 54664
rect 0 54136 800 54256
rect 59200 54136 60000 54256
rect 0 53592 800 53712
rect 59200 53728 60000 53848
rect 59200 53320 60000 53440
rect 0 53048 800 53168
rect 59200 52912 60000 53032
rect 0 52504 800 52624
rect 59200 52504 60000 52624
rect 0 51960 800 52080
rect 59200 52096 60000 52216
rect 59200 51688 60000 51808
rect 0 51416 800 51536
rect 59200 51280 60000 51400
rect 0 50872 800 50992
rect 59200 50872 60000 50992
rect 0 50328 800 50448
rect 59200 50464 60000 50584
rect 59200 50056 60000 50176
rect 0 49784 800 49904
rect 59200 49648 60000 49768
rect 0 49240 800 49360
rect 59200 49240 60000 49360
rect 0 48696 800 48816
rect 59200 48832 60000 48952
rect 59200 48424 60000 48544
rect 0 48152 800 48272
rect 59200 48016 60000 48136
rect 0 47608 800 47728
rect 59200 47608 60000 47728
rect 0 47064 800 47184
rect 59200 47200 60000 47320
rect 59200 46792 60000 46912
rect 0 46520 800 46640
rect 59200 46384 60000 46504
rect 0 45976 800 46096
rect 59200 45976 60000 46096
rect 0 45432 800 45552
rect 59200 45568 60000 45688
rect 59200 45160 60000 45280
rect 0 44888 800 45008
rect 59200 44752 60000 44872
rect 0 44344 800 44464
rect 59200 44344 60000 44464
rect 0 43800 800 43920
rect 59200 43936 60000 44056
rect 59200 43528 60000 43648
rect 0 43256 800 43376
rect 59200 43120 60000 43240
rect 0 42712 800 42832
rect 59200 42712 60000 42832
rect 0 42168 800 42288
rect 59200 42304 60000 42424
rect 59200 41896 60000 42016
rect 0 41624 800 41744
rect 59200 41488 60000 41608
rect 0 41080 800 41200
rect 59200 41080 60000 41200
rect 0 40536 800 40656
rect 59200 40672 60000 40792
rect 59200 40264 60000 40384
rect 0 39992 800 40112
rect 59200 39856 60000 39976
rect 0 39448 800 39568
rect 59200 39448 60000 39568
rect 0 38904 800 39024
rect 59200 39040 60000 39160
rect 59200 38632 60000 38752
rect 0 38360 800 38480
rect 59200 38224 60000 38344
rect 0 37816 800 37936
rect 59200 37816 60000 37936
rect 0 37272 800 37392
rect 59200 37408 60000 37528
rect 59200 37000 60000 37120
rect 0 36728 800 36848
rect 59200 36592 60000 36712
rect 0 36184 800 36304
rect 59200 36184 60000 36304
rect 0 35640 800 35760
rect 59200 35776 60000 35896
rect 59200 35368 60000 35488
rect 0 35096 800 35216
rect 59200 34960 60000 35080
rect 0 34552 800 34672
rect 59200 34552 60000 34672
rect 0 34008 800 34128
rect 59200 34144 60000 34264
rect 59200 33736 60000 33856
rect 0 33464 800 33584
rect 59200 33328 60000 33448
rect 0 32920 800 33040
rect 59200 32920 60000 33040
rect 0 32376 800 32496
rect 59200 32512 60000 32632
rect 59200 32104 60000 32224
rect 0 31832 800 31952
rect 59200 31696 60000 31816
rect 0 31288 800 31408
rect 59200 31288 60000 31408
rect 0 30744 800 30864
rect 59200 30880 60000 31000
rect 59200 30472 60000 30592
rect 0 30200 800 30320
rect 59200 30064 60000 30184
rect 0 29656 800 29776
rect 59200 29656 60000 29776
rect 0 29112 800 29232
rect 59200 29248 60000 29368
rect 59200 28840 60000 28960
rect 0 28568 800 28688
rect 59200 28432 60000 28552
rect 0 28024 800 28144
rect 59200 28024 60000 28144
rect 0 27480 800 27600
rect 59200 27616 60000 27736
rect 59200 27208 60000 27328
rect 0 26936 800 27056
rect 59200 26800 60000 26920
rect 0 26392 800 26512
rect 59200 26392 60000 26512
rect 0 25848 800 25968
rect 59200 25984 60000 26104
rect 59200 25576 60000 25696
rect 0 25304 800 25424
rect 59200 25168 60000 25288
rect 0 24760 800 24880
rect 59200 24760 60000 24880
rect 0 24216 800 24336
rect 59200 24352 60000 24472
rect 59200 23944 60000 24064
rect 0 23672 800 23792
rect 59200 23536 60000 23656
rect 0 23128 800 23248
rect 59200 23128 60000 23248
rect 0 22584 800 22704
rect 59200 22720 60000 22840
rect 59200 22312 60000 22432
rect 0 22040 800 22160
rect 59200 21904 60000 22024
rect 0 21496 800 21616
rect 59200 21496 60000 21616
rect 0 20952 800 21072
rect 59200 21088 60000 21208
rect 59200 20680 60000 20800
rect 0 20408 800 20528
rect 59200 20272 60000 20392
rect 0 19864 800 19984
rect 59200 19864 60000 19984
rect 0 19320 800 19440
rect 59200 19456 60000 19576
rect 59200 19048 60000 19168
rect 0 18776 800 18896
rect 59200 18640 60000 18760
rect 0 18232 800 18352
rect 59200 18232 60000 18352
rect 0 17688 800 17808
rect 59200 17824 60000 17944
rect 59200 17416 60000 17536
rect 0 17144 800 17264
rect 59200 17008 60000 17128
rect 0 16600 800 16720
rect 59200 16600 60000 16720
rect 0 16056 800 16176
rect 59200 16192 60000 16312
rect 59200 15784 60000 15904
rect 0 15512 800 15632
rect 59200 15376 60000 15496
rect 0 14968 800 15088
rect 59200 14968 60000 15088
rect 0 14424 800 14544
rect 59200 14560 60000 14680
rect 59200 14152 60000 14272
rect 0 13880 800 14000
rect 59200 13744 60000 13864
rect 0 13336 800 13456
rect 59200 13336 60000 13456
rect 0 12792 800 12912
rect 59200 12928 60000 13048
rect 59200 12520 60000 12640
rect 0 12248 800 12368
rect 59200 12112 60000 12232
rect 0 11704 800 11824
rect 59200 11704 60000 11824
rect 0 11160 800 11280
rect 59200 11296 60000 11416
rect 59200 10888 60000 11008
rect 0 10616 800 10736
rect 59200 10480 60000 10600
rect 0 10072 800 10192
rect 59200 10072 60000 10192
rect 0 9528 800 9648
rect 59200 9664 60000 9784
rect 59200 9256 60000 9376
rect 0 8984 800 9104
rect 59200 8848 60000 8968
rect 0 8440 800 8560
rect 59200 8440 60000 8560
rect 0 7896 800 8016
rect 59200 8032 60000 8152
rect 59200 7624 60000 7744
rect 0 7352 800 7472
rect 59200 7216 60000 7336
rect 0 6808 800 6928
rect 59200 6808 60000 6928
rect 0 6264 800 6384
rect 59200 6400 60000 6520
rect 59200 5992 60000 6112
rect 0 5720 800 5840
rect 59200 5584 60000 5704
rect 0 5176 800 5296
rect 59200 5176 60000 5296
rect 0 4632 800 4752
rect 59200 4768 60000 4888
rect 59200 4360 60000 4480
rect 0 4088 800 4208
rect 59200 3952 60000 4072
rect 59200 3544 60000 3664
rect 59200 3136 60000 3256
rect 59200 2728 60000 2848
rect 59200 2320 60000 2440
rect 59200 1912 60000 2032
rect 59200 1504 60000 1624
rect 59200 1096 60000 1216
<< obsm3 >>
rect 800 58544 59120 58717
rect 800 58416 59200 58544
rect 800 58136 59120 58416
rect 800 58008 59200 58136
rect 800 57728 59120 58008
rect 800 57600 59200 57728
rect 800 57320 59120 57600
rect 800 57192 59200 57320
rect 800 56912 59120 57192
rect 800 56784 59200 56912
rect 800 56504 59120 56784
rect 800 56376 59200 56504
rect 800 56096 59120 56376
rect 800 55968 59200 56096
rect 880 55688 59120 55968
rect 800 55560 59200 55688
rect 800 55424 59120 55560
rect 880 55280 59120 55424
rect 880 55152 59200 55280
rect 880 55144 59120 55152
rect 800 54880 59120 55144
rect 880 54872 59120 54880
rect 880 54744 59200 54872
rect 880 54600 59120 54744
rect 800 54464 59120 54600
rect 800 54336 59200 54464
rect 880 54056 59120 54336
rect 800 53928 59200 54056
rect 800 53792 59120 53928
rect 880 53648 59120 53792
rect 880 53520 59200 53648
rect 880 53512 59120 53520
rect 800 53248 59120 53512
rect 880 53240 59120 53248
rect 880 53112 59200 53240
rect 880 52968 59120 53112
rect 800 52832 59120 52968
rect 800 52704 59200 52832
rect 880 52424 59120 52704
rect 800 52296 59200 52424
rect 800 52160 59120 52296
rect 880 52016 59120 52160
rect 880 51888 59200 52016
rect 880 51880 59120 51888
rect 800 51616 59120 51880
rect 880 51608 59120 51616
rect 880 51480 59200 51608
rect 880 51336 59120 51480
rect 800 51200 59120 51336
rect 800 51072 59200 51200
rect 880 50792 59120 51072
rect 800 50664 59200 50792
rect 800 50528 59120 50664
rect 880 50384 59120 50528
rect 880 50256 59200 50384
rect 880 50248 59120 50256
rect 800 49984 59120 50248
rect 880 49976 59120 49984
rect 880 49848 59200 49976
rect 880 49704 59120 49848
rect 800 49568 59120 49704
rect 800 49440 59200 49568
rect 880 49160 59120 49440
rect 800 49032 59200 49160
rect 800 48896 59120 49032
rect 880 48752 59120 48896
rect 880 48624 59200 48752
rect 880 48616 59120 48624
rect 800 48352 59120 48616
rect 880 48344 59120 48352
rect 880 48216 59200 48344
rect 880 48072 59120 48216
rect 800 47936 59120 48072
rect 800 47808 59200 47936
rect 880 47528 59120 47808
rect 800 47400 59200 47528
rect 800 47264 59120 47400
rect 880 47120 59120 47264
rect 880 46992 59200 47120
rect 880 46984 59120 46992
rect 800 46720 59120 46984
rect 880 46712 59120 46720
rect 880 46584 59200 46712
rect 880 46440 59120 46584
rect 800 46304 59120 46440
rect 800 46176 59200 46304
rect 880 45896 59120 46176
rect 800 45768 59200 45896
rect 800 45632 59120 45768
rect 880 45488 59120 45632
rect 880 45360 59200 45488
rect 880 45352 59120 45360
rect 800 45088 59120 45352
rect 880 45080 59120 45088
rect 880 44952 59200 45080
rect 880 44808 59120 44952
rect 800 44672 59120 44808
rect 800 44544 59200 44672
rect 880 44264 59120 44544
rect 800 44136 59200 44264
rect 800 44000 59120 44136
rect 880 43856 59120 44000
rect 880 43728 59200 43856
rect 880 43720 59120 43728
rect 800 43456 59120 43720
rect 880 43448 59120 43456
rect 880 43320 59200 43448
rect 880 43176 59120 43320
rect 800 43040 59120 43176
rect 800 42912 59200 43040
rect 880 42632 59120 42912
rect 800 42504 59200 42632
rect 800 42368 59120 42504
rect 880 42224 59120 42368
rect 880 42096 59200 42224
rect 880 42088 59120 42096
rect 800 41824 59120 42088
rect 880 41816 59120 41824
rect 880 41688 59200 41816
rect 880 41544 59120 41688
rect 800 41408 59120 41544
rect 800 41280 59200 41408
rect 880 41000 59120 41280
rect 800 40872 59200 41000
rect 800 40736 59120 40872
rect 880 40592 59120 40736
rect 880 40464 59200 40592
rect 880 40456 59120 40464
rect 800 40192 59120 40456
rect 880 40184 59120 40192
rect 880 40056 59200 40184
rect 880 39912 59120 40056
rect 800 39776 59120 39912
rect 800 39648 59200 39776
rect 880 39368 59120 39648
rect 800 39240 59200 39368
rect 800 39104 59120 39240
rect 880 38960 59120 39104
rect 880 38832 59200 38960
rect 880 38824 59120 38832
rect 800 38560 59120 38824
rect 880 38552 59120 38560
rect 880 38424 59200 38552
rect 880 38280 59120 38424
rect 800 38144 59120 38280
rect 800 38016 59200 38144
rect 880 37736 59120 38016
rect 800 37608 59200 37736
rect 800 37472 59120 37608
rect 880 37328 59120 37472
rect 880 37200 59200 37328
rect 880 37192 59120 37200
rect 800 36928 59120 37192
rect 880 36920 59120 36928
rect 880 36792 59200 36920
rect 880 36648 59120 36792
rect 800 36512 59120 36648
rect 800 36384 59200 36512
rect 880 36104 59120 36384
rect 800 35976 59200 36104
rect 800 35840 59120 35976
rect 880 35696 59120 35840
rect 880 35568 59200 35696
rect 880 35560 59120 35568
rect 800 35296 59120 35560
rect 880 35288 59120 35296
rect 880 35160 59200 35288
rect 880 35016 59120 35160
rect 800 34880 59120 35016
rect 800 34752 59200 34880
rect 880 34472 59120 34752
rect 800 34344 59200 34472
rect 800 34208 59120 34344
rect 880 34064 59120 34208
rect 880 33936 59200 34064
rect 880 33928 59120 33936
rect 800 33664 59120 33928
rect 880 33656 59120 33664
rect 880 33528 59200 33656
rect 880 33384 59120 33528
rect 800 33248 59120 33384
rect 800 33120 59200 33248
rect 880 32840 59120 33120
rect 800 32712 59200 32840
rect 800 32576 59120 32712
rect 880 32432 59120 32576
rect 880 32304 59200 32432
rect 880 32296 59120 32304
rect 800 32032 59120 32296
rect 880 32024 59120 32032
rect 880 31896 59200 32024
rect 880 31752 59120 31896
rect 800 31616 59120 31752
rect 800 31488 59200 31616
rect 880 31208 59120 31488
rect 800 31080 59200 31208
rect 800 30944 59120 31080
rect 880 30800 59120 30944
rect 880 30672 59200 30800
rect 880 30664 59120 30672
rect 800 30400 59120 30664
rect 880 30392 59120 30400
rect 880 30264 59200 30392
rect 880 30120 59120 30264
rect 800 29984 59120 30120
rect 800 29856 59200 29984
rect 880 29576 59120 29856
rect 800 29448 59200 29576
rect 800 29312 59120 29448
rect 880 29168 59120 29312
rect 880 29040 59200 29168
rect 880 29032 59120 29040
rect 800 28768 59120 29032
rect 880 28760 59120 28768
rect 880 28632 59200 28760
rect 880 28488 59120 28632
rect 800 28352 59120 28488
rect 800 28224 59200 28352
rect 880 27944 59120 28224
rect 800 27816 59200 27944
rect 800 27680 59120 27816
rect 880 27536 59120 27680
rect 880 27408 59200 27536
rect 880 27400 59120 27408
rect 800 27136 59120 27400
rect 880 27128 59120 27136
rect 880 27000 59200 27128
rect 880 26856 59120 27000
rect 800 26720 59120 26856
rect 800 26592 59200 26720
rect 880 26312 59120 26592
rect 800 26184 59200 26312
rect 800 26048 59120 26184
rect 880 25904 59120 26048
rect 880 25776 59200 25904
rect 880 25768 59120 25776
rect 800 25504 59120 25768
rect 880 25496 59120 25504
rect 880 25368 59200 25496
rect 880 25224 59120 25368
rect 800 25088 59120 25224
rect 800 24960 59200 25088
rect 880 24680 59120 24960
rect 800 24552 59200 24680
rect 800 24416 59120 24552
rect 880 24272 59120 24416
rect 880 24144 59200 24272
rect 880 24136 59120 24144
rect 800 23872 59120 24136
rect 880 23864 59120 23872
rect 880 23736 59200 23864
rect 880 23592 59120 23736
rect 800 23456 59120 23592
rect 800 23328 59200 23456
rect 880 23048 59120 23328
rect 800 22920 59200 23048
rect 800 22784 59120 22920
rect 880 22640 59120 22784
rect 880 22512 59200 22640
rect 880 22504 59120 22512
rect 800 22240 59120 22504
rect 880 22232 59120 22240
rect 880 22104 59200 22232
rect 880 21960 59120 22104
rect 800 21824 59120 21960
rect 800 21696 59200 21824
rect 880 21416 59120 21696
rect 800 21288 59200 21416
rect 800 21152 59120 21288
rect 880 21008 59120 21152
rect 880 20880 59200 21008
rect 880 20872 59120 20880
rect 800 20608 59120 20872
rect 880 20600 59120 20608
rect 880 20472 59200 20600
rect 880 20328 59120 20472
rect 800 20192 59120 20328
rect 800 20064 59200 20192
rect 880 19784 59120 20064
rect 800 19656 59200 19784
rect 800 19520 59120 19656
rect 880 19376 59120 19520
rect 880 19248 59200 19376
rect 880 19240 59120 19248
rect 800 18976 59120 19240
rect 880 18968 59120 18976
rect 880 18840 59200 18968
rect 880 18696 59120 18840
rect 800 18560 59120 18696
rect 800 18432 59200 18560
rect 880 18152 59120 18432
rect 800 18024 59200 18152
rect 800 17888 59120 18024
rect 880 17744 59120 17888
rect 880 17616 59200 17744
rect 880 17608 59120 17616
rect 800 17344 59120 17608
rect 880 17336 59120 17344
rect 880 17208 59200 17336
rect 880 17064 59120 17208
rect 800 16928 59120 17064
rect 800 16800 59200 16928
rect 880 16520 59120 16800
rect 800 16392 59200 16520
rect 800 16256 59120 16392
rect 880 16112 59120 16256
rect 880 15984 59200 16112
rect 880 15976 59120 15984
rect 800 15712 59120 15976
rect 880 15704 59120 15712
rect 880 15576 59200 15704
rect 880 15432 59120 15576
rect 800 15296 59120 15432
rect 800 15168 59200 15296
rect 880 14888 59120 15168
rect 800 14760 59200 14888
rect 800 14624 59120 14760
rect 880 14480 59120 14624
rect 880 14352 59200 14480
rect 880 14344 59120 14352
rect 800 14080 59120 14344
rect 880 14072 59120 14080
rect 880 13944 59200 14072
rect 880 13800 59120 13944
rect 800 13664 59120 13800
rect 800 13536 59200 13664
rect 880 13256 59120 13536
rect 800 13128 59200 13256
rect 800 12992 59120 13128
rect 880 12848 59120 12992
rect 880 12720 59200 12848
rect 880 12712 59120 12720
rect 800 12448 59120 12712
rect 880 12440 59120 12448
rect 880 12312 59200 12440
rect 880 12168 59120 12312
rect 800 12032 59120 12168
rect 800 11904 59200 12032
rect 880 11624 59120 11904
rect 800 11496 59200 11624
rect 800 11360 59120 11496
rect 880 11216 59120 11360
rect 880 11088 59200 11216
rect 880 11080 59120 11088
rect 800 10816 59120 11080
rect 880 10808 59120 10816
rect 880 10680 59200 10808
rect 880 10536 59120 10680
rect 800 10400 59120 10536
rect 800 10272 59200 10400
rect 880 9992 59120 10272
rect 800 9864 59200 9992
rect 800 9728 59120 9864
rect 880 9584 59120 9728
rect 880 9456 59200 9584
rect 880 9448 59120 9456
rect 800 9184 59120 9448
rect 880 9176 59120 9184
rect 880 9048 59200 9176
rect 880 8904 59120 9048
rect 800 8768 59120 8904
rect 800 8640 59200 8768
rect 880 8360 59120 8640
rect 800 8232 59200 8360
rect 800 8096 59120 8232
rect 880 7952 59120 8096
rect 880 7824 59200 7952
rect 880 7816 59120 7824
rect 800 7552 59120 7816
rect 880 7544 59120 7552
rect 880 7416 59200 7544
rect 880 7272 59120 7416
rect 800 7136 59120 7272
rect 800 7008 59200 7136
rect 880 6728 59120 7008
rect 800 6600 59200 6728
rect 800 6464 59120 6600
rect 880 6320 59120 6464
rect 880 6192 59200 6320
rect 880 6184 59120 6192
rect 800 5920 59120 6184
rect 880 5912 59120 5920
rect 880 5784 59200 5912
rect 880 5640 59120 5784
rect 800 5504 59120 5640
rect 800 5376 59200 5504
rect 880 5096 59120 5376
rect 800 4968 59200 5096
rect 800 4832 59120 4968
rect 880 4688 59120 4832
rect 880 4560 59200 4688
rect 880 4552 59120 4560
rect 800 4288 59120 4552
rect 880 4280 59120 4288
rect 880 4152 59200 4280
rect 880 4008 59120 4152
rect 800 3872 59120 4008
rect 800 3744 59200 3872
rect 800 3464 59120 3744
rect 800 3336 59200 3464
rect 800 3056 59120 3336
rect 800 2928 59200 3056
rect 800 2648 59120 2928
rect 800 2520 59200 2648
rect 800 2240 59120 2520
rect 800 2112 59200 2240
rect 800 1832 59120 2112
rect 800 1704 59200 1832
rect 800 1424 59120 1704
rect 800 1296 59200 1424
rect 800 1123 59120 1296
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< obsm4 >>
rect 29499 2347 34848 56677
rect 35328 2347 48885 56677
<< labels >>
rlabel metal3 s 0 19320 800 19440 6 design_clk_o
port 1 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 dsi_all[0]
port 2 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 dsi_all[10]
port 3 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 dsi_all[11]
port 4 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 dsi_all[12]
port 5 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 dsi_all[13]
port 6 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 dsi_all[14]
port 7 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 dsi_all[15]
port 8 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 dsi_all[16]
port 9 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 dsi_all[17]
port 10 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 dsi_all[18]
port 11 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 dsi_all[19]
port 12 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 dsi_all[1]
port 13 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 dsi_all[20]
port 14 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 dsi_all[21]
port 15 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 dsi_all[22]
port 16 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 dsi_all[23]
port 17 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 dsi_all[24]
port 18 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 dsi_all[25]
port 19 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 dsi_all[26]
port 20 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 dsi_all[27]
port 21 nsew signal output
rlabel metal3 s 0 5176 800 5296 6 dsi_all[2]
port 22 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 dsi_all[3]
port 23 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 dsi_all[4]
port 24 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 dsi_all[5]
port 25 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 dsi_all[6]
port 26 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 dsi_all[7]
port 27 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 dsi_all[8]
port 28 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 dsi_all[9]
port 29 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 dso_6502[0]
port 30 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 dso_6502[10]
port 31 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 dso_6502[11]
port 32 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 dso_6502[12]
port 33 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 dso_6502[13]
port 34 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 dso_6502[14]
port 35 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 dso_6502[15]
port 36 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 dso_6502[16]
port 37 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 dso_6502[17]
port 38 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 dso_6502[18]
port 39 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 dso_6502[19]
port 40 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 dso_6502[1]
port 41 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 dso_6502[20]
port 42 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 dso_6502[21]
port 43 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 dso_6502[22]
port 44 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 dso_6502[23]
port 45 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 dso_6502[24]
port 46 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 dso_6502[25]
port 47 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 dso_6502[26]
port 48 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 dso_6502[2]
port 49 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 dso_6502[3]
port 50 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 dso_6502[4]
port 51 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 dso_6502[5]
port 52 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 dso_6502[6]
port 53 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 dso_6502[7]
port 54 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 dso_6502[8]
port 55 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 dso_6502[9]
port 56 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 dso_LCD[0]
port 57 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 dso_LCD[1]
port 58 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 dso_LCD[2]
port 59 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 dso_LCD[3]
port 60 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 dso_LCD[4]
port 61 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 dso_LCD[5]
port 62 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 dso_LCD[6]
port 63 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 dso_LCD[7]
port 64 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 dso_as1802[0]
port 65 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 dso_as1802[10]
port 66 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 dso_as1802[11]
port 67 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 dso_as1802[12]
port 68 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 dso_as1802[13]
port 69 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 dso_as1802[14]
port 70 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 dso_as1802[15]
port 71 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 dso_as1802[16]
port 72 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 dso_as1802[17]
port 73 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 dso_as1802[18]
port 74 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 dso_as1802[19]
port 75 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 dso_as1802[1]
port 76 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 dso_as1802[20]
port 77 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 dso_as1802[21]
port 78 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 dso_as1802[22]
port 79 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 dso_as1802[23]
port 80 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 dso_as1802[24]
port 81 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 dso_as1802[25]
port 82 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 dso_as1802[26]
port 83 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 dso_as1802[2]
port 84 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 dso_as1802[3]
port 85 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 dso_as1802[4]
port 86 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 dso_as1802[5]
port 87 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 dso_as1802[6]
port 88 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 dso_as1802[7]
port 89 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 dso_as1802[8]
port 90 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 dso_as1802[9]
port 91 nsew signal input
rlabel metal2 s 24122 59200 24178 60000 6 dso_as2650[0]
port 92 nsew signal input
rlabel metal2 s 37002 59200 37058 60000 6 dso_as2650[10]
port 93 nsew signal input
rlabel metal2 s 38290 59200 38346 60000 6 dso_as2650[11]
port 94 nsew signal input
rlabel metal2 s 39578 59200 39634 60000 6 dso_as2650[12]
port 95 nsew signal input
rlabel metal2 s 40866 59200 40922 60000 6 dso_as2650[13]
port 96 nsew signal input
rlabel metal2 s 42154 59200 42210 60000 6 dso_as2650[14]
port 97 nsew signal input
rlabel metal2 s 43442 59200 43498 60000 6 dso_as2650[15]
port 98 nsew signal input
rlabel metal2 s 44730 59200 44786 60000 6 dso_as2650[16]
port 99 nsew signal input
rlabel metal2 s 46018 59200 46074 60000 6 dso_as2650[17]
port 100 nsew signal input
rlabel metal2 s 47306 59200 47362 60000 6 dso_as2650[18]
port 101 nsew signal input
rlabel metal2 s 48594 59200 48650 60000 6 dso_as2650[19]
port 102 nsew signal input
rlabel metal2 s 25410 59200 25466 60000 6 dso_as2650[1]
port 103 nsew signal input
rlabel metal2 s 49882 59200 49938 60000 6 dso_as2650[20]
port 104 nsew signal input
rlabel metal2 s 51170 59200 51226 60000 6 dso_as2650[21]
port 105 nsew signal input
rlabel metal2 s 52458 59200 52514 60000 6 dso_as2650[22]
port 106 nsew signal input
rlabel metal2 s 53746 59200 53802 60000 6 dso_as2650[23]
port 107 nsew signal input
rlabel metal2 s 55034 59200 55090 60000 6 dso_as2650[24]
port 108 nsew signal input
rlabel metal2 s 56322 59200 56378 60000 6 dso_as2650[25]
port 109 nsew signal input
rlabel metal2 s 57610 59200 57666 60000 6 dso_as2650[26]
port 110 nsew signal input
rlabel metal2 s 26698 59200 26754 60000 6 dso_as2650[2]
port 111 nsew signal input
rlabel metal2 s 27986 59200 28042 60000 6 dso_as2650[3]
port 112 nsew signal input
rlabel metal2 s 29274 59200 29330 60000 6 dso_as2650[4]
port 113 nsew signal input
rlabel metal2 s 30562 59200 30618 60000 6 dso_as2650[5]
port 114 nsew signal input
rlabel metal2 s 31850 59200 31906 60000 6 dso_as2650[6]
port 115 nsew signal input
rlabel metal2 s 33138 59200 33194 60000 6 dso_as2650[7]
port 116 nsew signal input
rlabel metal2 s 34426 59200 34482 60000 6 dso_as2650[8]
port 117 nsew signal input
rlabel metal2 s 35714 59200 35770 60000 6 dso_as2650[9]
port 118 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 dso_as512512512[0]
port 119 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 dso_as512512512[10]
port 120 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 dso_as512512512[11]
port 121 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 dso_as512512512[12]
port 122 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 dso_as512512512[13]
port 123 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 dso_as512512512[14]
port 124 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 dso_as512512512[15]
port 125 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 dso_as512512512[16]
port 126 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 dso_as512512512[17]
port 127 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 dso_as512512512[18]
port 128 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 dso_as512512512[19]
port 129 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 dso_as512512512[1]
port 130 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 dso_as512512512[20]
port 131 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 dso_as512512512[21]
port 132 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 dso_as512512512[22]
port 133 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 dso_as512512512[23]
port 134 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 dso_as512512512[24]
port 135 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 dso_as512512512[25]
port 136 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 dso_as512512512[26]
port 137 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 dso_as512512512[27]
port 138 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 dso_as512512512[2]
port 139 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 dso_as512512512[3]
port 140 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 dso_as512512512[4]
port 141 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 dso_as512512512[5]
port 142 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 dso_as512512512[6]
port 143 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 dso_as512512512[7]
port 144 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 dso_as512512512[8]
port 145 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 dso_as512512512[9]
port 146 nsew signal input
rlabel metal3 s 59200 47608 60000 47728 6 dso_as5401[0]
port 147 nsew signal input
rlabel metal3 s 59200 51688 60000 51808 6 dso_as5401[10]
port 148 nsew signal input
rlabel metal3 s 59200 52096 60000 52216 6 dso_as5401[11]
port 149 nsew signal input
rlabel metal3 s 59200 52504 60000 52624 6 dso_as5401[12]
port 150 nsew signal input
rlabel metal3 s 59200 52912 60000 53032 6 dso_as5401[13]
port 151 nsew signal input
rlabel metal3 s 59200 53320 60000 53440 6 dso_as5401[14]
port 152 nsew signal input
rlabel metal3 s 59200 53728 60000 53848 6 dso_as5401[15]
port 153 nsew signal input
rlabel metal3 s 59200 54136 60000 54256 6 dso_as5401[16]
port 154 nsew signal input
rlabel metal3 s 59200 54544 60000 54664 6 dso_as5401[17]
port 155 nsew signal input
rlabel metal3 s 59200 54952 60000 55072 6 dso_as5401[18]
port 156 nsew signal input
rlabel metal3 s 59200 55360 60000 55480 6 dso_as5401[19]
port 157 nsew signal input
rlabel metal3 s 59200 48016 60000 48136 6 dso_as5401[1]
port 158 nsew signal input
rlabel metal3 s 59200 55768 60000 55888 6 dso_as5401[20]
port 159 nsew signal input
rlabel metal3 s 59200 56176 60000 56296 6 dso_as5401[21]
port 160 nsew signal input
rlabel metal3 s 59200 56584 60000 56704 6 dso_as5401[22]
port 161 nsew signal input
rlabel metal3 s 59200 56992 60000 57112 6 dso_as5401[23]
port 162 nsew signal input
rlabel metal3 s 59200 57400 60000 57520 6 dso_as5401[24]
port 163 nsew signal input
rlabel metal3 s 59200 57808 60000 57928 6 dso_as5401[25]
port 164 nsew signal input
rlabel metal3 s 59200 58216 60000 58336 6 dso_as5401[26]
port 165 nsew signal input
rlabel metal3 s 59200 48424 60000 48544 6 dso_as5401[2]
port 166 nsew signal input
rlabel metal3 s 59200 48832 60000 48952 6 dso_as5401[3]
port 167 nsew signal input
rlabel metal3 s 59200 49240 60000 49360 6 dso_as5401[4]
port 168 nsew signal input
rlabel metal3 s 59200 49648 60000 49768 6 dso_as5401[5]
port 169 nsew signal input
rlabel metal3 s 59200 50056 60000 50176 6 dso_as5401[6]
port 170 nsew signal input
rlabel metal3 s 59200 50464 60000 50584 6 dso_as5401[7]
port 171 nsew signal input
rlabel metal3 s 59200 50872 60000 50992 6 dso_as5401[8]
port 172 nsew signal input
rlabel metal3 s 59200 51280 60000 51400 6 dso_as5401[9]
port 173 nsew signal input
rlabel metal3 s 59200 42712 60000 42832 6 dso_counter[0]
port 174 nsew signal input
rlabel metal3 s 59200 46792 60000 46912 6 dso_counter[10]
port 175 nsew signal input
rlabel metal3 s 59200 47200 60000 47320 6 dso_counter[11]
port 176 nsew signal input
rlabel metal3 s 59200 43120 60000 43240 6 dso_counter[1]
port 177 nsew signal input
rlabel metal3 s 59200 43528 60000 43648 6 dso_counter[2]
port 178 nsew signal input
rlabel metal3 s 59200 43936 60000 44056 6 dso_counter[3]
port 179 nsew signal input
rlabel metal3 s 59200 44344 60000 44464 6 dso_counter[4]
port 180 nsew signal input
rlabel metal3 s 59200 44752 60000 44872 6 dso_counter[5]
port 181 nsew signal input
rlabel metal3 s 59200 45160 60000 45280 6 dso_counter[6]
port 182 nsew signal input
rlabel metal3 s 59200 45568 60000 45688 6 dso_counter[7]
port 183 nsew signal input
rlabel metal3 s 59200 45976 60000 46096 6 dso_counter[8]
port 184 nsew signal input
rlabel metal3 s 59200 46384 60000 46504 6 dso_counter[9]
port 185 nsew signal input
rlabel metal2 s 12530 59200 12586 60000 6 dso_diceroll[0]
port 186 nsew signal input
rlabel metal2 s 13818 59200 13874 60000 6 dso_diceroll[1]
port 187 nsew signal input
rlabel metal2 s 15106 59200 15162 60000 6 dso_diceroll[2]
port 188 nsew signal input
rlabel metal2 s 16394 59200 16450 60000 6 dso_diceroll[3]
port 189 nsew signal input
rlabel metal2 s 17682 59200 17738 60000 6 dso_diceroll[4]
port 190 nsew signal input
rlabel metal2 s 18970 59200 19026 60000 6 dso_diceroll[5]
port 191 nsew signal input
rlabel metal2 s 20258 59200 20314 60000 6 dso_diceroll[6]
port 192 nsew signal input
rlabel metal2 s 21546 59200 21602 60000 6 dso_diceroll[7]
port 193 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 dso_mc14500[0]
port 194 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 dso_mc14500[1]
port 195 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 dso_mc14500[2]
port 196 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 dso_mc14500[3]
port 197 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 dso_mc14500[4]
port 198 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 dso_mc14500[5]
port 199 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 dso_mc14500[6]
port 200 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 dso_mc14500[7]
port 201 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 dso_mc14500[8]
port 202 nsew signal input
rlabel metal2 s 2226 59200 2282 60000 6 dso_multiplier[0]
port 203 nsew signal input
rlabel metal2 s 3514 59200 3570 60000 6 dso_multiplier[1]
port 204 nsew signal input
rlabel metal2 s 4802 59200 4858 60000 6 dso_multiplier[2]
port 205 nsew signal input
rlabel metal2 s 6090 59200 6146 60000 6 dso_multiplier[3]
port 206 nsew signal input
rlabel metal2 s 7378 59200 7434 60000 6 dso_multiplier[4]
port 207 nsew signal input
rlabel metal2 s 8666 59200 8722 60000 6 dso_multiplier[5]
port 208 nsew signal input
rlabel metal2 s 9954 59200 10010 60000 6 dso_multiplier[6]
port 209 nsew signal input
rlabel metal2 s 11242 59200 11298 60000 6 dso_multiplier[7]
port 210 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 dso_posit[0]
port 211 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 dso_posit[1]
port 212 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 dso_posit[2]
port 213 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 dso_posit[3]
port 214 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 dso_tbb1143[0]
port 215 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 dso_tbb1143[1]
port 216 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 dso_tbb1143[2]
port 217 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 dso_tbb1143[3]
port 218 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 dso_tbb1143[4]
port 219 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 dso_tbb1143[5]
port 220 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 dso_tbb1143[6]
port 221 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 dso_tbb1143[7]
port 222 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 dso_tune
port 223 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 io_in[0]
port 224 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 io_in[10]
port 225 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 io_in[11]
port 226 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 io_in[12]
port 227 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 io_in[13]
port 228 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 io_in[14]
port 229 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 io_in[15]
port 230 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 io_in[16]
port 231 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 io_in[17]
port 232 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 io_in[18]
port 233 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 io_in[19]
port 234 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 io_in[1]
port 235 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 io_in[20]
port 236 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 io_in[21]
port 237 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 io_in[22]
port 238 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 io_in[23]
port 239 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 io_in[24]
port 240 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 io_in[25]
port 241 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 io_in[26]
port 242 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 io_in[27]
port 243 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 io_in[28]
port 244 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 io_in[29]
port 245 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_in[2]
port 246 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_in[30]
port 247 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 io_in[31]
port 248 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 io_in[32]
port 249 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 io_in[33]
port 250 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 io_in[34]
port 251 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 io_in[35]
port 252 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 io_in[36]
port 253 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 io_in[37]
port 254 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 io_in[3]
port 255 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 io_in[4]
port 256 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 io_in[5]
port 257 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 io_in[6]
port 258 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 io_in[7]
port 259 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 io_in[8]
port 260 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 io_in[9]
port 261 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 io_oeb[0]
port 262 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 io_oeb[10]
port 263 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 io_oeb[11]
port 264 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 io_oeb[12]
port 265 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 io_oeb[13]
port 266 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 io_oeb[14]
port 267 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 io_oeb[15]
port 268 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 io_oeb[16]
port 269 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 io_oeb[17]
port 270 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 io_oeb[18]
port 271 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 io_oeb[19]
port 272 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 io_oeb[1]
port 273 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 io_oeb[20]
port 274 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 io_oeb[21]
port 275 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 io_oeb[22]
port 276 nsew signal output
rlabel metal2 s 33230 0 33286 800 6 io_oeb[23]
port 277 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 io_oeb[24]
port 278 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 io_oeb[25]
port 279 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 io_oeb[26]
port 280 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 io_oeb[27]
port 281 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 io_oeb[28]
port 282 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 io_oeb[29]
port 283 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 io_oeb[2]
port 284 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 io_oeb[30]
port 285 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 io_oeb[31]
port 286 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 io_oeb[32]
port 287 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 io_oeb[33]
port 288 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 io_oeb[34]
port 289 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 io_oeb[35]
port 290 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 io_oeb[36]
port 291 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 io_oeb[37]
port 292 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 io_oeb[3]
port 293 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 io_oeb[4]
port 294 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 io_oeb[5]
port 295 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 io_oeb[6]
port 296 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 io_oeb[7]
port 297 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 io_oeb[8]
port 298 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 io_oeb[9]
port 299 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 io_out[0]
port 300 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 io_out[10]
port 301 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 io_out[11]
port 302 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 io_out[12]
port 303 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 io_out[13]
port 304 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 io_out[14]
port 305 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 io_out[15]
port 306 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 io_out[16]
port 307 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 io_out[17]
port 308 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 io_out[18]
port 309 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 io_out[19]
port 310 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 io_out[1]
port 311 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 io_out[20]
port 312 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 io_out[21]
port 313 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 io_out[22]
port 314 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 io_out[23]
port 315 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 io_out[24]
port 316 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 io_out[25]
port 317 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 io_out[26]
port 318 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 io_out[27]
port 319 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 io_out[28]
port 320 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 io_out[29]
port 321 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 io_out[2]
port 322 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 io_out[30]
port 323 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 io_out[31]
port 324 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 io_out[32]
port 325 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 io_out[33]
port 326 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 io_out[34]
port 327 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 io_out[35]
port 328 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 io_out[36]
port 329 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 io_out[37]
port 330 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 io_out[3]
port 331 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 io_out[4]
port 332 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 io_out[5]
port 333 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 io_out[6]
port 334 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 io_out[7]
port 335 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 io_out[8]
port 336 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 io_out[9]
port 337 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 oeb_6502
port 338 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 oeb_as1802
port 339 nsew signal input
rlabel metal2 s 22834 59200 22890 60000 6 oeb_as2650
port 340 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 oeb_as512512512
port 341 nsew signal input
rlabel metal3 s 59200 58624 60000 58744 6 oeb_as5401
port 342 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 oeb_mc14500
port 343 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 rst_6502
port 344 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 rst_LCD
port 345 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 rst_as1802
port 346 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 rst_as2650
port 347 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 rst_as512512512
port 348 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 rst_as5401
port 349 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 rst_counter
port 350 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 rst_diceroll
port 351 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 rst_mc14500
port 352 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 rst_posit
port 353 nsew signal output
rlabel metal3 s 0 25304 800 25424 6 rst_tbb1143
port 354 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 rst_tune
port 355 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 356 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 356 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 357 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 357 nsew ground bidirectional
rlabel metal3 s 59200 1096 60000 1216 6 wb_clk_i
port 358 nsew signal input
rlabel metal3 s 59200 1504 60000 1624 6 wb_rst_i
port 359 nsew signal input
rlabel metal3 s 59200 1912 60000 2032 6 wbs_ack_o
port 360 nsew signal output
rlabel metal3 s 59200 3544 60000 3664 6 wbs_adr_i[0]
port 361 nsew signal input
rlabel metal3 s 59200 15784 60000 15904 6 wbs_adr_i[10]
port 362 nsew signal input
rlabel metal3 s 59200 17008 60000 17128 6 wbs_adr_i[11]
port 363 nsew signal input
rlabel metal3 s 59200 18232 60000 18352 6 wbs_adr_i[12]
port 364 nsew signal input
rlabel metal3 s 59200 19456 60000 19576 6 wbs_adr_i[13]
port 365 nsew signal input
rlabel metal3 s 59200 20680 60000 20800 6 wbs_adr_i[14]
port 366 nsew signal input
rlabel metal3 s 59200 21904 60000 22024 6 wbs_adr_i[15]
port 367 nsew signal input
rlabel metal3 s 59200 23128 60000 23248 6 wbs_adr_i[16]
port 368 nsew signal input
rlabel metal3 s 59200 24352 60000 24472 6 wbs_adr_i[17]
port 369 nsew signal input
rlabel metal3 s 59200 25576 60000 25696 6 wbs_adr_i[18]
port 370 nsew signal input
rlabel metal3 s 59200 26800 60000 26920 6 wbs_adr_i[19]
port 371 nsew signal input
rlabel metal3 s 59200 4768 60000 4888 6 wbs_adr_i[1]
port 372 nsew signal input
rlabel metal3 s 59200 28024 60000 28144 6 wbs_adr_i[20]
port 373 nsew signal input
rlabel metal3 s 59200 29248 60000 29368 6 wbs_adr_i[21]
port 374 nsew signal input
rlabel metal3 s 59200 30472 60000 30592 6 wbs_adr_i[22]
port 375 nsew signal input
rlabel metal3 s 59200 31696 60000 31816 6 wbs_adr_i[23]
port 376 nsew signal input
rlabel metal3 s 59200 32920 60000 33040 6 wbs_adr_i[24]
port 377 nsew signal input
rlabel metal3 s 59200 34144 60000 34264 6 wbs_adr_i[25]
port 378 nsew signal input
rlabel metal3 s 59200 35368 60000 35488 6 wbs_adr_i[26]
port 379 nsew signal input
rlabel metal3 s 59200 36592 60000 36712 6 wbs_adr_i[27]
port 380 nsew signal input
rlabel metal3 s 59200 37816 60000 37936 6 wbs_adr_i[28]
port 381 nsew signal input
rlabel metal3 s 59200 39040 60000 39160 6 wbs_adr_i[29]
port 382 nsew signal input
rlabel metal3 s 59200 5992 60000 6112 6 wbs_adr_i[2]
port 383 nsew signal input
rlabel metal3 s 59200 40264 60000 40384 6 wbs_adr_i[30]
port 384 nsew signal input
rlabel metal3 s 59200 41488 60000 41608 6 wbs_adr_i[31]
port 385 nsew signal input
rlabel metal3 s 59200 7216 60000 7336 6 wbs_adr_i[3]
port 386 nsew signal input
rlabel metal3 s 59200 8440 60000 8560 6 wbs_adr_i[4]
port 387 nsew signal input
rlabel metal3 s 59200 9664 60000 9784 6 wbs_adr_i[5]
port 388 nsew signal input
rlabel metal3 s 59200 10888 60000 11008 6 wbs_adr_i[6]
port 389 nsew signal input
rlabel metal3 s 59200 12112 60000 12232 6 wbs_adr_i[7]
port 390 nsew signal input
rlabel metal3 s 59200 13336 60000 13456 6 wbs_adr_i[8]
port 391 nsew signal input
rlabel metal3 s 59200 14560 60000 14680 6 wbs_adr_i[9]
port 392 nsew signal input
rlabel metal3 s 59200 2320 60000 2440 6 wbs_cyc_i
port 393 nsew signal input
rlabel metal3 s 59200 3952 60000 4072 6 wbs_dat_i[0]
port 394 nsew signal input
rlabel metal3 s 59200 16192 60000 16312 6 wbs_dat_i[10]
port 395 nsew signal input
rlabel metal3 s 59200 17416 60000 17536 6 wbs_dat_i[11]
port 396 nsew signal input
rlabel metal3 s 59200 18640 60000 18760 6 wbs_dat_i[12]
port 397 nsew signal input
rlabel metal3 s 59200 19864 60000 19984 6 wbs_dat_i[13]
port 398 nsew signal input
rlabel metal3 s 59200 21088 60000 21208 6 wbs_dat_i[14]
port 399 nsew signal input
rlabel metal3 s 59200 22312 60000 22432 6 wbs_dat_i[15]
port 400 nsew signal input
rlabel metal3 s 59200 23536 60000 23656 6 wbs_dat_i[16]
port 401 nsew signal input
rlabel metal3 s 59200 24760 60000 24880 6 wbs_dat_i[17]
port 402 nsew signal input
rlabel metal3 s 59200 25984 60000 26104 6 wbs_dat_i[18]
port 403 nsew signal input
rlabel metal3 s 59200 27208 60000 27328 6 wbs_dat_i[19]
port 404 nsew signal input
rlabel metal3 s 59200 5176 60000 5296 6 wbs_dat_i[1]
port 405 nsew signal input
rlabel metal3 s 59200 28432 60000 28552 6 wbs_dat_i[20]
port 406 nsew signal input
rlabel metal3 s 59200 29656 60000 29776 6 wbs_dat_i[21]
port 407 nsew signal input
rlabel metal3 s 59200 30880 60000 31000 6 wbs_dat_i[22]
port 408 nsew signal input
rlabel metal3 s 59200 32104 60000 32224 6 wbs_dat_i[23]
port 409 nsew signal input
rlabel metal3 s 59200 33328 60000 33448 6 wbs_dat_i[24]
port 410 nsew signal input
rlabel metal3 s 59200 34552 60000 34672 6 wbs_dat_i[25]
port 411 nsew signal input
rlabel metal3 s 59200 35776 60000 35896 6 wbs_dat_i[26]
port 412 nsew signal input
rlabel metal3 s 59200 37000 60000 37120 6 wbs_dat_i[27]
port 413 nsew signal input
rlabel metal3 s 59200 38224 60000 38344 6 wbs_dat_i[28]
port 414 nsew signal input
rlabel metal3 s 59200 39448 60000 39568 6 wbs_dat_i[29]
port 415 nsew signal input
rlabel metal3 s 59200 6400 60000 6520 6 wbs_dat_i[2]
port 416 nsew signal input
rlabel metal3 s 59200 40672 60000 40792 6 wbs_dat_i[30]
port 417 nsew signal input
rlabel metal3 s 59200 41896 60000 42016 6 wbs_dat_i[31]
port 418 nsew signal input
rlabel metal3 s 59200 7624 60000 7744 6 wbs_dat_i[3]
port 419 nsew signal input
rlabel metal3 s 59200 8848 60000 8968 6 wbs_dat_i[4]
port 420 nsew signal input
rlabel metal3 s 59200 10072 60000 10192 6 wbs_dat_i[5]
port 421 nsew signal input
rlabel metal3 s 59200 11296 60000 11416 6 wbs_dat_i[6]
port 422 nsew signal input
rlabel metal3 s 59200 12520 60000 12640 6 wbs_dat_i[7]
port 423 nsew signal input
rlabel metal3 s 59200 13744 60000 13864 6 wbs_dat_i[8]
port 424 nsew signal input
rlabel metal3 s 59200 14968 60000 15088 6 wbs_dat_i[9]
port 425 nsew signal input
rlabel metal3 s 59200 4360 60000 4480 6 wbs_dat_o[0]
port 426 nsew signal output
rlabel metal3 s 59200 16600 60000 16720 6 wbs_dat_o[10]
port 427 nsew signal output
rlabel metal3 s 59200 17824 60000 17944 6 wbs_dat_o[11]
port 428 nsew signal output
rlabel metal3 s 59200 19048 60000 19168 6 wbs_dat_o[12]
port 429 nsew signal output
rlabel metal3 s 59200 20272 60000 20392 6 wbs_dat_o[13]
port 430 nsew signal output
rlabel metal3 s 59200 21496 60000 21616 6 wbs_dat_o[14]
port 431 nsew signal output
rlabel metal3 s 59200 22720 60000 22840 6 wbs_dat_o[15]
port 432 nsew signal output
rlabel metal3 s 59200 23944 60000 24064 6 wbs_dat_o[16]
port 433 nsew signal output
rlabel metal3 s 59200 25168 60000 25288 6 wbs_dat_o[17]
port 434 nsew signal output
rlabel metal3 s 59200 26392 60000 26512 6 wbs_dat_o[18]
port 435 nsew signal output
rlabel metal3 s 59200 27616 60000 27736 6 wbs_dat_o[19]
port 436 nsew signal output
rlabel metal3 s 59200 5584 60000 5704 6 wbs_dat_o[1]
port 437 nsew signal output
rlabel metal3 s 59200 28840 60000 28960 6 wbs_dat_o[20]
port 438 nsew signal output
rlabel metal3 s 59200 30064 60000 30184 6 wbs_dat_o[21]
port 439 nsew signal output
rlabel metal3 s 59200 31288 60000 31408 6 wbs_dat_o[22]
port 440 nsew signal output
rlabel metal3 s 59200 32512 60000 32632 6 wbs_dat_o[23]
port 441 nsew signal output
rlabel metal3 s 59200 33736 60000 33856 6 wbs_dat_o[24]
port 442 nsew signal output
rlabel metal3 s 59200 34960 60000 35080 6 wbs_dat_o[25]
port 443 nsew signal output
rlabel metal3 s 59200 36184 60000 36304 6 wbs_dat_o[26]
port 444 nsew signal output
rlabel metal3 s 59200 37408 60000 37528 6 wbs_dat_o[27]
port 445 nsew signal output
rlabel metal3 s 59200 38632 60000 38752 6 wbs_dat_o[28]
port 446 nsew signal output
rlabel metal3 s 59200 39856 60000 39976 6 wbs_dat_o[29]
port 447 nsew signal output
rlabel metal3 s 59200 6808 60000 6928 6 wbs_dat_o[2]
port 448 nsew signal output
rlabel metal3 s 59200 41080 60000 41200 6 wbs_dat_o[30]
port 449 nsew signal output
rlabel metal3 s 59200 42304 60000 42424 6 wbs_dat_o[31]
port 450 nsew signal output
rlabel metal3 s 59200 8032 60000 8152 6 wbs_dat_o[3]
port 451 nsew signal output
rlabel metal3 s 59200 9256 60000 9376 6 wbs_dat_o[4]
port 452 nsew signal output
rlabel metal3 s 59200 10480 60000 10600 6 wbs_dat_o[5]
port 453 nsew signal output
rlabel metal3 s 59200 11704 60000 11824 6 wbs_dat_o[6]
port 454 nsew signal output
rlabel metal3 s 59200 12928 60000 13048 6 wbs_dat_o[7]
port 455 nsew signal output
rlabel metal3 s 59200 14152 60000 14272 6 wbs_dat_o[8]
port 456 nsew signal output
rlabel metal3 s 59200 15376 60000 15496 6 wbs_dat_o[9]
port 457 nsew signal output
rlabel metal3 s 59200 2728 60000 2848 6 wbs_stb_i
port 458 nsew signal input
rlabel metal3 s 59200 3136 60000 3256 6 wbs_we_i
port 459 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4541726
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/Multiplexer/runs/23_03_28_15_02/results/signoff/multiplexer.magic.gds
string GDS_START 721888
<< end >>

