magic
tech sky130B
magscale 1 2
timestamp 1676316617
<< obsli1 >>
rect 1104 2159 63848 62577
<< obsm1 >>
rect 1104 1708 63848 62608
<< metal2 >>
rect 1370 0 1482 800
rect 3670 0 3782 800
rect 5970 0 6082 800
rect 8270 0 8382 800
rect 10570 0 10682 800
rect 12870 0 12982 800
rect 15170 0 15282 800
rect 17470 0 17582 800
rect 19770 0 19882 800
rect 22070 0 22182 800
rect 24370 0 24482 800
rect 26670 0 26782 800
rect 28970 0 29082 800
rect 31270 0 31382 800
rect 33570 0 33682 800
rect 35870 0 35982 800
rect 38170 0 38282 800
rect 40470 0 40582 800
rect 42770 0 42882 800
rect 45070 0 45182 800
rect 47370 0 47482 800
rect 49670 0 49782 800
rect 51970 0 52082 800
rect 54270 0 54382 800
rect 56570 0 56682 800
rect 58870 0 58982 800
rect 61170 0 61282 800
rect 63470 0 63582 800
<< obsm2 >>
rect 1398 856 63552 62597
rect 1538 800 3614 856
rect 3838 800 5914 856
rect 6138 800 8214 856
rect 8438 800 10514 856
rect 10738 800 12814 856
rect 13038 800 15114 856
rect 15338 800 17414 856
rect 17638 800 19714 856
rect 19938 800 22014 856
rect 22238 800 24314 856
rect 24538 800 26614 856
rect 26838 800 28914 856
rect 29138 800 31214 856
rect 31438 800 33514 856
rect 33738 800 35814 856
rect 36038 800 38114 856
rect 38338 800 40414 856
rect 40638 800 42714 856
rect 42938 800 45014 856
rect 45238 800 47314 856
rect 47538 800 49614 856
rect 49838 800 51914 856
rect 52138 800 54214 856
rect 54438 800 56514 856
rect 56738 800 58814 856
rect 59038 800 61114 856
rect 61338 800 63414 856
<< metal3 >>
rect 0 61828 800 62068
rect 0 57612 800 57852
rect 0 53396 800 53636
rect 0 49180 800 49420
rect 0 44964 800 45204
rect 0 40748 800 40988
rect 0 36532 800 36772
rect 0 32316 800 32556
rect 0 28100 800 28340
rect 0 23884 800 24124
rect 0 19668 800 19908
rect 0 15452 800 15692
rect 0 11236 800 11476
rect 0 7020 800 7260
rect 0 2804 800 3044
<< obsm3 >>
rect 614 62148 60799 62593
rect 880 61748 60799 62148
rect 614 57932 60799 61748
rect 880 57532 60799 57932
rect 614 53716 60799 57532
rect 880 53316 60799 53716
rect 614 49500 60799 53316
rect 880 49100 60799 49500
rect 614 45284 60799 49100
rect 880 44884 60799 45284
rect 614 41068 60799 44884
rect 880 40668 60799 41068
rect 614 36852 60799 40668
rect 880 36452 60799 36852
rect 614 32636 60799 36452
rect 880 32236 60799 32636
rect 614 28420 60799 32236
rect 880 28020 60799 28420
rect 614 24204 60799 28020
rect 880 23804 60799 24204
rect 614 19988 60799 23804
rect 880 19588 60799 19988
rect 614 15772 60799 19588
rect 880 15372 60799 15772
rect 614 11556 60799 15372
rect 880 11156 60799 11556
rect 614 7340 60799 11156
rect 880 6940 60799 7340
rect 614 3124 60799 6940
rect 880 2724 60799 3124
rect 614 1939 60799 2724
<< metal4 >>
rect 4208 2128 4528 62608
rect 19568 2128 19888 62608
rect 34928 2128 35248 62608
rect 50288 2128 50608 62608
<< obsm4 >>
rect 1899 2048 4128 57765
rect 4608 2048 19488 57765
rect 19968 2048 34848 57765
rect 35328 2048 50208 57765
rect 50688 2048 58269 57765
rect 1899 1939 58269 2048
<< labels >>
rlabel metal3 s 0 57612 800 57852 6 clk
port 1 nsew signal input
rlabel metal3 s 0 2804 800 3044 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 0 44964 800 45204 6 io_in[10]
port 3 nsew signal input
rlabel metal3 s 0 49180 800 49420 6 io_in[11]
port 4 nsew signal input
rlabel metal3 s 0 53396 800 53636 6 io_in[12]
port 5 nsew signal input
rlabel metal3 s 0 7020 800 7260 6 io_in[1]
port 6 nsew signal input
rlabel metal3 s 0 11236 800 11476 6 io_in[2]
port 7 nsew signal input
rlabel metal3 s 0 15452 800 15692 6 io_in[3]
port 8 nsew signal input
rlabel metal3 s 0 19668 800 19908 6 io_in[4]
port 9 nsew signal input
rlabel metal3 s 0 23884 800 24124 6 io_in[5]
port 10 nsew signal input
rlabel metal3 s 0 28100 800 28340 6 io_in[6]
port 11 nsew signal input
rlabel metal3 s 0 32316 800 32556 6 io_in[7]
port 12 nsew signal input
rlabel metal3 s 0 36532 800 36772 6 io_in[8]
port 13 nsew signal input
rlabel metal3 s 0 40748 800 40988 6 io_in[9]
port 14 nsew signal input
rlabel metal2 s 63470 0 63582 800 6 io_oeb
port 15 nsew signal output
rlabel metal2 s 1370 0 1482 800 6 io_out[0]
port 16 nsew signal output
rlabel metal2 s 24370 0 24482 800 6 io_out[10]
port 17 nsew signal output
rlabel metal2 s 26670 0 26782 800 6 io_out[11]
port 18 nsew signal output
rlabel metal2 s 28970 0 29082 800 6 io_out[12]
port 19 nsew signal output
rlabel metal2 s 31270 0 31382 800 6 io_out[13]
port 20 nsew signal output
rlabel metal2 s 33570 0 33682 800 6 io_out[14]
port 21 nsew signal output
rlabel metal2 s 35870 0 35982 800 6 io_out[15]
port 22 nsew signal output
rlabel metal2 s 38170 0 38282 800 6 io_out[16]
port 23 nsew signal output
rlabel metal2 s 40470 0 40582 800 6 io_out[17]
port 24 nsew signal output
rlabel metal2 s 42770 0 42882 800 6 io_out[18]
port 25 nsew signal output
rlabel metal2 s 45070 0 45182 800 6 io_out[19]
port 26 nsew signal output
rlabel metal2 s 3670 0 3782 800 6 io_out[1]
port 27 nsew signal output
rlabel metal2 s 47370 0 47482 800 6 io_out[20]
port 28 nsew signal output
rlabel metal2 s 49670 0 49782 800 6 io_out[21]
port 29 nsew signal output
rlabel metal2 s 51970 0 52082 800 6 io_out[22]
port 30 nsew signal output
rlabel metal2 s 54270 0 54382 800 6 io_out[23]
port 31 nsew signal output
rlabel metal2 s 56570 0 56682 800 6 io_out[24]
port 32 nsew signal output
rlabel metal2 s 58870 0 58982 800 6 io_out[25]
port 33 nsew signal output
rlabel metal2 s 61170 0 61282 800 6 io_out[26]
port 34 nsew signal output
rlabel metal2 s 5970 0 6082 800 6 io_out[2]
port 35 nsew signal output
rlabel metal2 s 8270 0 8382 800 6 io_out[3]
port 36 nsew signal output
rlabel metal2 s 10570 0 10682 800 6 io_out[4]
port 37 nsew signal output
rlabel metal2 s 12870 0 12982 800 6 io_out[5]
port 38 nsew signal output
rlabel metal2 s 15170 0 15282 800 6 io_out[6]
port 39 nsew signal output
rlabel metal2 s 17470 0 17582 800 6 io_out[7]
port 40 nsew signal output
rlabel metal2 s 19770 0 19882 800 6 io_out[8]
port 41 nsew signal output
rlabel metal2 s 22070 0 22182 800 6 io_out[9]
port 42 nsew signal output
rlabel metal3 s 0 61828 800 62068 6 rst
port 43 nsew signal input
rlabel metal4 s 4208 2128 4528 62608 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 62608 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 62608 6 vssd1
port 45 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 62608 6 vssd1
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 65000 65000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13107830
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/AS1802/runs/23_02_13_20_22/results/signoff/wrapped_as1802.magic.gds
string GDS_START 960974
<< end >>

