VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt2_tholin_multiplexed_counter
  CLASS BLOCK ;
  FOREIGN tt2_tholin_multiplexed_counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 90.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 86.000 22.450 90.000 ;
    END
  END clk
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END io_out[11]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 86.000 67.530 90.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.550 10.640 16.150 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.215 10.640 35.815 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.880 10.640 55.480 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.545 10.640 75.145 79.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.380 10.640 25.980 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.045 10.640 45.645 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.710 10.640 65.310 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.375 10.640 84.975 79.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 84.180 78.965 ;
      LAYER met1 ;
        RECT 4.210 10.640 85.490 79.120 ;
      LAYER met2 ;
        RECT 4.240 85.720 21.890 86.000 ;
        RECT 22.730 85.720 66.970 86.000 ;
        RECT 67.810 85.720 85.460 86.000 ;
        RECT 4.240 4.280 85.460 85.720 ;
        RECT 4.790 4.000 11.310 4.280 ;
        RECT 12.150 4.000 18.670 4.280 ;
        RECT 19.510 4.000 26.030 4.280 ;
        RECT 26.870 4.000 33.390 4.280 ;
        RECT 34.230 4.000 40.750 4.280 ;
        RECT 41.590 4.000 48.110 4.280 ;
        RECT 48.950 4.000 55.470 4.280 ;
        RECT 56.310 4.000 62.830 4.280 ;
        RECT 63.670 4.000 70.190 4.280 ;
        RECT 71.030 4.000 77.550 4.280 ;
        RECT 78.390 4.000 84.910 4.280 ;
      LAYER met3 ;
        RECT 14.560 10.715 84.965 79.045 ;
  END
END tt2_tholin_multiplexed_counter
END LIBRARY

