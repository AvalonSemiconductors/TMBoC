magic
tech sky130B
magscale 1 2
timestamp 1680267168
<< viali >>
rect 1961 61285 1995 61319
rect 9689 61285 9723 61319
rect 20729 61285 20763 61319
rect 49525 61217 49559 61251
rect 2513 61149 2547 61183
rect 4353 61149 4387 61183
rect 5089 61149 5123 61183
rect 5825 61149 5859 61183
rect 6745 61149 6779 61183
rect 7573 61149 7607 61183
rect 7849 61149 7883 61183
rect 9505 61149 9539 61183
rect 10241 61149 10275 61183
rect 10977 61149 11011 61183
rect 12449 61149 12483 61183
rect 13277 61149 13311 61183
rect 14381 61149 14415 61183
rect 15393 61149 15427 61183
rect 16129 61149 16163 61183
rect 17233 61149 17267 61183
rect 17969 61149 18003 61183
rect 18705 61149 18739 61183
rect 19809 61149 19843 61183
rect 20545 61149 20579 61183
rect 21281 61149 21315 61183
rect 22385 61149 22419 61183
rect 23121 61149 23155 61183
rect 23857 61149 23891 61183
rect 25329 61149 25363 61183
rect 26065 61149 26099 61183
rect 27537 61149 27571 61183
rect 28365 61149 28399 61183
rect 29837 61149 29871 61183
rect 31217 61149 31251 61183
rect 32413 61149 32447 61183
rect 33057 61149 33091 61183
rect 33793 61149 33827 61183
rect 34989 61149 35023 61183
rect 35909 61149 35943 61183
rect 37565 61149 37599 61183
rect 38301 61149 38335 61183
rect 39037 61149 39071 61183
rect 40785 61149 40819 61183
rect 41613 61149 41647 61183
rect 42717 61149 42751 61183
rect 43637 61149 43671 61183
rect 44373 61149 44407 61183
rect 45293 61149 45327 61183
rect 46029 61149 46063 61183
rect 46765 61149 46799 61183
rect 47869 61149 47903 61183
rect 48605 61149 48639 61183
rect 49341 61149 49375 61183
rect 51089 61149 51123 61183
rect 52009 61149 52043 61183
rect 53205 61149 53239 61183
rect 54217 61149 54251 61183
rect 56149 61149 56183 61183
rect 57161 61149 57195 61183
rect 58081 61149 58115 61183
rect 1685 61081 1719 61115
rect 2789 61081 2823 61115
rect 4537 61081 4571 61115
rect 13553 61081 13587 61115
rect 15577 61081 15611 61115
rect 16313 61081 16347 61115
rect 18153 61081 18187 61115
rect 19993 61081 20027 61115
rect 26433 61081 26467 61115
rect 37749 61081 37783 61115
rect 40141 61081 40175 61115
rect 46949 61081 46983 61115
rect 53481 61081 53515 61115
rect 54401 61081 54435 61115
rect 56425 61081 56459 61115
rect 5181 61013 5215 61047
rect 5917 61013 5951 61047
rect 7021 61013 7055 61047
rect 10333 61013 10367 61047
rect 11069 61013 11103 61047
rect 12541 61013 12575 61047
rect 14473 61013 14507 61047
rect 17325 61013 17359 61047
rect 18797 61013 18831 61047
rect 21373 61013 21407 61047
rect 22477 61013 22511 61047
rect 23213 61013 23247 61047
rect 23949 61013 23983 61047
rect 25421 61013 25455 61047
rect 27629 61013 27663 61047
rect 28549 61013 28583 61047
rect 29929 61013 29963 61047
rect 31309 61013 31343 61047
rect 32505 61013 32539 61047
rect 33241 61013 33275 61047
rect 33977 61013 34011 61047
rect 35081 61013 35115 61047
rect 36001 61013 36035 61047
rect 38393 61013 38427 61047
rect 39129 61013 39163 61047
rect 40233 61013 40267 61047
rect 40969 61013 41003 61047
rect 41705 61013 41739 61047
rect 42809 61013 42843 61047
rect 43729 61013 43763 61047
rect 44465 61013 44499 61047
rect 45385 61013 45419 61047
rect 46121 61013 46155 61047
rect 47961 61013 47995 61047
rect 48697 61013 48731 61047
rect 51181 61013 51215 61047
rect 52101 61013 52135 61047
rect 57253 61013 57287 61047
rect 58265 61013 58299 61047
rect 1685 60741 1719 60775
rect 3249 60741 3283 60775
rect 3985 60741 4019 60775
rect 8401 60741 8435 60775
rect 9137 60741 9171 60775
rect 12081 60741 12115 60775
rect 15025 60741 15059 60775
rect 19441 60741 19475 60775
rect 24593 60741 24627 60775
rect 34161 60741 34195 60775
rect 36369 60741 36403 60775
rect 46673 60741 46707 60775
rect 50353 60741 50387 60775
rect 53021 60741 53055 60775
rect 54769 60741 54803 60775
rect 55505 60741 55539 60775
rect 57161 60741 57195 60775
rect 58173 60741 58207 60775
rect 27169 60673 27203 60707
rect 29653 60673 29687 60707
rect 30389 60673 30423 60707
rect 41429 60673 41463 60707
rect 49525 60673 49559 60707
rect 56149 60673 56183 60707
rect 9321 60605 9355 60639
rect 56333 60605 56367 60639
rect 4169 60537 4203 60571
rect 8585 60537 8619 60571
rect 15209 60537 15243 60571
rect 19625 60537 19659 60571
rect 24777 60537 24811 60571
rect 1961 60469 1995 60503
rect 3341 60469 3375 60503
rect 12173 60469 12207 60503
rect 27353 60469 27387 60503
rect 29837 60469 29871 60503
rect 30573 60469 30607 60503
rect 34253 60469 34287 60503
rect 36461 60469 36495 60503
rect 41613 60469 41647 60503
rect 46765 60469 46799 60503
rect 49709 60469 49743 60503
rect 50445 60469 50479 60503
rect 53113 60469 53147 60503
rect 54861 60469 54895 60503
rect 55597 60469 55631 60503
rect 57253 60469 57287 60503
rect 58265 60469 58299 60503
rect 57253 60197 57287 60231
rect 1777 60061 1811 60095
rect 2513 60061 2547 60095
rect 56241 60061 56275 60095
rect 1961 59993 1995 60027
rect 57069 59993 57103 60027
rect 57989 59993 58023 60027
rect 58357 59993 58391 60027
rect 2605 59925 2639 59959
rect 56333 59925 56367 59959
rect 2421 59653 2455 59687
rect 1593 59585 1627 59619
rect 57069 59585 57103 59619
rect 58081 59585 58115 59619
rect 57253 59517 57287 59551
rect 2605 59449 2639 59483
rect 1777 59381 1811 59415
rect 58265 59381 58299 59415
rect 43913 59041 43947 59075
rect 44373 59041 44407 59075
rect 1593 58973 1627 59007
rect 44097 58973 44131 59007
rect 44465 58973 44499 59007
rect 57253 58973 57287 59007
rect 57989 58905 58023 58939
rect 1777 58837 1811 58871
rect 43729 58837 43763 58871
rect 57345 58837 57379 58871
rect 58081 58837 58115 58871
rect 15117 58565 15151 58599
rect 17141 58565 17175 58599
rect 17233 58565 17267 58599
rect 1685 58497 1719 58531
rect 14841 58497 14875 58531
rect 15025 58497 15059 58531
rect 15261 58497 15295 58531
rect 16957 58497 16991 58531
rect 17377 58497 17411 58531
rect 39497 58497 39531 58531
rect 39681 58497 39715 58531
rect 39773 58497 39807 58531
rect 39917 58497 39951 58531
rect 58173 58497 58207 58531
rect 14565 58429 14599 58463
rect 1961 58361 1995 58395
rect 15393 58293 15427 58327
rect 17509 58293 17543 58327
rect 40049 58293 40083 58327
rect 58265 58293 58299 58327
rect 43913 57953 43947 57987
rect 44373 57953 44407 57987
rect 1593 57885 1627 57919
rect 21281 57885 21315 57919
rect 21373 57885 21407 57919
rect 21649 57885 21683 57919
rect 21925 57885 21959 57919
rect 22109 57885 22143 57919
rect 22753 57885 22787 57919
rect 22846 57885 22880 57919
rect 23029 57885 23063 57919
rect 23218 57885 23252 57919
rect 24593 57885 24627 57919
rect 24966 57885 25000 57919
rect 31861 57885 31895 57919
rect 31953 57885 31987 57919
rect 32229 57885 32263 57919
rect 32505 57885 32539 57919
rect 32689 57885 32723 57919
rect 38669 57885 38703 57919
rect 44097 57885 44131 57919
rect 44465 57885 44499 57919
rect 54125 57885 54159 57919
rect 54545 57885 54579 57919
rect 23121 57817 23155 57851
rect 24777 57817 24811 57851
rect 24869 57817 24903 57851
rect 38485 57817 38519 57851
rect 38945 57817 38979 57851
rect 54309 57817 54343 57851
rect 54401 57817 54435 57851
rect 58173 57817 58207 57851
rect 1777 57749 1811 57783
rect 20913 57749 20947 57783
rect 23397 57749 23431 57783
rect 25162 57749 25196 57783
rect 31493 57749 31527 57783
rect 38853 57749 38887 57783
rect 43729 57749 43763 57783
rect 54685 57749 54719 57783
rect 58265 57749 58299 57783
rect 20729 57545 20763 57579
rect 38669 57545 38703 57579
rect 20453 57477 20487 57511
rect 38393 57477 38427 57511
rect 19901 57409 19935 57443
rect 20177 57409 20211 57443
rect 20361 57409 20395 57443
rect 20545 57409 20579 57443
rect 30757 57409 30791 57443
rect 31033 57409 31067 57443
rect 31125 57409 31159 57443
rect 31401 57409 31435 57443
rect 31585 57409 31619 57443
rect 35725 57409 35759 57443
rect 36001 57409 36035 57443
rect 36093 57409 36127 57443
rect 36369 57409 36403 57443
rect 36645 57409 36679 57443
rect 38117 57409 38151 57443
rect 38301 57409 38335 57443
rect 38485 57409 38519 57443
rect 54445 57409 54479 57443
rect 54861 57409 54895 57443
rect 55045 57409 55079 57443
rect 58173 57409 58207 57443
rect 53941 57341 53975 57375
rect 54309 57341 54343 57375
rect 58357 57273 58391 57307
rect 30389 57205 30423 57239
rect 35357 57205 35391 57239
rect 22293 56933 22327 56967
rect 54125 56865 54159 56899
rect 58357 56865 58391 56899
rect 1685 56797 1719 56831
rect 21649 56797 21683 56831
rect 21742 56797 21776 56831
rect 21925 56797 21959 56831
rect 22155 56797 22189 56831
rect 43913 56797 43947 56831
rect 44097 56797 44131 56831
rect 44465 56797 44499 56831
rect 44557 56797 44591 56831
rect 54033 56797 54067 56831
rect 54401 56797 54435 56831
rect 54585 56797 54619 56831
rect 22017 56729 22051 56763
rect 58173 56729 58207 56763
rect 1961 56661 1995 56695
rect 43729 56661 43763 56695
rect 53481 56661 53515 56695
rect 15669 56389 15703 56423
rect 33793 56389 33827 56423
rect 34621 56389 34655 56423
rect 1685 56321 1719 56355
rect 15393 56321 15427 56355
rect 15577 56321 15611 56355
rect 15761 56321 15795 56355
rect 29469 56321 29503 56355
rect 29653 56321 29687 56355
rect 29745 56321 29779 56355
rect 29889 56321 29923 56355
rect 33609 56321 33643 56355
rect 33885 56321 33919 56355
rect 33977 56321 34011 56355
rect 34989 56253 35023 56287
rect 15945 56185 15979 56219
rect 34897 56185 34931 56219
rect 1777 56117 1811 56151
rect 30021 56117 30055 56151
rect 34161 56117 34195 56151
rect 34759 56117 34793 56151
rect 35265 56117 35299 56151
rect 58357 56117 58391 56151
rect 1685 55641 1719 55675
rect 1961 55573 1995 55607
rect 1777 55369 1811 55403
rect 43269 55369 43303 55403
rect 1593 55233 1627 55267
rect 43453 55233 43487 55267
rect 43637 55233 43671 55267
rect 44005 55233 44039 55267
rect 43913 55165 43947 55199
rect 58357 54621 58391 54655
rect 1685 54145 1719 54179
rect 43269 54145 43303 54179
rect 43637 54145 43671 54179
rect 42717 54077 42751 54111
rect 43085 54077 43119 54111
rect 43545 54077 43579 54111
rect 1961 53941 1995 53975
rect 1593 53533 1627 53567
rect 1777 53397 1811 53431
rect 1593 53057 1627 53091
rect 1777 52853 1811 52887
rect 58357 52853 58391 52887
rect 1869 52445 1903 52479
rect 1685 52377 1719 52411
rect 5457 52037 5491 52071
rect 5181 51969 5215 52003
rect 5365 51969 5399 52003
rect 5601 51969 5635 52003
rect 5733 51765 5767 51799
rect 22477 51357 22511 51391
rect 22570 51357 22604 51391
rect 22983 51357 23017 51391
rect 58357 51357 58391 51391
rect 1685 51289 1719 51323
rect 22753 51289 22787 51323
rect 22845 51289 22879 51323
rect 1777 51221 1811 51255
rect 23121 51221 23155 51255
rect 1685 50881 1719 50915
rect 1869 50745 1903 50779
rect 57897 50269 57931 50303
rect 1685 50201 1719 50235
rect 58173 50201 58207 50235
rect 1777 50133 1811 50167
rect 20821 49861 20855 49895
rect 1685 49793 1719 49827
rect 20545 49793 20579 49827
rect 20729 49793 20763 49827
rect 20913 49793 20947 49827
rect 1869 49725 1903 49759
rect 21097 49589 21131 49623
rect 21741 49385 21775 49419
rect 21189 49181 21223 49215
rect 21557 49181 21591 49215
rect 21373 49113 21407 49147
rect 21465 49113 21499 49147
rect 57989 49113 58023 49147
rect 58357 49113 58391 49147
rect 19993 48773 20027 48807
rect 1685 48705 1719 48739
rect 19717 48705 19751 48739
rect 19901 48705 19935 48739
rect 20085 48705 20119 48739
rect 22017 48705 22051 48739
rect 22110 48705 22144 48739
rect 22293 48705 22327 48739
rect 22385 48705 22419 48739
rect 22482 48705 22516 48739
rect 23029 48637 23063 48671
rect 1777 48501 1811 48535
rect 20269 48501 20303 48535
rect 22661 48501 22695 48535
rect 56977 48093 57011 48127
rect 1685 48025 1719 48059
rect 57253 48025 57287 48059
rect 57989 48025 58023 48059
rect 58357 48025 58391 48059
rect 1777 47957 1811 47991
rect 1685 47617 1719 47651
rect 1777 47413 1811 47447
rect 1869 47005 1903 47039
rect 57897 47005 57931 47039
rect 1685 46937 1719 46971
rect 58173 46937 58207 46971
rect 22845 45917 22879 45951
rect 23029 45917 23063 45951
rect 23213 45917 23247 45951
rect 1685 45849 1719 45883
rect 23121 45849 23155 45883
rect 57989 45849 58023 45883
rect 58357 45849 58391 45883
rect 1777 45781 1811 45815
rect 22569 45781 22603 45815
rect 23397 45781 23431 45815
rect 1593 45441 1627 45475
rect 1777 45237 1811 45271
rect 1869 44965 1903 44999
rect 56977 44829 57011 44863
rect 1685 44761 1719 44795
rect 57253 44761 57287 44795
rect 57989 44761 58023 44795
rect 58357 44761 58391 44795
rect 1685 44353 1719 44387
rect 1777 44149 1811 44183
rect 15485 43809 15519 43843
rect 15669 43741 15703 43775
rect 16037 43741 16071 43775
rect 16221 43741 16255 43775
rect 57897 43741 57931 43775
rect 58173 43673 58207 43707
rect 15117 43605 15151 43639
rect 1593 43265 1627 43299
rect 1777 43061 1811 43095
rect 23305 42721 23339 42755
rect 23029 42653 23063 42687
rect 56977 42653 57011 42687
rect 57897 42653 57931 42687
rect 1685 42585 1719 42619
rect 2053 42585 2087 42619
rect 57253 42585 57287 42619
rect 58173 42585 58207 42619
rect 1869 42245 1903 42279
rect 4721 42245 4755 42279
rect 1685 42177 1719 42211
rect 4445 42177 4479 42211
rect 4629 42177 4663 42211
rect 4813 42177 4847 42211
rect 22937 42177 22971 42211
rect 23121 42177 23155 42211
rect 23489 42109 23523 42143
rect 4997 41973 5031 42007
rect 22661 41769 22695 41803
rect 22845 41565 22879 41599
rect 22937 41565 22971 41599
rect 23121 41565 23155 41599
rect 23213 41565 23247 41599
rect 56977 41565 57011 41599
rect 1685 41497 1719 41531
rect 1869 41497 1903 41531
rect 57253 41497 57287 41531
rect 57989 41497 58023 41531
rect 58357 41497 58391 41531
rect 3985 41157 4019 41191
rect 1685 41089 1719 41123
rect 3709 41089 3743 41123
rect 3893 41089 3927 41123
rect 4082 41089 4116 41123
rect 1869 40953 1903 40987
rect 4261 40885 4295 40919
rect 22661 40477 22695 40511
rect 23029 40477 23063 40511
rect 57897 40477 57931 40511
rect 1685 40409 1719 40443
rect 22845 40409 22879 40443
rect 22937 40409 22971 40443
rect 58173 40409 58207 40443
rect 1777 40341 1811 40375
rect 23213 40341 23247 40375
rect 1685 40069 1719 40103
rect 2789 40069 2823 40103
rect 58173 40069 58207 40103
rect 2513 40001 2547 40035
rect 2697 40001 2731 40035
rect 2933 40001 2967 40035
rect 1869 39865 1903 39899
rect 3065 39797 3099 39831
rect 58265 39797 58299 39831
rect 23397 39457 23431 39491
rect 23121 39389 23155 39423
rect 1685 39321 1719 39355
rect 1869 39321 1903 39355
rect 57069 39321 57103 39355
rect 57989 39321 58023 39355
rect 58357 39321 58391 39355
rect 57161 39253 57195 39287
rect 20821 38981 20855 39015
rect 22937 38981 22971 39015
rect 1685 38913 1719 38947
rect 20453 38913 20487 38947
rect 20601 38913 20635 38947
rect 20729 38913 20763 38947
rect 20959 38913 20993 38947
rect 22661 38913 22695 38947
rect 22845 38913 22879 38947
rect 23034 38913 23068 38947
rect 1777 38709 1811 38743
rect 21097 38709 21131 38743
rect 23213 38709 23247 38743
rect 21465 38437 21499 38471
rect 20269 38369 20303 38403
rect 2421 38301 2455 38335
rect 2513 38301 2547 38335
rect 2789 38301 2823 38335
rect 3065 38301 3099 38335
rect 3249 38301 3283 38335
rect 20085 38301 20119 38335
rect 21373 38301 21407 38335
rect 21649 38301 21683 38335
rect 56977 38301 57011 38335
rect 57897 38301 57931 38335
rect 57253 38233 57287 38267
rect 58173 38233 58207 38267
rect 2053 38165 2087 38199
rect 21833 38165 21867 38199
rect 2697 37961 2731 37995
rect 2421 37893 2455 37927
rect 11989 37893 12023 37927
rect 2145 37825 2179 37859
rect 2329 37825 2363 37859
rect 2513 37825 2547 37859
rect 11713 37825 11747 37859
rect 11897 37825 11931 37859
rect 12081 37825 12115 37859
rect 18705 37825 18739 37859
rect 18889 37825 18923 37859
rect 18981 37825 19015 37859
rect 19119 37825 19153 37859
rect 19717 37825 19751 37859
rect 21465 37825 21499 37859
rect 22293 37825 22327 37859
rect 22753 37825 22787 37859
rect 22845 37825 22879 37859
rect 23213 37825 23247 37859
rect 1869 37757 1903 37791
rect 18429 37757 18463 37791
rect 23489 37757 23523 37791
rect 12265 37689 12299 37723
rect 19257 37689 19291 37723
rect 22477 37417 22511 37451
rect 2605 37281 2639 37315
rect 1593 37213 1627 37247
rect 19441 37213 19475 37247
rect 19717 37213 19751 37247
rect 19809 37213 19843 37247
rect 20545 37213 20579 37247
rect 21925 37213 21959 37247
rect 22293 37213 22327 37247
rect 45201 37213 45235 37247
rect 45477 37213 45511 37247
rect 45569 37213 45603 37247
rect 46489 37213 46523 37247
rect 46765 37213 46799 37247
rect 57897 37213 57931 37247
rect 2421 37145 2455 37179
rect 19625 37145 19659 37179
rect 21281 37145 21315 37179
rect 22109 37145 22143 37179
rect 22201 37145 22235 37179
rect 45385 37145 45419 37179
rect 46305 37145 46339 37179
rect 58173 37145 58207 37179
rect 1777 37077 1811 37111
rect 19993 37077 20027 37111
rect 45753 37077 45787 37111
rect 46673 37077 46707 37111
rect 21373 36873 21407 36907
rect 20453 36805 20487 36839
rect 21097 36805 21131 36839
rect 45661 36805 45695 36839
rect 1685 36737 1719 36771
rect 20729 36737 20763 36771
rect 20877 36737 20911 36771
rect 21005 36737 21039 36771
rect 21194 36737 21228 36771
rect 23121 36737 23155 36771
rect 23213 36737 23247 36771
rect 23397 36737 23431 36771
rect 23489 36737 23523 36771
rect 45385 36737 45419 36771
rect 1777 36533 1811 36567
rect 22937 36533 22971 36567
rect 1777 36329 1811 36363
rect 21925 36261 21959 36295
rect 22477 36261 22511 36295
rect 25145 36261 25179 36295
rect 18245 36125 18279 36159
rect 18613 36125 18647 36159
rect 21373 36125 21407 36159
rect 21649 36125 21683 36159
rect 21741 36125 21775 36159
rect 22385 36125 22419 36159
rect 22661 36125 22695 36159
rect 24593 36125 24627 36159
rect 24961 36125 24995 36159
rect 1685 36057 1719 36091
rect 21557 36057 21591 36091
rect 23121 36057 23155 36091
rect 24777 36057 24811 36091
rect 24869 36057 24903 36091
rect 57989 36057 58023 36091
rect 58357 36057 58391 36091
rect 21465 35785 21499 35819
rect 2329 35717 2363 35751
rect 18245 35717 18279 35751
rect 21097 35717 21131 35751
rect 2053 35649 2087 35683
rect 2237 35649 2271 35683
rect 2426 35649 2460 35683
rect 18429 35649 18463 35683
rect 18521 35649 18555 35683
rect 18705 35649 18739 35683
rect 18797 35649 18831 35683
rect 20821 35649 20855 35683
rect 20914 35649 20948 35683
rect 21189 35649 21223 35683
rect 21286 35649 21320 35683
rect 22017 35649 22051 35683
rect 24961 35649 24995 35683
rect 25053 35649 25087 35683
rect 25329 35649 25363 35683
rect 23213 35581 23247 35615
rect 25421 35581 25455 35615
rect 20545 35513 20579 35547
rect 2605 35445 2639 35479
rect 24409 35445 24443 35479
rect 22247 35241 22281 35275
rect 22385 35241 22419 35275
rect 24869 35241 24903 35275
rect 2605 35173 2639 35207
rect 23765 35173 23799 35207
rect 22477 35105 22511 35139
rect 2053 35037 2087 35071
rect 2237 35037 2271 35071
rect 2426 35037 2460 35071
rect 16221 35037 16255 35071
rect 16313 35037 16347 35071
rect 16589 35037 16623 35071
rect 16865 35037 16899 35071
rect 17049 35037 17083 35071
rect 21373 35037 21407 35071
rect 21649 35037 21683 35071
rect 22109 35037 22143 35071
rect 23765 35037 23799 35071
rect 24041 35037 24075 35071
rect 25053 35037 25087 35071
rect 25145 35037 25179 35071
rect 25329 35037 25363 35071
rect 25421 35037 25455 35071
rect 57897 35037 57931 35071
rect 2329 34969 2363 35003
rect 20913 34969 20947 35003
rect 21557 34969 21591 35003
rect 23949 34969 23983 35003
rect 58173 34969 58207 35003
rect 15853 34901 15887 34935
rect 21189 34901 21223 34935
rect 22753 34901 22787 34935
rect 23489 34901 23523 34935
rect 1869 34629 1903 34663
rect 1685 34561 1719 34595
rect 22017 34561 22051 34595
rect 22293 34561 22327 34595
rect 23673 34561 23707 34595
rect 23857 34561 23891 34595
rect 24409 34561 24443 34595
rect 24961 34561 24995 34595
rect 22753 34493 22787 34527
rect 24593 34493 24627 34527
rect 22109 34425 22143 34459
rect 22569 34153 22603 34187
rect 1869 34085 1903 34119
rect 17693 34017 17727 34051
rect 17233 33949 17267 33983
rect 17417 33949 17451 33983
rect 20177 33949 20211 33983
rect 20545 33949 20579 33983
rect 22293 33949 22327 33983
rect 22385 33949 22419 33983
rect 23121 33949 23155 33983
rect 24593 33949 24627 33983
rect 24686 33949 24720 33983
rect 24869 33949 24903 33983
rect 25099 33949 25133 33983
rect 40141 33949 40175 33983
rect 40289 33949 40323 33983
rect 40417 33949 40451 33983
rect 40606 33949 40640 33983
rect 41337 33949 41371 33983
rect 57989 33949 58023 33983
rect 1685 33881 1719 33915
rect 17325 33881 17359 33915
rect 17555 33881 17589 33915
rect 23489 33881 23523 33915
rect 24961 33881 24995 33915
rect 40509 33881 40543 33915
rect 58357 33881 58391 33915
rect 17049 33813 17083 33847
rect 20085 33813 20119 33847
rect 20269 33813 20303 33847
rect 20361 33813 20395 33847
rect 25237 33813 25271 33847
rect 40785 33813 40819 33847
rect 41521 33813 41555 33847
rect 20269 33609 20303 33643
rect 20361 33609 20395 33643
rect 1869 33541 1903 33575
rect 25329 33541 25363 33575
rect 1685 33473 1719 33507
rect 17785 33473 17819 33507
rect 20177 33473 20211 33507
rect 20545 33473 20579 33507
rect 23581 33473 23615 33507
rect 25053 33473 25087 33507
rect 25201 33473 25235 33507
rect 25421 33473 25455 33507
rect 25559 33473 25593 33507
rect 27353 33473 27387 33507
rect 27537 33473 27571 33507
rect 27905 33473 27939 33507
rect 28457 33473 28491 33507
rect 29193 33473 29227 33507
rect 32781 33473 32815 33507
rect 32965 33473 32999 33507
rect 33065 33473 33099 33507
rect 33195 33473 33229 33507
rect 17969 33405 18003 33439
rect 23949 33405 23983 33439
rect 29469 33405 29503 33439
rect 19993 33337 20027 33371
rect 25697 33269 25731 33303
rect 28641 33269 28675 33303
rect 33333 33269 33367 33303
rect 16773 33065 16807 33099
rect 16957 33065 16991 33099
rect 22385 33065 22419 33099
rect 34069 33065 34103 33099
rect 26157 32997 26191 33031
rect 26801 32997 26835 33031
rect 58173 32929 58207 32963
rect 16589 32861 16623 32895
rect 16773 32861 16807 32895
rect 17601 32861 17635 32895
rect 17877 32861 17911 32895
rect 17969 32861 18003 32895
rect 18429 32861 18463 32895
rect 19625 32861 19659 32895
rect 19791 32861 19825 32895
rect 19902 32839 19936 32873
rect 19994 32861 20028 32895
rect 20269 32861 20303 32895
rect 21005 32861 21039 32895
rect 21189 32861 21223 32895
rect 21557 32861 21591 32895
rect 21741 32861 21775 32895
rect 21925 32861 21959 32895
rect 25513 32861 25547 32895
rect 25606 32861 25640 32895
rect 25978 32861 26012 32895
rect 26709 32861 26743 32895
rect 26985 32861 27019 32895
rect 27445 32861 27479 32895
rect 33057 32861 33091 32895
rect 33149 32861 33183 32895
rect 33333 32861 33367 32895
rect 33425 32861 33459 32895
rect 42901 32861 42935 32895
rect 43049 32861 43083 32895
rect 43366 32861 43400 32895
rect 57897 32861 57931 32895
rect 25789 32793 25823 32827
rect 25881 32793 25915 32827
rect 33977 32793 34011 32827
rect 43177 32793 43211 32827
rect 43269 32793 43303 32827
rect 57069 32793 57103 32827
rect 17509 32725 17543 32759
rect 32873 32725 32907 32759
rect 43545 32725 43579 32759
rect 57161 32725 57195 32759
rect 1869 32453 1903 32487
rect 18245 32453 18279 32487
rect 19809 32453 19843 32487
rect 20453 32453 20487 32487
rect 25421 32453 25455 32487
rect 25973 32453 26007 32487
rect 44925 32453 44959 32487
rect 45017 32453 45051 32487
rect 1685 32385 1719 32419
rect 18705 32385 18739 32419
rect 18797 32385 18831 32419
rect 20269 32385 20303 32419
rect 20361 32385 20395 32419
rect 22201 32385 22235 32419
rect 22293 32385 22327 32419
rect 22385 32385 22419 32419
rect 22569 32385 22603 32419
rect 22661 32385 22695 32419
rect 25605 32385 25639 32419
rect 33057 32385 33091 32419
rect 33517 32385 33551 32419
rect 44741 32385 44775 32419
rect 45114 32385 45148 32419
rect 18337 32317 18371 32351
rect 19257 32317 19291 32351
rect 19901 32317 19935 32351
rect 33149 32317 33183 32351
rect 33885 32249 33919 32283
rect 22017 32181 22051 32215
rect 45293 32181 45327 32215
rect 23121 31977 23155 32011
rect 44649 31977 44683 32011
rect 21373 31909 21407 31943
rect 23581 31909 23615 31943
rect 42901 31909 42935 31943
rect 1869 31841 1903 31875
rect 23213 31841 23247 31875
rect 1685 31773 1719 31807
rect 17417 31773 17451 31807
rect 17877 31773 17911 31807
rect 18061 31773 18095 31807
rect 18889 31773 18923 31807
rect 19901 31773 19935 31807
rect 20453 31773 20487 31807
rect 21557 31773 21591 31807
rect 21925 31773 21959 31807
rect 22017 31773 22051 31807
rect 23121 31773 23155 31807
rect 23397 31773 23431 31807
rect 25145 31773 25179 31807
rect 32873 31773 32907 31807
rect 42257 31773 42291 31807
rect 42405 31773 42439 31807
rect 42625 31773 42659 31807
rect 42722 31773 42756 31807
rect 44005 31773 44039 31807
rect 44098 31773 44132 31807
rect 44281 31773 44315 31807
rect 44470 31773 44504 31807
rect 57897 31773 57931 31807
rect 58173 31773 58207 31807
rect 25697 31705 25731 31739
rect 33701 31705 33735 31739
rect 42533 31705 42567 31739
rect 44373 31705 44407 31739
rect 17325 31637 17359 31671
rect 19257 31365 19291 31399
rect 25145 31365 25179 31399
rect 25881 31365 25915 31399
rect 35265 31365 35299 31399
rect 1685 31297 1719 31331
rect 18153 31297 18187 31331
rect 18521 31297 18555 31331
rect 19073 31297 19107 31331
rect 19625 31297 19659 31331
rect 20269 31297 20303 31331
rect 22293 31297 22327 31331
rect 24777 31297 24811 31331
rect 24925 31297 24959 31331
rect 25053 31297 25087 31331
rect 25283 31297 25317 31331
rect 26065 31297 26099 31331
rect 33793 31297 33827 31331
rect 34069 31297 34103 31331
rect 34989 31297 35023 31331
rect 35137 31297 35171 31331
rect 35357 31297 35391 31331
rect 35454 31297 35488 31331
rect 36369 31297 36403 31331
rect 20545 31229 20579 31263
rect 22569 31229 22603 31263
rect 26341 31229 26375 31263
rect 34253 31229 34287 31263
rect 36553 31229 36587 31263
rect 33885 31161 33919 31195
rect 35633 31161 35667 31195
rect 1777 31093 1811 31127
rect 25421 31093 25455 31127
rect 38301 30889 38335 30923
rect 23581 30821 23615 30855
rect 17509 30753 17543 30787
rect 21557 30753 21591 30787
rect 30481 30753 30515 30787
rect 17969 30685 18003 30719
rect 18061 30685 18095 30719
rect 18521 30685 18555 30719
rect 19717 30685 19751 30719
rect 19993 30685 20027 30719
rect 20453 30685 20487 30719
rect 20729 30685 20763 30719
rect 22017 30685 22051 30719
rect 22201 30685 22235 30719
rect 22385 30685 22419 30719
rect 23029 30685 23063 30719
rect 23305 30685 23339 30719
rect 23397 30685 23431 30719
rect 24593 30685 24627 30719
rect 24777 30685 24811 30719
rect 30389 30685 30423 30719
rect 30757 30685 30791 30719
rect 30941 30685 30975 30719
rect 35817 30685 35851 30719
rect 35910 30685 35944 30719
rect 36093 30685 36127 30719
rect 36282 30685 36316 30719
rect 36921 30685 36955 30719
rect 37014 30685 37048 30719
rect 37197 30685 37231 30719
rect 37289 30685 37323 30719
rect 37427 30685 37461 30719
rect 38209 30685 38243 30719
rect 57989 30685 58023 30719
rect 1685 30617 1719 30651
rect 17601 30617 17635 30651
rect 23213 30617 23247 30651
rect 29745 30617 29779 30651
rect 36185 30617 36219 30651
rect 38025 30617 38059 30651
rect 1777 30549 1811 30583
rect 20637 30549 20671 30583
rect 24869 30549 24903 30583
rect 36461 30549 36495 30583
rect 37565 30549 37599 30583
rect 58081 30549 58115 30583
rect 19625 30345 19659 30379
rect 17785 30277 17819 30311
rect 17877 30277 17911 30311
rect 20637 30277 20671 30311
rect 22569 30277 22603 30311
rect 37473 30277 37507 30311
rect 18245 30209 18279 30243
rect 18337 30209 18371 30243
rect 19349 30209 19383 30243
rect 20269 30209 20303 30243
rect 22109 30209 22143 30243
rect 37657 30209 37691 30243
rect 18797 30141 18831 30175
rect 22017 30141 22051 30175
rect 37749 30005 37783 30039
rect 21741 29801 21775 29835
rect 35449 29801 35483 29835
rect 43821 29801 43855 29835
rect 58173 29665 58207 29699
rect 1593 29597 1627 29631
rect 15209 29597 15243 29631
rect 15363 29597 15397 29631
rect 19533 29597 19567 29631
rect 19901 29597 19935 29631
rect 20453 29597 20487 29631
rect 21005 29597 21039 29631
rect 34897 29597 34931 29631
rect 35173 29597 35207 29631
rect 35265 29597 35299 29631
rect 43177 29597 43211 29631
rect 43325 29597 43359 29631
rect 43453 29597 43487 29631
rect 43683 29597 43717 29631
rect 57897 29597 57931 29631
rect 1869 29529 1903 29563
rect 15577 29529 15611 29563
rect 21649 29529 21683 29563
rect 35081 29529 35115 29563
rect 43545 29529 43579 29563
rect 57069 29529 57103 29563
rect 19533 29461 19567 29495
rect 57161 29461 57195 29495
rect 19625 29257 19659 29291
rect 24409 29257 24443 29291
rect 18613 29189 18647 29223
rect 1593 29121 1627 29155
rect 18705 29121 18739 29155
rect 18797 29121 18831 29155
rect 19441 29121 19475 29155
rect 20637 29121 20671 29155
rect 23765 29121 23799 29155
rect 24133 29121 24167 29155
rect 24225 29121 24259 29155
rect 1777 29053 1811 29087
rect 18061 29053 18095 29087
rect 18245 29053 18279 29087
rect 20821 28985 20855 29019
rect 2881 28645 2915 28679
rect 1593 28509 1627 28543
rect 2513 28509 2547 28543
rect 2667 28509 2701 28543
rect 57897 28509 57931 28543
rect 1869 28441 1903 28475
rect 58173 28441 58207 28475
rect 2881 28169 2915 28203
rect 2237 28101 2271 28135
rect 1409 28033 1443 28067
rect 2513 28033 2547 28067
rect 2667 28033 2701 28067
rect 1593 27965 1627 27999
rect 2237 27625 2271 27659
rect 18061 27489 18095 27523
rect 2053 27421 2087 27455
rect 2207 27421 2241 27455
rect 18153 27421 18187 27455
rect 18521 27421 18555 27455
rect 57989 27421 58023 27455
rect 18613 27353 18647 27387
rect 18705 27353 18739 27387
rect 58081 27285 58115 27319
rect 2881 27013 2915 27047
rect 18061 27013 18095 27047
rect 1593 26945 1627 26979
rect 2513 26945 2547 26979
rect 2667 26945 2701 26979
rect 17969 26945 18003 26979
rect 18429 26945 18463 26979
rect 18521 26945 18555 26979
rect 18981 26945 19015 26979
rect 19993 26945 20027 26979
rect 20085 26945 20119 26979
rect 20545 26945 20579 26979
rect 1777 26877 1811 26911
rect 19533 26877 19567 26911
rect 19625 26877 19659 26911
rect 2881 26401 2915 26435
rect 18613 26401 18647 26435
rect 20177 26401 20211 26435
rect 26249 26401 26283 26435
rect 58173 26401 58207 26435
rect 1593 26333 1627 26367
rect 2513 26333 2547 26367
rect 2606 26333 2640 26367
rect 18245 26333 18279 26367
rect 19441 26333 19475 26367
rect 25421 26333 25455 26367
rect 26065 26333 26099 26367
rect 27169 26333 27203 26367
rect 27261 26333 27295 26367
rect 57897 26333 57931 26367
rect 1869 26265 1903 26299
rect 26157 26265 26191 26299
rect 27445 26265 27479 26299
rect 25697 26197 25731 26231
rect 28273 25993 28307 26027
rect 28365 25925 28399 25959
rect 29285 25925 29319 25959
rect 1593 25857 1627 25891
rect 19901 25857 19935 25891
rect 20545 25857 20579 25891
rect 20637 25857 20671 25891
rect 25973 25857 26007 25891
rect 29469 25857 29503 25891
rect 58081 25857 58115 25891
rect 1777 25789 1811 25823
rect 20729 25789 20763 25823
rect 26065 25789 26099 25823
rect 26249 25789 26283 25823
rect 28273 25789 28307 25823
rect 25329 25721 25363 25755
rect 20177 25653 20211 25687
rect 25605 25653 25639 25687
rect 27813 25653 27847 25687
rect 29653 25653 29687 25687
rect 58265 25653 58299 25687
rect 2697 25449 2731 25483
rect 16497 25313 16531 25347
rect 21925 25313 21959 25347
rect 29101 25313 29135 25347
rect 56701 25313 56735 25347
rect 1593 25245 1627 25279
rect 2513 25245 2547 25279
rect 2667 25245 2701 25279
rect 16129 25245 16163 25279
rect 19349 25245 19383 25279
rect 21097 25245 21131 25279
rect 21741 25245 21775 25279
rect 24961 25245 24995 25279
rect 27169 25245 27203 25279
rect 29009 25245 29043 25279
rect 29193 25245 29227 25279
rect 29745 25245 29779 25279
rect 55873 25245 55907 25279
rect 56057 25245 56091 25279
rect 56885 25245 56919 25279
rect 57897 25245 57931 25279
rect 1869 25177 1903 25211
rect 19616 25177 19650 25211
rect 21833 25177 21867 25211
rect 25228 25177 25262 25211
rect 27414 25177 27448 25211
rect 29929 25177 29963 25211
rect 58173 25177 58207 25211
rect 20729 25109 20763 25143
rect 21373 25109 21407 25143
rect 26341 25109 26375 25143
rect 28549 25109 28583 25143
rect 30113 25109 30147 25143
rect 56241 25109 56275 25143
rect 57069 25109 57103 25143
rect 16221 24905 16255 24939
rect 56057 24905 56091 24939
rect 57069 24905 57103 24939
rect 31401 24837 31435 24871
rect 31769 24837 31803 24871
rect 56793 24837 56827 24871
rect 15853 24769 15887 24803
rect 16007 24769 16041 24803
rect 19349 24769 19383 24803
rect 19533 24769 19567 24803
rect 19625 24769 19659 24803
rect 20085 24769 20119 24803
rect 20352 24769 20386 24803
rect 22477 24769 22511 24803
rect 23581 24769 23615 24803
rect 26433 24769 26467 24803
rect 26617 24769 26651 24803
rect 27977 24769 28011 24803
rect 29828 24769 29862 24803
rect 31585 24769 31619 24803
rect 32597 24769 32631 24803
rect 32689 24769 32723 24803
rect 32781 24769 32815 24803
rect 32965 24769 32999 24803
rect 45477 24769 45511 24803
rect 45845 24769 45879 24803
rect 54309 24769 54343 24803
rect 55505 24769 55539 24803
rect 55689 24769 55723 24803
rect 55781 24769 55815 24803
rect 55873 24769 55907 24803
rect 56517 24769 56551 24803
rect 56701 24769 56735 24803
rect 56885 24769 56919 24803
rect 58081 24769 58115 24803
rect 22293 24701 22327 24735
rect 27721 24701 27755 24735
rect 29561 24701 29595 24735
rect 45385 24701 45419 24735
rect 45937 24701 45971 24735
rect 54585 24701 54619 24735
rect 33241 24633 33275 24667
rect 19349 24565 19383 24599
rect 21465 24565 21499 24599
rect 22661 24565 22695 24599
rect 24777 24565 24811 24599
rect 26525 24565 26559 24599
rect 29101 24565 29135 24599
rect 30941 24565 30975 24599
rect 32321 24565 32355 24599
rect 44925 24565 44959 24599
rect 58265 24565 58299 24599
rect 23029 24293 23063 24327
rect 44649 24293 44683 24327
rect 53941 24293 53975 24327
rect 57437 24293 57471 24327
rect 17601 24225 17635 24259
rect 19533 24225 19567 24259
rect 24593 24225 24627 24259
rect 52101 24225 52135 24259
rect 54493 24225 54527 24259
rect 1593 24157 1627 24191
rect 17509 24157 17543 24191
rect 17877 24157 17911 24191
rect 18061 24157 18095 24191
rect 19800 24157 19834 24191
rect 21373 24157 21407 24191
rect 21557 24157 21591 24191
rect 23581 24157 23615 24191
rect 24860 24157 24894 24191
rect 26433 24157 26467 24191
rect 30021 24157 30055 24191
rect 31953 24157 31987 24191
rect 43269 24157 43303 24191
rect 50353 24157 50387 24191
rect 50537 24157 50571 24191
rect 51641 24157 51675 24191
rect 51943 24157 51977 24191
rect 52561 24157 52595 24191
rect 54677 24157 54711 24191
rect 56057 24157 56091 24191
rect 56324 24157 56358 24191
rect 57897 24157 57931 24191
rect 1869 24089 1903 24123
rect 16865 24089 16899 24123
rect 23397 24089 23431 24123
rect 30288 24089 30322 24123
rect 32220 24089 32254 24123
rect 43536 24089 43570 24123
rect 51733 24089 51767 24123
rect 51825 24089 51859 24123
rect 52828 24089 52862 24123
rect 58173 24089 58207 24123
rect 20913 24021 20947 24055
rect 21741 24021 21775 24055
rect 23213 24021 23247 24055
rect 23305 24021 23339 24055
rect 25973 24021 26007 24055
rect 27629 24021 27663 24055
rect 31401 24021 31435 24055
rect 33333 24021 33367 24055
rect 50721 24021 50755 24055
rect 51457 24021 51491 24055
rect 54861 24021 54895 24055
rect 20177 23817 20211 23851
rect 20637 23817 20671 23851
rect 22293 23817 22327 23851
rect 27261 23817 27295 23851
rect 29561 23817 29595 23851
rect 31125 23817 31159 23851
rect 32873 23817 32907 23851
rect 40417 23817 40451 23851
rect 57529 23817 57563 23851
rect 19165 23749 19199 23783
rect 20545 23749 20579 23783
rect 32689 23749 32723 23783
rect 41981 23749 42015 23783
rect 42870 23749 42904 23783
rect 1593 23681 1627 23715
rect 13553 23681 13587 23715
rect 13707 23681 13741 23715
rect 15577 23681 15611 23715
rect 15731 23681 15765 23715
rect 18153 23681 18187 23715
rect 22234 23681 22268 23715
rect 22753 23681 22787 23715
rect 23305 23681 23339 23715
rect 23949 23681 23983 23715
rect 27537 23681 27571 23715
rect 27629 23681 27663 23715
rect 27721 23681 27755 23715
rect 27905 23681 27939 23715
rect 28365 23681 28399 23715
rect 31401 23681 31435 23715
rect 31490 23681 31524 23715
rect 31585 23681 31619 23715
rect 31769 23681 31803 23715
rect 33968 23681 34002 23715
rect 36461 23681 36495 23715
rect 36645 23681 36679 23715
rect 38393 23681 38427 23715
rect 39293 23681 39327 23715
rect 41889 23681 41923 23715
rect 42073 23681 42107 23715
rect 44465 23681 44499 23715
rect 44649 23681 44683 23715
rect 50353 23681 50387 23715
rect 50620 23681 50654 23715
rect 53113 23681 53147 23715
rect 53297 23681 53331 23715
rect 53757 23681 53791 23715
rect 54024 23681 54058 23715
rect 56149 23681 56183 23715
rect 56416 23681 56450 23715
rect 1777 23613 1811 23647
rect 13921 23613 13955 23647
rect 20729 23613 20763 23647
rect 22661 23613 22695 23647
rect 32965 23613 32999 23647
rect 33701 23613 33735 23647
rect 38209 23613 38243 23647
rect 39037 23613 39071 23647
rect 42625 23613 42659 23647
rect 52929 23613 52963 23647
rect 15945 23545 15979 23579
rect 25145 23545 25179 23579
rect 28273 23545 28307 23579
rect 35081 23545 35115 23579
rect 51733 23545 51767 23579
rect 22109 23477 22143 23511
rect 23397 23477 23431 23511
rect 32413 23477 32447 23511
rect 36829 23477 36863 23511
rect 38577 23477 38611 23511
rect 44005 23477 44039 23511
rect 44465 23477 44499 23511
rect 55137 23477 55171 23511
rect 19809 23273 19843 23307
rect 19993 23273 20027 23307
rect 25605 23273 25639 23307
rect 28089 23273 28123 23307
rect 29745 23273 29779 23307
rect 35357 23273 35391 23307
rect 38485 23273 38519 23307
rect 41981 23273 42015 23307
rect 42533 23273 42567 23307
rect 43269 23273 43303 23307
rect 50905 23273 50939 23307
rect 53757 23273 53791 23307
rect 58265 23273 58299 23307
rect 20453 23205 20487 23239
rect 24961 23205 24995 23239
rect 37933 23205 37967 23239
rect 18429 23137 18463 23171
rect 18889 23137 18923 23171
rect 24685 23137 24719 23171
rect 39129 23137 39163 23171
rect 40693 23137 40727 23171
rect 54401 23137 54435 23171
rect 56241 23137 56275 23171
rect 56885 23137 56919 23171
rect 1593 23069 1627 23103
rect 15945 23069 15979 23103
rect 18521 23069 18555 23103
rect 20637 23069 20671 23103
rect 21005 23069 21039 23103
rect 21741 23069 21775 23103
rect 24593 23069 24627 23103
rect 25329 23069 25363 23103
rect 25835 23069 25869 23103
rect 25973 23069 26007 23103
rect 26065 23069 26099 23103
rect 26249 23069 26283 23103
rect 26709 23069 26743 23103
rect 30021 23069 30055 23103
rect 30110 23069 30144 23103
rect 30210 23069 30244 23103
rect 30389 23069 30423 23103
rect 31033 23069 31067 23103
rect 35909 23069 35943 23103
rect 36553 23069 36587 23103
rect 38669 23069 38703 23103
rect 38991 23069 39025 23103
rect 40233 23063 40267 23097
rect 40325 23069 40359 23103
rect 42162 23069 42196 23103
rect 42625 23069 42659 23103
rect 43394 23069 43428 23103
rect 43821 23069 43855 23103
rect 43913 23069 43947 23103
rect 47961 23069 47995 23103
rect 50353 23069 50387 23103
rect 50721 23069 50755 23103
rect 53941 23069 53975 23103
rect 54125 23069 54159 23103
rect 54243 23069 54277 23103
rect 56149 23069 56183 23103
rect 56338 23069 56372 23103
rect 57152 23069 57186 23103
rect 1869 23001 1903 23035
rect 16212 23001 16246 23035
rect 19625 23001 19659 23035
rect 20729 23001 20763 23035
rect 33793 23001 33827 23035
rect 33977 23001 34011 23035
rect 35633 23001 35667 23035
rect 35817 23001 35851 23035
rect 36798 23001 36832 23035
rect 38761 23001 38795 23035
rect 38853 23001 38887 23035
rect 40049 23001 40083 23035
rect 40417 23001 40451 23035
rect 40535 23001 40569 23035
rect 48237 23001 48271 23035
rect 50537 23001 50571 23035
rect 50629 23001 50663 23035
rect 54033 23001 54067 23035
rect 55965 23001 55999 23035
rect 56241 23001 56275 23035
rect 17325 22933 17359 22967
rect 19825 22933 19859 22967
rect 20821 22933 20855 22967
rect 22937 22933 22971 22967
rect 32229 22933 32263 22967
rect 34161 22933 34195 22967
rect 42165 22933 42199 22967
rect 43453 22933 43487 22967
rect 53389 22933 53423 22967
rect 17509 22729 17543 22763
rect 23857 22729 23891 22763
rect 25513 22729 25547 22763
rect 35081 22729 35115 22763
rect 36277 22729 36311 22763
rect 37841 22729 37875 22763
rect 40325 22729 40359 22763
rect 45845 22729 45879 22763
rect 49157 22729 49191 22763
rect 21189 22661 21223 22695
rect 22744 22661 22778 22695
rect 37657 22661 37691 22695
rect 1593 22593 1627 22627
rect 17049 22593 17083 22627
rect 17417 22593 17451 22627
rect 17785 22593 17819 22627
rect 18429 22593 18463 22627
rect 21373 22593 21407 22627
rect 21465 22593 21499 22627
rect 24317 22593 24351 22627
rect 27445 22593 27479 22627
rect 27721 22593 27755 22627
rect 27997 22593 28031 22627
rect 28365 22593 28399 22627
rect 29469 22593 29503 22627
rect 32321 22593 32355 22627
rect 35311 22593 35345 22627
rect 35449 22593 35483 22627
rect 35541 22593 35575 22627
rect 35725 22593 35759 22627
rect 36533 22593 36567 22627
rect 36645 22593 36679 22627
rect 36758 22599 36792 22633
rect 36921 22593 36955 22627
rect 37473 22593 37507 22627
rect 39201 22593 39235 22627
rect 43821 22593 43855 22627
rect 44005 22593 44039 22627
rect 44465 22593 44499 22627
rect 44732 22593 44766 22627
rect 48044 22593 48078 22627
rect 56517 22593 56551 22627
rect 56701 22593 56735 22627
rect 58081 22593 58115 22627
rect 1777 22525 1811 22559
rect 22477 22525 22511 22559
rect 27629 22525 27663 22559
rect 38945 22525 38979 22559
rect 47777 22525 47811 22559
rect 56517 22457 56551 22491
rect 19625 22389 19659 22423
rect 21189 22389 21223 22423
rect 30665 22389 30699 22423
rect 33517 22389 33551 22423
rect 43821 22389 43855 22423
rect 58265 22389 58299 22423
rect 13553 22185 13587 22219
rect 34161 22117 34195 22151
rect 37105 22117 37139 22151
rect 44373 22117 44407 22151
rect 45201 22117 45235 22151
rect 45753 22117 45787 22151
rect 46121 22117 46155 22151
rect 34897 22049 34931 22083
rect 37289 22049 37323 22083
rect 39129 22049 39163 22083
rect 48881 22049 48915 22083
rect 13369 21981 13403 22015
rect 13523 21981 13557 22015
rect 14381 21981 14415 22015
rect 16589 21981 16623 22015
rect 19441 21981 19475 22015
rect 21741 21981 21775 22015
rect 24593 21981 24627 22015
rect 26893 21981 26927 22015
rect 30067 21981 30101 22015
rect 30205 21981 30239 22015
rect 30318 21981 30352 22015
rect 30481 21981 30515 22015
rect 31033 21981 31067 22015
rect 33966 21981 34000 22015
rect 35173 21981 35207 22015
rect 37013 21981 37047 22015
rect 37933 21981 37967 22015
rect 38117 21981 38151 22015
rect 38853 21981 38887 22015
rect 38945 21981 38979 22015
rect 40049 21981 40083 22015
rect 40325 21981 40359 22015
rect 43177 21981 43211 22015
rect 43361 21981 43395 22015
rect 44002 21981 44036 22015
rect 44465 21981 44499 22015
rect 45382 21981 45416 22015
rect 45845 21981 45879 22015
rect 47501 21981 47535 22015
rect 47869 21981 47903 22015
rect 48513 21981 48547 22015
rect 48697 21981 48731 22015
rect 57897 21981 57931 22015
rect 14933 21913 14967 21947
rect 19708 21913 19742 21947
rect 24860 21913 24894 21947
rect 33793 21913 33827 21947
rect 37289 21913 37323 21947
rect 38301 21913 38335 21947
rect 43269 21913 43303 21947
rect 47685 21913 47719 21947
rect 47777 21913 47811 21947
rect 58173 21913 58207 21947
rect 17785 21845 17819 21879
rect 20821 21845 20855 21879
rect 22937 21845 22971 21879
rect 25973 21845 26007 21879
rect 28089 21845 28123 21879
rect 29837 21845 29871 21879
rect 32229 21845 32263 21879
rect 36277 21845 36311 21879
rect 43821 21845 43855 21879
rect 44005 21845 44039 21879
rect 45385 21845 45419 21879
rect 48053 21845 48087 21879
rect 14197 21641 14231 21675
rect 20361 21641 20395 21675
rect 25513 21641 25547 21675
rect 27169 21641 27203 21675
rect 27353 21641 27387 21675
rect 31769 21641 31803 21675
rect 35449 21641 35483 21675
rect 22652 21573 22686 21607
rect 32566 21573 32600 21607
rect 34805 21573 34839 21607
rect 1685 21505 1719 21539
rect 13921 21505 13955 21539
rect 15485 21505 15519 21539
rect 15669 21505 15703 21539
rect 16129 21505 16163 21539
rect 16313 21505 16347 21539
rect 17233 21505 17267 21539
rect 17500 21505 17534 21539
rect 19165 21505 19199 21539
rect 22385 21505 22419 21539
rect 24317 21505 24351 21539
rect 27350 21505 27384 21539
rect 27813 21505 27847 21539
rect 28641 21505 28675 21539
rect 31401 21505 31435 21539
rect 31585 21505 31619 21539
rect 34621 21505 34655 21539
rect 35725 21505 35759 21539
rect 35817 21505 35851 21539
rect 35909 21505 35943 21539
rect 36093 21505 36127 21539
rect 36553 21505 36587 21539
rect 36737 21505 36771 21539
rect 37841 21505 37875 21539
rect 40417 21505 40451 21539
rect 40673 21505 40707 21539
rect 44272 21505 44306 21539
rect 50261 21505 50295 21539
rect 56425 21505 56459 21539
rect 56609 21505 56643 21539
rect 57161 21505 57195 21539
rect 1869 21437 1903 21471
rect 32321 21437 32355 21471
rect 34897 21437 34931 21471
rect 37933 21437 37967 21471
rect 38025 21437 38059 21471
rect 44005 21437 44039 21471
rect 50077 21437 50111 21471
rect 15577 21369 15611 21403
rect 33701 21369 33735 21403
rect 16129 21301 16163 21335
rect 18613 21301 18647 21335
rect 23765 21301 23799 21335
rect 27721 21301 27755 21335
rect 29837 21301 29871 21335
rect 34345 21301 34379 21335
rect 36921 21301 36955 21335
rect 37473 21301 37507 21335
rect 41797 21301 41831 21335
rect 45385 21301 45419 21335
rect 50445 21301 50479 21335
rect 56425 21301 56459 21335
rect 57253 21301 57287 21335
rect 17785 21097 17819 21131
rect 29837 21097 29871 21131
rect 40969 21097 41003 21131
rect 48145 21097 48179 21131
rect 51733 21097 51767 21131
rect 58265 21097 58299 21131
rect 16037 21029 16071 21063
rect 20821 21029 20855 21063
rect 26801 21029 26835 21063
rect 28365 21029 28399 21063
rect 14473 20961 14507 20995
rect 24685 20961 24719 20995
rect 31493 20961 31527 20995
rect 33885 20961 33919 20995
rect 43361 20961 43395 20995
rect 56241 20961 56275 20995
rect 56885 20961 56919 20995
rect 1593 20893 1627 20927
rect 14749 20893 14783 20927
rect 16589 20893 16623 20927
rect 19441 20893 19475 20927
rect 21741 20893 21775 20927
rect 24777 20893 24811 20927
rect 25605 20893 25639 20927
rect 28549 20893 28583 20927
rect 28825 20893 28859 20927
rect 29745 20893 29779 20927
rect 30389 20893 30423 20927
rect 35081 20893 35115 20927
rect 36507 20893 36541 20927
rect 36645 20893 36679 20927
rect 36758 20890 36792 20924
rect 36921 20893 36955 20927
rect 38209 20893 38243 20927
rect 40598 20893 40632 20927
rect 41073 20893 41107 20927
rect 50353 20893 50387 20927
rect 56338 20893 56372 20927
rect 57141 20893 57175 20927
rect 1869 20825 1903 20859
rect 19708 20825 19742 20859
rect 28733 20825 28767 20859
rect 33149 20825 33183 20859
rect 34897 20825 34931 20859
rect 35449 20825 35483 20859
rect 37381 20825 37415 20859
rect 37565 20825 37599 20859
rect 41613 20825 41647 20859
rect 46857 20825 46891 20859
rect 50598 20825 50632 20859
rect 55965 20825 55999 20859
rect 56149 20825 56183 20859
rect 56241 20825 56275 20859
rect 22937 20757 22971 20791
rect 25145 20757 25179 20791
rect 36277 20757 36311 20791
rect 37749 20757 37783 20791
rect 38393 20757 38427 20791
rect 40417 20757 40451 20791
rect 40601 20757 40635 20791
rect 17417 20553 17451 20587
rect 23765 20553 23799 20587
rect 29837 20553 29871 20587
rect 40417 20553 40451 20587
rect 50353 20553 50387 20587
rect 22652 20485 22686 20519
rect 27445 20485 27479 20519
rect 36185 20485 36219 20519
rect 37749 20485 37783 20519
rect 1593 20417 1627 20451
rect 15945 20417 15979 20451
rect 17049 20417 17083 20451
rect 18337 20417 18371 20451
rect 18429 20417 18463 20451
rect 19165 20417 19199 20451
rect 22385 20417 22419 20451
rect 24317 20417 24351 20451
rect 27353 20417 27387 20451
rect 27537 20417 27571 20451
rect 28641 20417 28675 20451
rect 31401 20417 31435 20451
rect 31677 20417 31711 20451
rect 32321 20417 32355 20451
rect 36001 20417 36035 20451
rect 37473 20417 37507 20451
rect 38853 20417 38887 20451
rect 40325 20417 40359 20451
rect 40509 20417 40543 20451
rect 45385 20417 45419 20451
rect 45569 20417 45603 20451
rect 45661 20417 45695 20451
rect 45753 20417 45787 20451
rect 49801 20417 49835 20451
rect 49985 20417 50019 20451
rect 50077 20417 50111 20451
rect 50169 20417 50203 20451
rect 52929 20417 52963 20451
rect 53196 20417 53230 20451
rect 1777 20349 1811 20383
rect 16037 20349 16071 20383
rect 16957 20349 16991 20383
rect 18521 20349 18555 20383
rect 18613 20349 18647 20383
rect 20729 20349 20763 20383
rect 36277 20349 36311 20383
rect 39037 20349 39071 20383
rect 25513 20281 25547 20315
rect 27169 20281 27203 20315
rect 27721 20281 27755 20315
rect 31677 20281 31711 20315
rect 35725 20281 35759 20315
rect 16313 20213 16347 20247
rect 18153 20213 18187 20247
rect 33517 20213 33551 20247
rect 45937 20213 45971 20247
rect 54309 20213 54343 20247
rect 17141 20009 17175 20043
rect 21005 20009 21039 20043
rect 24685 20009 24719 20043
rect 26525 20009 26559 20043
rect 28549 20009 28583 20043
rect 29101 20009 29135 20043
rect 40233 20009 40267 20043
rect 32689 19941 32723 19975
rect 22661 19873 22695 19907
rect 29193 19873 29227 19907
rect 30481 19873 30515 19907
rect 36001 19873 36035 19907
rect 39037 19873 39071 19907
rect 41521 19873 41555 19907
rect 45937 19873 45971 19907
rect 46305 19873 46339 19907
rect 52653 19873 52687 19907
rect 57345 19873 57379 19907
rect 58173 19873 58207 19907
rect 1593 19805 1627 19839
rect 15945 19805 15979 19839
rect 18705 19805 18739 19839
rect 18889 19805 18923 19839
rect 19809 19805 19843 19839
rect 24685 19805 24719 19839
rect 24869 19805 24903 19839
rect 25329 19805 25363 19839
rect 28674 19805 28708 19839
rect 30389 19805 30423 19839
rect 30757 19805 30791 19839
rect 30941 19805 30975 19839
rect 31493 19805 31527 19839
rect 34897 19805 34931 19839
rect 37657 19805 37691 19839
rect 37933 19805 37967 19839
rect 40141 19805 40175 19839
rect 41061 19805 41095 19839
rect 41245 19805 41279 19839
rect 45845 19805 45879 19839
rect 46213 19805 46247 19839
rect 52193 19805 52227 19839
rect 57897 19805 57931 19839
rect 1869 19737 1903 19771
rect 22928 19737 22962 19771
rect 29745 19737 29779 19771
rect 45201 19737 45235 19771
rect 52285 19737 52319 19771
rect 52377 19737 52411 19771
rect 52515 19737 52549 19771
rect 57069 19737 57103 19771
rect 18797 19669 18831 19703
rect 24041 19669 24075 19703
rect 28733 19669 28767 19703
rect 52009 19669 52043 19703
rect 15117 19465 15151 19499
rect 18337 19465 18371 19499
rect 25513 19465 25547 19499
rect 36461 19465 36495 19499
rect 37473 19465 37507 19499
rect 45385 19465 45419 19499
rect 52377 19465 52411 19499
rect 56977 19465 57011 19499
rect 18061 19397 18095 19431
rect 23857 19397 23891 19431
rect 28646 19397 28680 19431
rect 17417 19329 17451 19363
rect 17601 19329 17635 19363
rect 18245 19329 18279 19363
rect 18429 19329 18463 19363
rect 19165 19329 19199 19363
rect 24317 19329 24351 19363
rect 27354 19329 27388 19363
rect 28365 19329 28399 19363
rect 28549 19329 28583 19363
rect 28779 19329 28813 19363
rect 29469 19329 29503 19363
rect 32321 19329 32355 19363
rect 35081 19329 35115 19363
rect 35348 19329 35382 19363
rect 37749 19329 37783 19363
rect 37841 19329 37875 19363
rect 37933 19329 37967 19363
rect 38117 19329 38151 19363
rect 38761 19329 38795 19363
rect 39017 19329 39051 19363
rect 44005 19329 44039 19363
rect 44272 19329 44306 19363
rect 52193 19329 52227 19363
rect 56793 19329 56827 19363
rect 57069 19329 57103 19363
rect 15301 19261 15335 19295
rect 15393 19261 15427 19295
rect 15485 19261 15519 19295
rect 15577 19261 15611 19295
rect 17509 19261 17543 19295
rect 22201 19261 22235 19295
rect 22477 19261 22511 19295
rect 27445 19261 27479 19295
rect 27537 19261 27571 19295
rect 27629 19261 27663 19295
rect 30665 19261 30699 19295
rect 33425 19261 33459 19295
rect 52009 19261 52043 19295
rect 28917 19193 28951 19227
rect 18613 19125 18647 19159
rect 21373 19125 21407 19159
rect 27169 19125 27203 19159
rect 40141 19125 40175 19159
rect 56793 19125 56827 19159
rect 10793 18921 10827 18955
rect 35449 18921 35483 18955
rect 37933 18921 37967 18955
rect 38393 18921 38427 18955
rect 58265 18921 58299 18955
rect 44373 18853 44407 18887
rect 11069 18785 11103 18819
rect 11161 18785 11195 18819
rect 18613 18785 18647 18819
rect 18889 18785 18923 18819
rect 19809 18785 19843 18819
rect 30757 18785 30791 18819
rect 43085 18785 43119 18819
rect 1593 18717 1627 18751
rect 10977 18717 11011 18751
rect 11253 18717 11287 18751
rect 16037 18717 16071 18751
rect 16191 18717 16225 18751
rect 16957 18717 16991 18751
rect 17325 18717 17359 18751
rect 17509 18717 17543 18751
rect 18521 18717 18555 18751
rect 21741 18717 21775 18751
rect 24593 18717 24627 18751
rect 24777 18717 24811 18751
rect 25237 18717 25271 18751
rect 28273 18717 28307 18751
rect 28365 18717 28399 18751
rect 28457 18717 28491 18751
rect 28641 18717 28675 18751
rect 30573 18717 30607 18751
rect 30849 18717 30883 18751
rect 31125 18717 31159 18751
rect 31585 18717 31619 18751
rect 32505 18717 32539 18751
rect 32597 18717 32631 18751
rect 32781 18717 32815 18751
rect 32873 18717 32907 18751
rect 33425 18717 33459 18751
rect 33609 18717 33643 18751
rect 33700 18717 33734 18751
rect 33885 18717 33919 18751
rect 33977 18717 34011 18751
rect 35725 18717 35759 18751
rect 35817 18717 35851 18751
rect 35909 18717 35943 18751
rect 36093 18717 36127 18751
rect 36553 18717 36587 18751
rect 38669 18717 38703 18751
rect 38758 18717 38792 18751
rect 38874 18711 38908 18745
rect 39037 18717 39071 18751
rect 42993 18717 43027 18751
rect 43177 18717 43211 18751
rect 44002 18717 44036 18751
rect 44465 18717 44499 18751
rect 56885 18717 56919 18751
rect 57141 18717 57175 18751
rect 1869 18649 1903 18683
rect 16405 18649 16439 18683
rect 20076 18649 20110 18683
rect 36798 18649 36832 18683
rect 17049 18581 17083 18615
rect 21189 18581 21223 18615
rect 22937 18581 22971 18615
rect 24777 18581 24811 18615
rect 26433 18581 26467 18615
rect 27997 18581 28031 18615
rect 32321 18581 32355 18615
rect 43453 18581 43487 18615
rect 43821 18581 43855 18615
rect 44005 18581 44039 18615
rect 10517 18377 10551 18411
rect 16221 18377 16255 18411
rect 20361 18377 20395 18411
rect 25513 18377 25547 18411
rect 32781 18377 32815 18411
rect 37933 18377 37967 18411
rect 56977 18377 57011 18411
rect 58173 18377 58207 18411
rect 10057 18309 10091 18343
rect 22652 18309 22686 18343
rect 32413 18309 32447 18343
rect 32597 18309 32631 18343
rect 34621 18309 34655 18343
rect 39221 18309 39255 18343
rect 41889 18309 41923 18343
rect 42870 18309 42904 18343
rect 1593 18241 1627 18275
rect 15209 18241 15243 18275
rect 15853 18241 15887 18275
rect 17141 18241 17175 18275
rect 17233 18241 17267 18275
rect 17417 18241 17451 18275
rect 18337 18241 18371 18275
rect 18613 18241 18647 18275
rect 19165 18241 19199 18275
rect 22385 18241 22419 18275
rect 24317 18241 24351 18275
rect 27169 18241 27203 18275
rect 27353 18241 27387 18275
rect 27813 18241 27847 18275
rect 28080 18241 28114 18275
rect 30389 18241 30423 18275
rect 30849 18241 30883 18275
rect 31125 18241 31159 18275
rect 31493 18241 31527 18275
rect 33517 18241 33551 18275
rect 33609 18241 33643 18275
rect 33793 18241 33827 18275
rect 33885 18241 33919 18275
rect 34345 18241 34379 18275
rect 34438 18241 34472 18275
rect 34713 18241 34747 18275
rect 34851 18241 34885 18275
rect 37749 18241 37783 18275
rect 38117 18241 38151 18275
rect 38393 18241 38427 18275
rect 38853 18241 38887 18275
rect 39037 18241 39071 18275
rect 39773 18241 39807 18275
rect 40233 18241 40267 18275
rect 41797 18241 41831 18275
rect 41981 18241 42015 18275
rect 42625 18241 42659 18275
rect 56885 18241 56919 18275
rect 58081 18241 58115 18275
rect 58265 18241 58299 18275
rect 1777 18173 1811 18207
rect 14841 18173 14875 18207
rect 15025 18173 15059 18207
rect 15117 18173 15151 18207
rect 15301 18173 15335 18207
rect 15945 18173 15979 18207
rect 17877 18173 17911 18207
rect 30757 18173 30791 18207
rect 40325 18173 40359 18207
rect 10333 18105 10367 18139
rect 16037 18037 16071 18071
rect 18429 18037 18463 18071
rect 23765 18037 23799 18071
rect 27261 18037 27295 18071
rect 29193 18037 29227 18071
rect 33333 18037 33367 18071
rect 34989 18037 35023 18071
rect 38117 18037 38151 18071
rect 44005 18037 44039 18071
rect 21005 17833 21039 17867
rect 41797 17833 41831 17867
rect 15761 17765 15795 17799
rect 25789 17765 25823 17799
rect 30297 17765 30331 17799
rect 32873 17765 32907 17799
rect 37657 17765 37691 17799
rect 17969 17697 18003 17731
rect 22569 17697 22603 17731
rect 25329 17697 25363 17731
rect 38209 17697 38243 17731
rect 58173 17697 58207 17731
rect 1593 17629 1627 17663
rect 15669 17629 15703 17663
rect 16497 17629 16531 17663
rect 17417 17629 17451 17663
rect 18521 17629 18555 17663
rect 18705 17629 18739 17663
rect 19809 17629 19843 17663
rect 24593 17629 24627 17663
rect 25421 17629 25455 17663
rect 26249 17629 26283 17663
rect 29765 17629 29799 17663
rect 30118 17629 30152 17663
rect 30849 17629 30883 17663
rect 31125 17629 31159 17663
rect 31769 17629 31803 17663
rect 32045 17629 32079 17663
rect 32137 17629 32171 17663
rect 33057 17629 33091 17663
rect 33149 17629 33183 17663
rect 33333 17629 33367 17663
rect 33425 17629 33459 17663
rect 35725 17629 35759 17663
rect 38025 17629 38059 17663
rect 41978 17629 42012 17663
rect 42349 17629 42383 17663
rect 42441 17629 42475 17663
rect 57897 17629 57931 17663
rect 1869 17561 1903 17595
rect 16313 17561 16347 17595
rect 22836 17561 22870 17595
rect 29929 17561 29963 17595
rect 30021 17561 30055 17595
rect 31953 17561 31987 17595
rect 35992 17561 36026 17595
rect 57069 17561 57103 17595
rect 16589 17493 16623 17527
rect 18889 17493 18923 17527
rect 23949 17493 23983 17527
rect 24685 17493 24719 17527
rect 27445 17493 27479 17527
rect 30941 17493 30975 17527
rect 32321 17493 32355 17527
rect 37105 17493 37139 17527
rect 38117 17493 38151 17527
rect 41981 17493 42015 17527
rect 57161 17493 57195 17527
rect 19993 17289 20027 17323
rect 21465 17289 21499 17323
rect 34897 17289 34931 17323
rect 21005 17221 21039 17255
rect 28917 17221 28951 17255
rect 32505 17221 32539 17255
rect 33609 17221 33643 17255
rect 40141 17221 40175 17255
rect 1593 17153 1627 17187
rect 15669 17153 15703 17187
rect 17417 17153 17451 17187
rect 17785 17153 17819 17187
rect 17877 17153 17911 17187
rect 18705 17153 18739 17187
rect 18981 17153 19015 17187
rect 19993 17153 20027 17187
rect 20177 17153 20211 17187
rect 20361 17153 20395 17187
rect 22017 17153 22051 17187
rect 22201 17153 22235 17187
rect 22845 17153 22879 17187
rect 26249 17153 26283 17187
rect 26341 17153 26375 17187
rect 26433 17153 26467 17187
rect 26617 17153 26651 17187
rect 27169 17153 27203 17187
rect 30001 17153 30035 17187
rect 30094 17153 30128 17187
rect 30205 17153 30239 17187
rect 30389 17153 30423 17187
rect 30849 17153 30883 17187
rect 32321 17153 32355 17187
rect 33333 17153 33367 17187
rect 33481 17153 33515 17187
rect 33698 17153 33732 17187
rect 33798 17153 33832 17187
rect 34437 17153 34471 17187
rect 34713 17153 34747 17187
rect 39037 17153 39071 17187
rect 39221 17153 39255 17187
rect 39865 17153 39899 17187
rect 57069 17153 57103 17187
rect 1777 17085 1811 17119
rect 19257 17085 19291 17119
rect 31033 17085 31067 17119
rect 32689 17085 32723 17119
rect 34529 17085 34563 17119
rect 57345 17085 57379 17119
rect 17233 17017 17267 17051
rect 18797 17017 18831 17051
rect 21373 17017 21407 17051
rect 24041 17017 24075 17051
rect 33977 17017 34011 17051
rect 15761 16949 15795 16983
rect 22385 16949 22419 16983
rect 25973 16949 26007 16983
rect 29745 16949 29779 16983
rect 39405 16949 39439 16983
rect 16681 16745 16715 16779
rect 22937 16745 22971 16779
rect 24593 16745 24627 16779
rect 31677 16745 31711 16779
rect 40049 16745 40083 16779
rect 17877 16677 17911 16711
rect 19579 16677 19613 16711
rect 21005 16677 21039 16711
rect 33057 16677 33091 16711
rect 11345 16609 11379 16643
rect 11713 16609 11747 16643
rect 14749 16609 14783 16643
rect 14841 16609 14875 16643
rect 15025 16609 15059 16643
rect 19809 16609 19843 16643
rect 25053 16609 25087 16643
rect 29837 16609 29871 16643
rect 32137 16609 32171 16643
rect 36829 16609 36863 16643
rect 39221 16609 39255 16643
rect 40233 16609 40267 16643
rect 40601 16609 40635 16643
rect 56057 16609 56091 16643
rect 56425 16609 56459 16643
rect 56885 16609 56919 16643
rect 11253 16541 11287 16575
rect 11621 16541 11655 16575
rect 14933 16541 14967 16575
rect 16037 16541 16071 16575
rect 16221 16541 16255 16575
rect 16681 16541 16715 16575
rect 16865 16541 16899 16575
rect 17325 16541 17359 16575
rect 17601 16541 17635 16575
rect 17693 16541 17727 16575
rect 18521 16541 18555 16575
rect 18613 16541 18647 16575
rect 18797 16541 18831 16575
rect 18889 16541 18923 16575
rect 19671 16541 19705 16575
rect 20637 16541 20671 16575
rect 21741 16541 21775 16575
rect 24777 16541 24811 16575
rect 24869 16541 24903 16575
rect 25145 16541 25179 16575
rect 26065 16541 26099 16575
rect 26157 16541 26191 16575
rect 26249 16541 26283 16575
rect 26433 16541 26467 16575
rect 26893 16541 26927 16575
rect 30093 16541 30127 16575
rect 31861 16541 31895 16575
rect 31953 16541 31987 16575
rect 32229 16541 32263 16575
rect 36645 16541 36679 16575
rect 39037 16541 39071 16575
rect 40325 16541 40359 16575
rect 56241 16541 56275 16575
rect 57141 16541 57175 16575
rect 10609 16473 10643 16507
rect 17509 16473 17543 16507
rect 19441 16473 19475 16507
rect 20177 16473 20211 16507
rect 32689 16473 32723 16507
rect 32873 16473 32907 16507
rect 40693 16473 40727 16507
rect 14565 16405 14599 16439
rect 16129 16405 16163 16439
rect 18337 16405 18371 16439
rect 21097 16405 21131 16439
rect 25421 16405 25455 16439
rect 25789 16405 25823 16439
rect 28089 16405 28123 16439
rect 31217 16405 31251 16439
rect 36277 16405 36311 16439
rect 36737 16405 36771 16439
rect 58265 16405 58299 16439
rect 16957 16201 16991 16235
rect 17877 16201 17911 16235
rect 23857 16201 23891 16235
rect 31309 16201 31343 16235
rect 34161 16201 34195 16235
rect 57253 16201 57287 16235
rect 15945 16133 15979 16167
rect 21373 16133 21407 16167
rect 22744 16133 22778 16167
rect 30174 16133 30208 16167
rect 56977 16133 57011 16167
rect 1593 16065 1627 16099
rect 16129 16065 16163 16099
rect 17141 16065 17175 16099
rect 17325 16065 17359 16099
rect 17417 16065 17451 16099
rect 18061 16065 18095 16099
rect 18245 16065 18279 16099
rect 18797 16065 18831 16099
rect 19073 16065 19107 16099
rect 20361 16065 20395 16099
rect 21189 16065 21223 16099
rect 21465 16065 21499 16099
rect 24317 16065 24351 16099
rect 27169 16065 27203 16099
rect 29929 16065 29963 16099
rect 32505 16065 32539 16099
rect 35449 16065 35483 16099
rect 35716 16065 35750 16099
rect 39497 16065 39531 16099
rect 39764 16065 39798 16099
rect 56701 16065 56735 16099
rect 56885 16065 56919 16099
rect 57069 16065 57103 16099
rect 1777 15997 1811 16031
rect 18337 15997 18371 16031
rect 19349 15997 19383 16031
rect 20453 15997 20487 16031
rect 22477 15997 22511 16031
rect 32689 15997 32723 16031
rect 34253 15997 34287 16031
rect 34345 15997 34379 16031
rect 18889 15929 18923 15963
rect 28365 15929 28399 15963
rect 40877 15929 40911 15963
rect 16313 15861 16347 15895
rect 20729 15861 20763 15895
rect 21189 15861 21223 15895
rect 25513 15861 25547 15895
rect 33793 15861 33827 15895
rect 36829 15861 36863 15895
rect 18705 15657 18739 15691
rect 19809 15657 19843 15691
rect 48145 15657 48179 15691
rect 17877 15589 17911 15623
rect 23029 15589 23063 15623
rect 19441 15521 19475 15555
rect 24593 15521 24627 15555
rect 30849 15521 30883 15555
rect 34253 15521 34287 15555
rect 35449 15521 35483 15555
rect 58265 15521 58299 15555
rect 1593 15453 1627 15487
rect 15117 15453 15151 15487
rect 17877 15453 17911 15487
rect 18061 15453 18095 15487
rect 19625 15453 19659 15487
rect 20269 15453 20303 15487
rect 23581 15453 23615 15487
rect 26893 15453 26927 15487
rect 29745 15453 29779 15487
rect 32505 15453 32539 15487
rect 56977 15453 57011 15487
rect 57989 15453 58023 15487
rect 1869 15385 1903 15419
rect 18521 15385 18555 15419
rect 18737 15385 18771 15419
rect 23397 15385 23431 15419
rect 24860 15385 24894 15419
rect 35265 15385 35299 15419
rect 46857 15385 46891 15419
rect 57253 15385 57287 15419
rect 16313 15317 16347 15351
rect 18889 15317 18923 15351
rect 21465 15317 21499 15351
rect 23213 15317 23247 15351
rect 23305 15317 23339 15351
rect 25973 15317 26007 15351
rect 29101 15317 29135 15351
rect 34897 15317 34931 15351
rect 35357 15317 35391 15351
rect 14197 15113 14231 15147
rect 18061 15045 18095 15079
rect 20260 15045 20294 15079
rect 22744 15045 22778 15079
rect 1593 14977 1627 15011
rect 19165 14977 19199 15011
rect 24317 14977 24351 15011
rect 27169 14977 27203 15011
rect 30297 14977 30331 15011
rect 30564 14977 30598 15011
rect 32873 14977 32907 15011
rect 33140 14977 33174 15011
rect 34713 14977 34747 15011
rect 34980 14977 35014 15011
rect 1777 14909 1811 14943
rect 13737 14909 13771 14943
rect 14657 14909 14691 14943
rect 14933 14909 14967 14943
rect 17141 14909 17175 14943
rect 19073 14909 19107 14943
rect 19993 14909 20027 14943
rect 22477 14909 22511 14943
rect 28273 14909 28307 14943
rect 14013 14841 14047 14875
rect 17509 14841 17543 14875
rect 18429 14841 18463 14875
rect 18521 14841 18555 14875
rect 23857 14841 23891 14875
rect 16221 14773 16255 14807
rect 17601 14773 17635 14807
rect 19441 14773 19475 14807
rect 21373 14773 21407 14807
rect 25513 14773 25547 14807
rect 31677 14773 31711 14807
rect 34253 14773 34287 14807
rect 36093 14773 36127 14807
rect 15485 14569 15519 14603
rect 22937 14569 22971 14603
rect 31217 14569 31251 14603
rect 58081 14569 58115 14603
rect 30297 14501 30331 14535
rect 15301 14433 15335 14467
rect 17141 14433 17175 14467
rect 24685 14433 24719 14467
rect 32689 14433 32723 14467
rect 1593 14365 1627 14399
rect 15209 14365 15243 14399
rect 16037 14365 16071 14399
rect 19625 14365 19659 14399
rect 19901 14365 19935 14399
rect 21741 14365 21775 14399
rect 24777 14365 24811 14399
rect 26157 14365 26191 14399
rect 28457 14365 28491 14399
rect 29101 14365 29135 14399
rect 29929 14365 29963 14399
rect 30113 14365 30147 14399
rect 30389 14365 30423 14399
rect 30757 14365 30791 14399
rect 31493 14365 31527 14399
rect 31585 14365 31619 14399
rect 31677 14365 31711 14399
rect 31861 14365 31895 14399
rect 32505 14365 32539 14399
rect 57989 14365 58023 14399
rect 1869 14297 1903 14331
rect 32321 14297 32355 14331
rect 21189 14229 21223 14263
rect 25145 14229 25179 14263
rect 29101 14229 29135 14263
rect 15209 14025 15243 14059
rect 20361 14025 20395 14059
rect 23397 14025 23431 14059
rect 28549 14025 28583 14059
rect 32413 14025 32447 14059
rect 40049 14025 40083 14059
rect 29377 13957 29411 13991
rect 33793 13957 33827 13991
rect 14013 13889 14047 13923
rect 19165 13889 19199 13923
rect 22017 13889 22051 13923
rect 22284 13889 22318 13923
rect 24041 13889 24075 13923
rect 27169 13889 27203 13923
rect 27436 13889 27470 13923
rect 30481 13889 30515 13923
rect 30941 13889 30975 13923
rect 31309 13889 31343 13923
rect 31401 13889 31435 13923
rect 32321 13889 32355 13923
rect 32505 13889 32539 13923
rect 33977 13889 34011 13923
rect 38761 13889 38795 13923
rect 57069 13889 57103 13923
rect 16865 13821 16899 13855
rect 17141 13821 17175 13855
rect 18521 13821 18555 13855
rect 25145 13821 25179 13855
rect 29469 13821 29503 13855
rect 29653 13821 29687 13855
rect 30757 13821 30791 13855
rect 57345 13821 57379 13855
rect 30573 13753 30607 13787
rect 29009 13685 29043 13719
rect 34161 13685 34195 13719
rect 20177 13481 20211 13515
rect 22293 13481 22327 13515
rect 23857 13481 23891 13515
rect 34253 13481 34287 13515
rect 58265 13481 58299 13515
rect 14473 13345 14507 13379
rect 14749 13345 14783 13379
rect 17693 13345 17727 13379
rect 19809 13345 19843 13379
rect 25697 13345 25731 13379
rect 27353 13345 27387 13379
rect 32873 13345 32907 13379
rect 56885 13345 56919 13379
rect 1593 13277 1627 13311
rect 1869 13277 1903 13311
rect 16589 13277 16623 13311
rect 19901 13277 19935 13311
rect 21097 13277 21131 13311
rect 23857 13277 23891 13311
rect 24041 13277 24075 13311
rect 24593 13277 24627 13311
rect 27620 13277 27654 13311
rect 29745 13277 29779 13311
rect 31861 13277 31895 13311
rect 31953 13277 31987 13311
rect 32137 13277 32171 13311
rect 32229 13277 32263 13311
rect 19533 13209 19567 13243
rect 19993 13209 20027 13243
rect 30012 13209 30046 13243
rect 33140 13209 33174 13243
rect 57130 13209 57164 13243
rect 16037 13141 16071 13175
rect 28733 13141 28767 13175
rect 31125 13141 31159 13175
rect 31677 13141 31711 13175
rect 18705 12937 18739 12971
rect 22201 12937 22235 12971
rect 27261 12937 27295 12971
rect 30849 12937 30883 12971
rect 31217 12937 31251 12971
rect 33701 12937 33735 12971
rect 58265 12937 58299 12971
rect 20913 12869 20947 12903
rect 22385 12869 22419 12903
rect 26341 12869 26375 12903
rect 49433 12869 49467 12903
rect 56977 12869 57011 12903
rect 1593 12801 1627 12835
rect 14657 12801 14691 12835
rect 17509 12801 17543 12835
rect 20729 12801 20763 12835
rect 22293 12801 22327 12835
rect 23397 12801 23431 12835
rect 26157 12801 26191 12835
rect 26433 12801 26467 12835
rect 27169 12801 27203 12835
rect 27353 12801 27387 12835
rect 28089 12801 28123 12835
rect 33977 12801 34011 12835
rect 34069 12801 34103 12835
rect 34161 12801 34195 12835
rect 34345 12801 34379 12835
rect 56793 12801 56827 12835
rect 57069 12801 57103 12835
rect 58081 12801 58115 12835
rect 58265 12801 58299 12835
rect 1777 12733 1811 12767
rect 14933 12733 14967 12767
rect 21005 12733 21039 12767
rect 22569 12733 22603 12767
rect 24869 12733 24903 12767
rect 31309 12733 31343 12767
rect 31401 12733 31435 12767
rect 22017 12665 22051 12699
rect 26157 12665 26191 12699
rect 56793 12665 56827 12699
rect 16037 12597 16071 12631
rect 20453 12597 20487 12631
rect 29285 12597 29319 12631
rect 50905 12597 50939 12631
rect 13093 12393 13127 12427
rect 17785 12393 17819 12427
rect 19993 12393 20027 12427
rect 27261 12393 27295 12427
rect 31033 12393 31067 12427
rect 13369 12257 13403 12291
rect 13461 12257 13495 12291
rect 15853 12257 15887 12291
rect 20361 12257 20395 12291
rect 25237 12257 25271 12291
rect 30297 12257 30331 12291
rect 1593 12189 1627 12223
rect 13277 12189 13311 12223
rect 13553 12189 13587 12223
rect 15761 12189 15795 12223
rect 16589 12189 16623 12223
rect 20545 12189 20579 12223
rect 21741 12189 21775 12223
rect 26065 12189 26099 12223
rect 30113 12189 30147 12223
rect 30941 12189 30975 12223
rect 56977 12189 57011 12223
rect 57989 12189 58023 12223
rect 1869 12121 1903 12155
rect 20453 12121 20487 12155
rect 24961 12121 24995 12155
rect 57253 12121 57287 12155
rect 16129 12053 16163 12087
rect 23121 12053 23155 12087
rect 24593 12053 24627 12087
rect 25053 12053 25087 12087
rect 29745 12053 29779 12087
rect 30205 12053 30239 12087
rect 58081 12053 58115 12087
rect 13001 11849 13035 11883
rect 15945 11849 15979 11883
rect 17049 11849 17083 11883
rect 17601 11849 17635 11883
rect 22661 11849 22695 11883
rect 23765 11849 23799 11883
rect 25513 11849 25547 11883
rect 30481 11849 30515 11883
rect 35173 11849 35207 11883
rect 27712 11781 27746 11815
rect 34077 11781 34111 11815
rect 1593 11713 1627 11747
rect 13185 11713 13219 11747
rect 13369 11713 13403 11747
rect 15577 11713 15611 11747
rect 15761 11713 15795 11747
rect 16957 11713 16991 11747
rect 17141 11713 17175 11747
rect 17877 11713 17911 11747
rect 19625 11713 19659 11747
rect 22845 11713 22879 11747
rect 23121 11713 23155 11747
rect 23673 11713 23707 11747
rect 23857 11713 23891 11747
rect 24317 11713 24351 11747
rect 27445 11713 27479 11747
rect 29285 11713 29319 11747
rect 33701 11713 33735 11747
rect 33849 11713 33883 11747
rect 33977 11713 34011 11747
rect 34166 11713 34200 11747
rect 38209 11713 38243 11747
rect 57161 11713 57195 11747
rect 1777 11645 1811 11679
rect 13277 11645 13311 11679
rect 13461 11645 13495 11679
rect 17785 11645 17819 11679
rect 17969 11645 18003 11679
rect 18061 11645 18095 11679
rect 18613 11645 18647 11679
rect 19809 11645 19843 11679
rect 22937 11645 22971 11679
rect 23029 11645 23063 11679
rect 35265 11645 35299 11679
rect 35357 11645 35391 11679
rect 38393 11645 38427 11679
rect 18889 11577 18923 11611
rect 19073 11509 19107 11543
rect 28825 11509 28859 11543
rect 34345 11509 34379 11543
rect 34805 11509 34839 11543
rect 57253 11509 57287 11543
rect 13461 11305 13495 11339
rect 20821 11305 20855 11339
rect 21281 11305 21315 11339
rect 23029 11305 23063 11339
rect 24593 11305 24627 11339
rect 36277 11305 36311 11339
rect 58265 11305 58299 11339
rect 13277 11237 13311 11271
rect 18245 11169 18279 11203
rect 21741 11169 21775 11203
rect 21925 11169 21959 11203
rect 22661 11169 22695 11203
rect 28917 11169 28951 11203
rect 34253 11169 34287 11203
rect 38669 11169 38703 11203
rect 56885 11169 56919 11203
rect 17969 11101 18003 11135
rect 19441 11101 19475 11135
rect 21649 11101 21683 11135
rect 22845 11101 22879 11135
rect 24593 11101 24627 11135
rect 24777 11101 24811 11135
rect 25605 11101 25639 11135
rect 32965 11101 32999 11135
rect 34897 11101 34931 11135
rect 35153 11101 35187 11135
rect 36737 11101 36771 11135
rect 38393 11101 38427 11135
rect 13001 11033 13035 11067
rect 19686 11033 19720 11067
rect 28825 11033 28859 11067
rect 32413 11033 32447 11067
rect 32597 11033 32631 11067
rect 32699 11033 32733 11067
rect 34069 11033 34103 11067
rect 37473 11033 37507 11067
rect 57130 11033 57164 11067
rect 17601 10965 17635 10999
rect 18061 10965 18095 10999
rect 26801 10965 26835 10999
rect 28365 10965 28399 10999
rect 28733 10965 28767 10999
rect 32781 10965 32815 10999
rect 33609 10965 33643 10999
rect 33977 10965 34011 10999
rect 14749 10761 14783 10795
rect 21465 10761 21499 10795
rect 22385 10761 22419 10795
rect 36001 10693 36035 10727
rect 56793 10693 56827 10727
rect 56977 10693 57011 10727
rect 58173 10693 58207 10727
rect 1593 10625 1627 10659
rect 2421 10625 2455 10659
rect 13093 10625 13127 10659
rect 13277 10625 13311 10659
rect 17693 10625 17727 10659
rect 20085 10625 20119 10659
rect 20352 10625 20386 10659
rect 23673 10625 23707 10659
rect 23940 10625 23974 10659
rect 26433 10625 26467 10659
rect 27169 10625 27203 10659
rect 29285 10625 29319 10659
rect 29469 10625 29503 10659
rect 33885 10625 33919 10659
rect 34141 10625 34175 10659
rect 35725 10625 35759 10659
rect 35909 10625 35943 10659
rect 36093 10625 36127 10659
rect 37740 10625 37774 10659
rect 57069 10625 57103 10659
rect 58081 10625 58115 10659
rect 58265 10625 58299 10659
rect 1777 10557 1811 10591
rect 13185 10557 13219 10591
rect 13369 10557 13403 10591
rect 14933 10557 14967 10591
rect 15025 10557 15059 10591
rect 15117 10557 15151 10591
rect 15209 10557 15243 10591
rect 17785 10557 17819 10591
rect 17877 10557 17911 10591
rect 22477 10557 22511 10591
rect 22661 10557 22695 10591
rect 26249 10557 26283 10591
rect 27445 10557 27479 10591
rect 37473 10557 37507 10591
rect 17325 10489 17359 10523
rect 28549 10489 28583 10523
rect 56793 10489 56827 10523
rect 12909 10421 12943 10455
rect 22017 10421 22051 10455
rect 25053 10421 25087 10455
rect 26617 10421 26651 10455
rect 29377 10421 29411 10455
rect 35265 10421 35299 10455
rect 36277 10421 36311 10455
rect 38853 10421 38887 10455
rect 13277 10217 13311 10251
rect 23949 10217 23983 10251
rect 25789 10217 25823 10251
rect 37841 10217 37875 10251
rect 13093 10149 13127 10183
rect 14565 10149 14599 10183
rect 21925 10149 21959 10183
rect 57253 10149 57287 10183
rect 30941 10081 30975 10115
rect 38301 10081 38335 10115
rect 38393 10081 38427 10115
rect 58173 10081 58207 10115
rect 1593 10013 1627 10047
rect 20545 10013 20579 10047
rect 20812 10013 20846 10047
rect 23673 10013 23707 10047
rect 23765 10013 23799 10047
rect 24593 10013 24627 10047
rect 27721 10013 27755 10047
rect 29745 10013 29779 10047
rect 29929 10013 29963 10047
rect 30021 10013 30055 10047
rect 30113 10013 30147 10047
rect 30297 10013 30331 10047
rect 31217 10013 31251 10047
rect 38209 10013 38243 10047
rect 40233 10013 40267 10047
rect 57897 10013 57931 10047
rect 1869 9945 1903 9979
rect 12817 9945 12851 9979
rect 14289 9945 14323 9979
rect 27966 9945 28000 9979
rect 40509 9945 40543 9979
rect 57069 9945 57103 9979
rect 14749 9877 14783 9911
rect 29101 9877 29135 9911
rect 30481 9877 30515 9911
rect 32321 9877 32355 9911
rect 27169 9673 27203 9707
rect 30757 9673 30791 9707
rect 12449 9605 12483 9639
rect 14013 9605 14047 9639
rect 29929 9605 29963 9639
rect 1593 9537 1627 9571
rect 19809 9537 19843 9571
rect 27425 9537 27459 9571
rect 27537 9537 27571 9571
rect 27650 9537 27684 9571
rect 27813 9537 27847 9571
rect 28273 9537 28307 9571
rect 28365 9537 28399 9571
rect 30113 9537 30147 9571
rect 30987 9537 31021 9571
rect 31125 9537 31159 9571
rect 31217 9543 31251 9577
rect 31401 9537 31435 9571
rect 34989 9537 35023 9571
rect 35081 9537 35115 9571
rect 35265 9537 35299 9571
rect 37933 9537 37967 9571
rect 38117 9537 38151 9571
rect 39589 9537 39623 9571
rect 40509 9537 40543 9571
rect 40776 9537 40810 9571
rect 57345 9537 57379 9571
rect 57529 9537 57563 9571
rect 1777 9469 1811 9503
rect 12909 9469 12943 9503
rect 14473 9469 14507 9503
rect 19901 9469 19935 9503
rect 20085 9469 20119 9503
rect 30297 9469 30331 9503
rect 35449 9469 35483 9503
rect 39865 9469 39899 9503
rect 12725 9401 12759 9435
rect 14289 9401 14323 9435
rect 19441 9333 19475 9367
rect 28181 9333 28215 9367
rect 38025 9333 38059 9367
rect 41889 9333 41923 9367
rect 57437 9333 57471 9367
rect 20821 9129 20855 9163
rect 37381 9129 37415 9163
rect 39037 9129 39071 9163
rect 41429 9129 41463 9163
rect 34989 9061 35023 9095
rect 23765 8993 23799 9027
rect 24593 8993 24627 9027
rect 30665 8993 30699 9027
rect 41061 8993 41095 9027
rect 56885 8993 56919 9027
rect 1593 8925 1627 8959
rect 19441 8925 19475 8959
rect 19697 8925 19731 8959
rect 23581 8925 23615 8959
rect 30849 8925 30883 8959
rect 30941 8925 30975 8959
rect 31125 8925 31159 8959
rect 31217 8925 31251 8959
rect 31861 8925 31895 8959
rect 32045 8925 32079 8959
rect 32137 8925 32171 8959
rect 32597 8925 32631 8959
rect 32781 8925 32815 8959
rect 35173 8925 35207 8959
rect 35265 8925 35299 8959
rect 35449 8925 35483 8959
rect 35541 8925 35575 8959
rect 37289 8925 37323 8959
rect 37749 8925 37783 8959
rect 40049 8925 40083 8959
rect 40325 8925 40359 8959
rect 40417 8925 40451 8959
rect 41245 8925 41279 8959
rect 1869 8857 1903 8891
rect 24860 8857 24894 8891
rect 38025 8857 38059 8891
rect 38485 8857 38519 8891
rect 38853 8857 38887 8891
rect 40233 8857 40267 8891
rect 57152 8857 57186 8891
rect 25973 8789 26007 8823
rect 31677 8789 31711 8823
rect 32689 8789 32723 8823
rect 39053 8789 39087 8823
rect 39221 8789 39255 8823
rect 40601 8789 40635 8823
rect 58265 8789 58299 8823
rect 11805 8585 11839 8619
rect 24317 8585 24351 8619
rect 25881 8585 25915 8619
rect 26249 8585 26283 8619
rect 29745 8585 29779 8619
rect 34989 8585 35023 8619
rect 56333 8585 56367 8619
rect 58265 8585 58299 8619
rect 18245 8517 18279 8551
rect 26341 8517 26375 8551
rect 27997 8517 28031 8551
rect 29009 8517 29043 8551
rect 30665 8517 30699 8551
rect 34621 8517 34655 8551
rect 34713 8517 34747 8551
rect 57345 8517 57379 8551
rect 58081 8517 58115 8551
rect 12081 8449 12115 8483
rect 13001 8449 13035 8483
rect 19073 8449 19107 8483
rect 19329 8449 19363 8483
rect 23121 8449 23155 8483
rect 28181 8449 28215 8483
rect 28825 8449 28859 8483
rect 29653 8449 29687 8483
rect 30481 8449 30515 8483
rect 30757 8449 30791 8483
rect 31493 8449 31527 8483
rect 31585 8449 31619 8483
rect 32597 8449 32631 8483
rect 32781 8449 32815 8483
rect 33425 8449 33459 8483
rect 34345 8449 34379 8483
rect 34438 8449 34472 8483
rect 34851 8449 34885 8483
rect 35449 8449 35483 8483
rect 37565 8449 37599 8483
rect 38301 8449 38335 8483
rect 38669 8449 38703 8483
rect 39773 8449 39807 8483
rect 56241 8449 56275 8483
rect 57069 8449 57103 8483
rect 58357 8449 58391 8483
rect 11989 8381 12023 8415
rect 12173 8381 12207 8415
rect 12265 8381 12299 8415
rect 12817 8381 12851 8415
rect 13093 8381 13127 8415
rect 13185 8381 13219 8415
rect 13277 8381 13311 8415
rect 18337 8381 18371 8415
rect 18521 8381 18555 8415
rect 26433 8381 26467 8415
rect 31401 8381 31435 8415
rect 31677 8381 31711 8415
rect 32689 8381 32723 8415
rect 33701 8381 33735 8415
rect 35633 8381 35667 8415
rect 40049 8381 40083 8415
rect 17877 8313 17911 8347
rect 29193 8313 29227 8347
rect 30297 8313 30331 8347
rect 31217 8313 31251 8347
rect 58081 8313 58115 8347
rect 20453 8245 20487 8279
rect 28365 8245 28399 8279
rect 37657 8245 37691 8279
rect 12081 8041 12115 8075
rect 17141 8041 17175 8075
rect 38393 8041 38427 8075
rect 38853 8041 38887 8075
rect 40141 8041 40175 8075
rect 11897 7973 11931 8007
rect 17325 7973 17359 8007
rect 28457 7973 28491 8007
rect 30757 7973 30791 8007
rect 38485 7973 38519 8007
rect 56149 7973 56183 8007
rect 19533 7905 19567 7939
rect 31033 7905 31067 7939
rect 31217 7905 31251 7939
rect 32137 7905 32171 7939
rect 32229 7905 32263 7939
rect 32965 7905 32999 7939
rect 33425 7905 33459 7939
rect 33517 7905 33551 7939
rect 34897 7905 34931 7939
rect 36277 7905 36311 7939
rect 38025 7905 38059 7939
rect 38577 7905 38611 7939
rect 56885 7905 56919 7939
rect 1593 7837 1627 7871
rect 16773 7837 16807 7871
rect 18337 7837 18371 7871
rect 23489 7837 23523 7871
rect 24041 7837 24075 7871
rect 25145 7837 25179 7871
rect 27077 7837 27111 7871
rect 30021 7837 30055 7871
rect 30297 7837 30331 7871
rect 30941 7837 30975 7871
rect 31125 7837 31159 7871
rect 31769 7837 31803 7871
rect 32321 7837 32355 7871
rect 35173 7837 35207 7871
rect 37197 7837 37231 7871
rect 37289 7837 37323 7871
rect 37473 7837 37507 7871
rect 37565 7837 37599 7871
rect 40049 7837 40083 7871
rect 40325 7837 40359 7871
rect 55505 7837 55539 7871
rect 55689 7837 55723 7871
rect 56425 7837 56459 7871
rect 57141 7837 57175 7871
rect 1869 7769 1903 7803
rect 11621 7769 11655 7803
rect 18613 7769 18647 7803
rect 19800 7769 19834 7803
rect 23673 7769 23707 7803
rect 25412 7769 25446 7803
rect 27445 7769 27479 7803
rect 28273 7769 28307 7803
rect 29837 7769 29871 7803
rect 56149 7769 56183 7803
rect 17150 7701 17184 7735
rect 20913 7701 20947 7735
rect 23765 7701 23799 7735
rect 23857 7701 23891 7735
rect 26525 7701 26559 7735
rect 30205 7701 30239 7735
rect 33149 7701 33183 7735
rect 37013 7701 37047 7735
rect 55689 7701 55723 7735
rect 56333 7701 56367 7735
rect 58265 7701 58299 7735
rect 11805 7497 11839 7531
rect 13277 7497 13311 7531
rect 17877 7497 17911 7531
rect 24685 7497 24719 7531
rect 28365 7497 28399 7531
rect 31217 7497 31251 7531
rect 32413 7497 32447 7531
rect 33793 7497 33827 7531
rect 34989 7497 35023 7531
rect 18245 7429 18279 7463
rect 18337 7429 18371 7463
rect 23397 7429 23431 7463
rect 29929 7429 29963 7463
rect 39773 7429 39807 7463
rect 57345 7429 57379 7463
rect 58265 7429 58299 7463
rect 1593 7361 1627 7395
rect 11989 7361 12023 7395
rect 12173 7361 12207 7395
rect 12817 7361 12851 7395
rect 20361 7361 20395 7395
rect 20453 7361 20487 7395
rect 27169 7361 27203 7395
rect 32321 7361 32355 7395
rect 32505 7361 32539 7395
rect 33149 7361 33183 7395
rect 33333 7361 33367 7395
rect 33609 7361 33643 7395
rect 34161 7361 34195 7395
rect 35265 7361 35299 7395
rect 35357 7361 35391 7395
rect 35449 7361 35483 7395
rect 35633 7361 35667 7395
rect 37565 7361 37599 7395
rect 37657 7361 37691 7395
rect 38761 7361 38795 7395
rect 39037 7361 39071 7395
rect 39681 7361 39715 7395
rect 56149 7361 56183 7395
rect 57069 7361 57103 7395
rect 58081 7361 58115 7395
rect 58357 7361 58391 7395
rect 1777 7293 1811 7327
rect 12081 7293 12115 7327
rect 12265 7293 12299 7327
rect 18521 7293 18555 7327
rect 20637 7293 20671 7327
rect 34069 7293 34103 7327
rect 37381 7293 37415 7327
rect 38853 7293 38887 7327
rect 56425 7293 56459 7327
rect 13093 7225 13127 7259
rect 19993 7225 20027 7259
rect 33149 7225 33183 7259
rect 39221 7225 39255 7259
rect 34621 7157 34655 7191
rect 37841 7157 37875 7191
rect 38393 7157 38427 7191
rect 38761 7157 38795 7191
rect 58081 7157 58115 7191
rect 13645 6885 13679 6919
rect 15209 6885 15243 6919
rect 22385 6885 22419 6919
rect 23489 6885 23523 6919
rect 11069 6817 11103 6851
rect 11253 6817 11287 6851
rect 11345 6817 11379 6851
rect 15393 6817 15427 6851
rect 20177 6817 20211 6851
rect 24593 6817 24627 6851
rect 31493 6817 31527 6851
rect 32689 6817 32723 6851
rect 34345 6817 34379 6851
rect 36001 6817 36035 6851
rect 37197 6817 37231 6851
rect 37841 6817 37875 6851
rect 39037 6817 39071 6851
rect 1593 6749 1627 6783
rect 9413 6749 9447 6783
rect 9505 6749 9539 6783
rect 9689 6749 9723 6783
rect 11437 6749 11471 6783
rect 11529 6749 11563 6783
rect 13277 6749 13311 6783
rect 22707 6749 22741 6783
rect 22937 6749 22971 6783
rect 23673 6749 23707 6783
rect 23764 6749 23798 6783
rect 23949 6749 23983 6783
rect 24036 6749 24070 6783
rect 25145 6749 25179 6783
rect 26433 6749 26467 6783
rect 28641 6749 28675 6783
rect 28733 6749 28767 6783
rect 28825 6749 28859 6783
rect 29009 6749 29043 6783
rect 31217 6749 31251 6783
rect 31310 6749 31344 6783
rect 31402 6749 31436 6783
rect 32873 6749 32907 6783
rect 35633 6749 35667 6783
rect 38117 6749 38151 6783
rect 38209 6749 38243 6783
rect 38301 6749 38335 6783
rect 38485 6749 38519 6783
rect 38945 6749 38979 6783
rect 39129 6749 39163 6783
rect 56885 6749 56919 6783
rect 57152 6749 57186 6783
rect 1869 6681 1903 6715
rect 10149 6681 10183 6715
rect 14933 6681 14967 6715
rect 19441 6681 19475 6715
rect 22569 6681 22603 6715
rect 24777 6681 24811 6715
rect 26700 6681 26734 6715
rect 33977 6681 34011 6715
rect 34161 6681 34195 6715
rect 35449 6681 35483 6715
rect 13737 6613 13771 6647
rect 22753 6613 22787 6647
rect 24869 6613 24903 6647
rect 24961 6613 24995 6647
rect 27813 6613 27847 6647
rect 28365 6613 28399 6647
rect 31033 6613 31067 6647
rect 33057 6613 33091 6647
rect 36553 6613 36587 6647
rect 36921 6613 36955 6647
rect 37013 6613 37047 6647
rect 58265 6613 58299 6647
rect 11161 6409 11195 6443
rect 12173 6409 12207 6443
rect 16313 6409 16347 6443
rect 17877 6409 17911 6443
rect 20453 6409 20487 6443
rect 23857 6409 23891 6443
rect 24961 6409 24995 6443
rect 25789 6409 25823 6443
rect 26249 6409 26283 6443
rect 27169 6409 27203 6443
rect 27537 6409 27571 6443
rect 30021 6409 30055 6443
rect 57529 6409 57563 6443
rect 13645 6341 13679 6375
rect 18245 6341 18279 6375
rect 19318 6341 19352 6375
rect 24041 6341 24075 6375
rect 33048 6341 33082 6375
rect 36645 6341 36679 6375
rect 37749 6341 37783 6375
rect 1593 6273 1627 6307
rect 19073 6273 19107 6307
rect 22569 6273 22603 6307
rect 23673 6273 23707 6307
rect 23811 6273 23845 6307
rect 24869 6273 24903 6307
rect 26157 6273 26191 6307
rect 28641 6273 28675 6307
rect 30849 6273 30883 6307
rect 31125 6273 31159 6307
rect 32781 6273 32815 6307
rect 36277 6273 36311 6307
rect 37473 6273 37507 6307
rect 57345 6273 57379 6307
rect 57529 6273 57563 6307
rect 1777 6205 1811 6239
rect 10701 6205 10735 6239
rect 11713 6205 11747 6239
rect 15853 6205 15887 6239
rect 18337 6205 18371 6239
rect 18521 6205 18555 6239
rect 22753 6205 22787 6239
rect 25145 6205 25179 6239
rect 26433 6205 26467 6239
rect 27629 6205 27663 6239
rect 27721 6205 27755 6239
rect 28917 6205 28951 6239
rect 10977 6137 11011 6171
rect 11989 6137 12023 6171
rect 14013 6137 14047 6171
rect 16129 6137 16163 6171
rect 23489 6137 23523 6171
rect 31125 6137 31159 6171
rect 14105 6069 14139 6103
rect 24501 6069 24535 6103
rect 34161 6069 34195 6103
rect 11989 5865 12023 5899
rect 13645 5865 13679 5899
rect 32873 5865 32907 5899
rect 37841 5865 37875 5899
rect 12909 5797 12943 5831
rect 18153 5797 18187 5831
rect 23489 5797 23523 5831
rect 18705 5729 18739 5763
rect 19441 5729 19475 5763
rect 22477 5729 22511 5763
rect 25605 5729 25639 5763
rect 33517 5729 33551 5763
rect 36461 5729 36495 5763
rect 17693 5661 17727 5695
rect 21465 5661 21499 5695
rect 22661 5661 22695 5695
rect 23811 5661 23845 5695
rect 24041 5661 24075 5695
rect 24915 5661 24949 5695
rect 25789 5661 25823 5695
rect 26157 5661 26191 5695
rect 28161 5661 28195 5695
rect 28270 5658 28304 5692
rect 28370 5661 28404 5695
rect 28549 5661 28583 5695
rect 30297 5661 30331 5695
rect 30481 5661 30515 5695
rect 33241 5661 33275 5695
rect 33333 5661 33367 5695
rect 56977 5661 57011 5695
rect 57989 5661 58023 5695
rect 11897 5593 11931 5627
rect 12725 5593 12759 5627
rect 13553 5593 13587 5627
rect 14381 5593 14415 5627
rect 19686 5593 19720 5627
rect 21741 5593 21775 5627
rect 23029 5593 23063 5627
rect 23673 5593 23707 5627
rect 24593 5593 24627 5627
rect 24777 5593 24811 5627
rect 25145 5593 25179 5627
rect 34989 5593 35023 5627
rect 35725 5593 35759 5627
rect 35909 5593 35943 5627
rect 36728 5593 36762 5627
rect 57253 5593 57287 5627
rect 14473 5525 14507 5559
rect 18521 5525 18555 5559
rect 18613 5525 18647 5559
rect 20821 5525 20855 5559
rect 22753 5525 22787 5559
rect 22845 5525 22879 5559
rect 23857 5525 23891 5559
rect 24961 5525 24995 5559
rect 25881 5525 25915 5559
rect 25973 5525 26007 5559
rect 27905 5525 27939 5559
rect 29009 5525 29043 5559
rect 30665 5525 30699 5559
rect 35081 5525 35115 5559
rect 58081 5525 58115 5559
rect 12357 5321 12391 5355
rect 18429 5321 18463 5355
rect 18889 5321 18923 5355
rect 29469 5321 29503 5355
rect 30389 5321 30423 5355
rect 32689 5321 32723 5355
rect 33701 5321 33735 5355
rect 35449 5321 35483 5355
rect 36737 5321 36771 5355
rect 38393 5321 38427 5355
rect 39865 5321 39899 5355
rect 40601 5321 40635 5355
rect 42809 5321 42843 5355
rect 11161 5253 11195 5287
rect 13829 5253 13863 5287
rect 18153 5253 18187 5287
rect 19901 5253 19935 5287
rect 23664 5253 23698 5287
rect 25973 5253 26007 5287
rect 38301 5253 38335 5287
rect 56885 5253 56919 5287
rect 1593 5185 1627 5219
rect 10241 5185 10275 5219
rect 10977 5185 11011 5219
rect 12173 5185 12207 5219
rect 13645 5185 13679 5219
rect 18797 5185 18831 5219
rect 19625 5185 19659 5219
rect 21005 5185 21039 5219
rect 22477 5185 22511 5219
rect 23397 5185 23431 5219
rect 25789 5185 25823 5219
rect 28089 5185 28123 5219
rect 28365 5185 28399 5219
rect 30757 5185 30791 5219
rect 32781 5185 32815 5219
rect 33517 5185 33551 5219
rect 34621 5185 34655 5219
rect 35265 5185 35299 5219
rect 36369 5185 36403 5219
rect 36553 5185 36587 5219
rect 37565 5185 37599 5219
rect 39037 5185 39071 5219
rect 39681 5185 39715 5219
rect 40417 5185 40451 5219
rect 42717 5185 42751 5219
rect 43821 5185 43855 5219
rect 44649 5185 44683 5219
rect 56517 5185 56551 5219
rect 58081 5185 58115 5219
rect 1777 5117 1811 5151
rect 14289 5117 14323 5151
rect 19073 5117 19107 5151
rect 21281 5117 21315 5151
rect 22753 5117 22787 5151
rect 25605 5117 25639 5151
rect 30849 5117 30883 5151
rect 31033 5117 31067 5151
rect 32965 5117 32999 5151
rect 39221 5117 39255 5151
rect 10425 5049 10459 5083
rect 14565 5049 14599 5083
rect 17785 5049 17819 5083
rect 34805 5049 34839 5083
rect 37749 5049 37783 5083
rect 44005 5049 44039 5083
rect 14749 4981 14783 5015
rect 17325 4981 17359 5015
rect 24777 4981 24811 5015
rect 27445 4981 27479 5015
rect 32321 4981 32355 5015
rect 44741 4981 44775 5015
rect 58265 4981 58299 5015
rect 10609 4777 10643 4811
rect 11621 4777 11655 4811
rect 12817 4777 12851 4811
rect 18153 4777 18187 4811
rect 21005 4777 21039 4811
rect 22017 4777 22051 4811
rect 40969 4777 41003 4811
rect 41705 4777 41739 4811
rect 45385 4777 45419 4811
rect 47593 4777 47627 4811
rect 58081 4777 58115 4811
rect 9689 4709 9723 4743
rect 16221 4709 16255 4743
rect 21833 4709 21867 4743
rect 22477 4709 22511 4743
rect 39129 4709 39163 4743
rect 43269 4709 43303 4743
rect 44189 4709 44223 4743
rect 48329 4709 48363 4743
rect 8585 4641 8619 4675
rect 10793 4641 10827 4675
rect 10885 4641 10919 4675
rect 10977 4641 11011 4675
rect 11797 4641 11831 4675
rect 11897 4641 11931 4675
rect 18797 4641 18831 4675
rect 20177 4641 20211 4675
rect 22937 4641 22971 4675
rect 23121 4641 23155 4675
rect 25053 4641 25087 4675
rect 25145 4641 25179 4675
rect 32137 4641 32171 4675
rect 38393 4641 38427 4675
rect 57345 4641 57379 4675
rect 1593 4573 1627 4607
rect 9413 4573 9447 4607
rect 11069 4573 11103 4607
rect 11989 4573 12023 4607
rect 12081 4573 12115 4607
rect 12725 4573 12759 4607
rect 17049 4573 17083 4607
rect 19901 4573 19935 4607
rect 20913 4573 20947 4607
rect 22845 4573 22879 4607
rect 24961 4573 24995 4607
rect 26617 4573 26651 4607
rect 29009 4573 29043 4607
rect 30297 4573 30331 4607
rect 32321 4573 32355 4607
rect 33609 4573 33643 4607
rect 34897 4573 34931 4607
rect 36093 4573 36127 4607
rect 37197 4573 37231 4607
rect 38209 4573 38243 4607
rect 40877 4573 40911 4607
rect 47409 4573 47443 4607
rect 48145 4573 48179 4607
rect 57989 4573 58023 4607
rect 58173 4573 58207 4607
rect 1869 4505 1903 4539
rect 7481 4505 7515 4539
rect 8401 4505 8435 4539
rect 14657 4505 14691 4539
rect 16037 4505 16071 4539
rect 17325 4505 17359 4539
rect 18613 4505 18647 4539
rect 21557 4505 21591 4539
rect 27721 4505 27755 4539
rect 30564 4505 30598 4539
rect 35173 4505 35207 4539
rect 36369 4505 36403 4539
rect 37473 4505 37507 4539
rect 38945 4505 38979 4539
rect 40141 4505 40175 4539
rect 41613 4505 41647 4539
rect 42349 4505 42383 4539
rect 42533 4505 42567 4539
rect 43085 4505 43119 4539
rect 44005 4505 44039 4539
rect 45293 4505 45327 4539
rect 46029 4505 46063 4539
rect 46765 4505 46799 4539
rect 56609 4505 56643 4539
rect 7573 4437 7607 4471
rect 9873 4437 9907 4471
rect 14749 4437 14783 4471
rect 18521 4437 18555 4471
rect 19533 4437 19567 4471
rect 19993 4437 20027 4471
rect 24593 4437 24627 4471
rect 27077 4437 27111 4471
rect 28365 4437 28399 4471
rect 29101 4437 29135 4471
rect 31677 4437 31711 4471
rect 32505 4437 32539 4471
rect 33701 4437 33735 4471
rect 40233 4437 40267 4471
rect 46121 4437 46155 4471
rect 46857 4437 46891 4471
rect 23397 4233 23431 4267
rect 25329 4233 25363 4267
rect 27537 4233 27571 4267
rect 29653 4233 29687 4267
rect 7297 4165 7331 4199
rect 8033 4165 8067 4199
rect 12541 4165 12575 4199
rect 24216 4165 24250 4199
rect 28457 4165 28491 4199
rect 30573 4165 30607 4199
rect 32413 4165 32447 4199
rect 33793 4165 33827 4199
rect 35081 4165 35115 4199
rect 38485 4165 38519 4199
rect 40693 4165 40727 4199
rect 46857 4165 46891 4199
rect 48605 4165 48639 4199
rect 1593 4097 1627 4131
rect 8769 4097 8803 4131
rect 8953 4097 8987 4131
rect 10701 4097 10735 4131
rect 12357 4097 12391 4131
rect 13277 4097 13311 4131
rect 14933 4097 14967 4131
rect 15853 4097 15887 4131
rect 16865 4097 16899 4131
rect 17785 4097 17819 4131
rect 19073 4097 19107 4131
rect 19165 4097 19199 4131
rect 20085 4097 20119 4131
rect 21005 4097 21039 4131
rect 22017 4097 22051 4131
rect 22284 4097 22318 4131
rect 23949 4097 23983 4131
rect 25789 4097 25823 4131
rect 28641 4097 28675 4131
rect 31585 4097 31619 4131
rect 33609 4097 33643 4131
rect 33877 4097 33911 4131
rect 34001 4097 34035 4131
rect 34713 4097 34747 4131
rect 35817 4097 35851 4131
rect 36001 4097 36035 4131
rect 36185 4097 36219 4131
rect 36277 4097 36311 4131
rect 37473 4097 37507 4131
rect 39221 4097 39255 4131
rect 39957 4097 39991 4131
rect 41613 4097 41647 4131
rect 42625 4097 42659 4131
rect 43269 4097 43303 4131
rect 43637 4097 43671 4131
rect 43821 4097 43855 4131
rect 45293 4097 45327 4131
rect 45385 4097 45419 4131
rect 45661 4097 45695 4131
rect 45937 4097 45971 4131
rect 46121 4097 46155 4131
rect 47869 4097 47903 4131
rect 55413 4097 55447 4131
rect 55597 4097 55631 4131
rect 56313 4097 56347 4131
rect 58081 4097 58115 4131
rect 1777 4029 1811 4063
rect 7481 4029 7515 4063
rect 9413 4029 9447 4063
rect 10333 4029 10367 4063
rect 10517 4029 10551 4063
rect 10609 4029 10643 4063
rect 10793 4029 10827 4063
rect 12725 4029 12759 4063
rect 14013 4029 14047 4063
rect 16129 4029 16163 4063
rect 17141 4029 17175 4063
rect 18061 4029 18095 4063
rect 18889 4029 18923 4063
rect 18981 4029 19015 4063
rect 20177 4029 20211 4063
rect 20361 4029 20395 4063
rect 21281 4029 21315 4063
rect 25973 4029 26007 4063
rect 27629 4029 27663 4063
rect 27721 4029 27755 4063
rect 29745 4029 29779 4063
rect 29837 4029 29871 4063
rect 37657 4029 37691 4063
rect 41797 4029 41831 4063
rect 43361 4029 43395 4063
rect 48789 4029 48823 4063
rect 55505 4029 55539 4063
rect 56057 4029 56091 4063
rect 8217 3961 8251 3995
rect 9689 3961 9723 3995
rect 14289 3961 14323 3995
rect 15209 3961 15243 3995
rect 15393 3961 15427 3995
rect 34161 3961 34195 3995
rect 9873 3893 9907 3927
rect 13461 3893 13495 3927
rect 14473 3893 14507 3927
rect 18705 3893 18739 3927
rect 19717 3893 19751 3927
rect 27169 3893 27203 3927
rect 28825 3893 28859 3927
rect 29285 3893 29319 3927
rect 30665 3893 30699 3927
rect 31677 3893 31711 3927
rect 32505 3893 32539 3927
rect 38577 3893 38611 3927
rect 39313 3893 39347 3927
rect 40049 3893 40083 3927
rect 40785 3893 40819 3927
rect 44925 3893 44959 3927
rect 46949 3893 46983 3927
rect 47961 3893 47995 3927
rect 57437 3893 57471 3927
rect 58265 3893 58299 3927
rect 7021 3689 7055 3723
rect 20821 3689 20855 3723
rect 22201 3689 22235 3723
rect 40233 3689 40267 3723
rect 44189 3689 44223 3723
rect 48053 3689 48087 3723
rect 49709 3689 49743 3723
rect 51273 3689 51307 3723
rect 52745 3689 52779 3723
rect 53481 3689 53515 3723
rect 6285 3621 6319 3655
rect 7849 3621 7883 3655
rect 9689 3621 9723 3655
rect 11437 3621 11471 3655
rect 12357 3621 12391 3655
rect 12541 3621 12575 3655
rect 13645 3621 13679 3655
rect 15025 3621 15059 3655
rect 22017 3621 22051 3655
rect 24593 3621 24627 3655
rect 27169 3621 27203 3655
rect 38669 3621 38703 3655
rect 39497 3621 39531 3655
rect 50629 3621 50663 3655
rect 52101 3621 52135 3655
rect 54309 3621 54343 3655
rect 9873 3553 9907 3587
rect 9965 3553 9999 3587
rect 10149 3553 10183 3587
rect 13277 3553 13311 3587
rect 13737 3553 13771 3587
rect 14749 3553 14783 3587
rect 15945 3553 15979 3587
rect 18705 3553 18739 3587
rect 19441 3553 19475 3587
rect 21741 3553 21775 3587
rect 23029 3553 23063 3587
rect 25053 3553 25087 3587
rect 25145 3553 25179 3587
rect 27721 3553 27755 3587
rect 32045 3553 32079 3587
rect 35081 3553 35115 3587
rect 36001 3553 36035 3587
rect 41153 3553 41187 3587
rect 41889 3553 41923 3587
rect 42625 3553 42659 3587
rect 56885 3553 56919 3587
rect 1593 3485 1627 3519
rect 6929 3485 6963 3519
rect 8401 3485 8435 3519
rect 10057 3485 10091 3519
rect 12081 3485 12115 3519
rect 15669 3485 15703 3519
rect 16589 3485 16623 3519
rect 16865 3485 16899 3519
rect 17509 3485 17543 3519
rect 18429 3485 18463 3519
rect 19708 3485 19742 3519
rect 23581 3485 23615 3519
rect 25789 3485 25823 3519
rect 26056 3485 26090 3519
rect 28549 3485 28583 3519
rect 28687 3485 28721 3519
rect 30297 3485 30331 3519
rect 32312 3485 32346 3519
rect 34069 3485 34103 3519
rect 34897 3485 34931 3519
rect 35817 3485 35851 3519
rect 36737 3485 36771 3519
rect 38117 3485 38151 3519
rect 38490 3485 38524 3519
rect 39313 3485 39347 3519
rect 40141 3485 40175 3519
rect 40969 3485 41003 3519
rect 42533 3485 42567 3519
rect 42901 3485 42935 3519
rect 42993 3485 43027 3519
rect 43545 3485 43579 3519
rect 43693 3485 43727 3519
rect 44010 3485 44044 3519
rect 45201 3485 45235 3519
rect 45661 3485 45695 3519
rect 45753 3485 45787 3519
rect 46029 3485 46063 3519
rect 46305 3485 46339 3519
rect 46581 3485 46615 3519
rect 48881 3485 48915 3519
rect 51089 3485 51123 3519
rect 52561 3485 52595 3519
rect 53297 3485 53331 3519
rect 56057 3485 56091 3519
rect 56241 3485 56275 3519
rect 1869 3417 1903 3451
rect 6101 3417 6135 3451
rect 7665 3417 7699 3451
rect 11161 3417 11195 3451
rect 17785 3417 17819 3451
rect 22753 3417 22787 3451
rect 23857 3417 23891 3451
rect 28365 3417 28399 3451
rect 28917 3417 28951 3451
rect 30573 3417 30607 3451
rect 31401 3417 31435 3451
rect 34253 3417 34287 3451
rect 37013 3417 37047 3451
rect 38301 3417 38335 3451
rect 38393 3417 38427 3451
rect 43821 3417 43855 3451
rect 43913 3417 43947 3451
rect 47225 3417 47259 3451
rect 47961 3417 47995 3451
rect 48697 3417 48731 3451
rect 49433 3417 49467 3451
rect 50445 3417 50479 3451
rect 51917 3417 51951 3451
rect 54125 3417 54159 3451
rect 56425 3417 56459 3451
rect 57130 3417 57164 3451
rect 8493 3349 8527 3383
rect 11621 3349 11655 3383
rect 15209 3349 15243 3383
rect 24961 3349 24995 3383
rect 28733 3349 28767 3383
rect 31493 3349 31527 3383
rect 33425 3349 33459 3383
rect 47317 3349 47351 3383
rect 58265 3349 58299 3383
rect 5917 3145 5951 3179
rect 6929 3145 6963 3179
rect 8401 3145 8435 3179
rect 9137 3145 9171 3179
rect 11161 3145 11195 3179
rect 12725 3145 12759 3179
rect 42809 3145 42843 3179
rect 46949 3145 46983 3179
rect 47961 3145 47995 3179
rect 48697 3145 48731 3179
rect 49801 3145 49835 3179
rect 50537 3145 50571 3179
rect 52009 3145 52043 3179
rect 53849 3145 53883 3179
rect 55321 3145 55355 3179
rect 58265 3145 58299 3179
rect 5825 3077 5859 3111
rect 10701 3077 10735 3111
rect 11897 3077 11931 3111
rect 12081 3077 12115 3111
rect 13369 3077 13403 3111
rect 15209 3077 15243 3111
rect 18429 3077 18463 3111
rect 19340 3077 19374 3111
rect 28816 3077 28850 3111
rect 34437 3077 34471 3111
rect 36277 3077 36311 3111
rect 40693 3077 40727 3111
rect 41613 3077 41647 3111
rect 53021 3077 53055 3111
rect 55229 3077 55263 3111
rect 56609 3077 56643 3111
rect 58173 3077 58207 3111
rect 6837 3009 6871 3043
rect 7573 3009 7607 3043
rect 8309 3009 8343 3043
rect 9045 3009 9079 3043
rect 10057 3009 10091 3043
rect 10149 3009 10183 3043
rect 12633 3009 12667 3043
rect 14013 3009 14047 3043
rect 14933 3009 14967 3043
rect 15853 3009 15887 3043
rect 17233 3009 17267 3043
rect 18153 3009 18187 3043
rect 19073 3009 19107 3043
rect 21005 3009 21039 3043
rect 22569 3009 22603 3043
rect 23489 3009 23523 3043
rect 23756 3009 23790 3043
rect 26157 3009 26191 3043
rect 27169 3009 27203 3043
rect 28549 3009 28583 3043
rect 30849 3009 30883 3043
rect 32321 3009 32355 3043
rect 33241 3009 33275 3043
rect 34161 3009 34195 3043
rect 35081 3009 35115 3043
rect 36001 3009 36035 3043
rect 37473 3009 37507 3043
rect 38393 3009 38427 3043
rect 39313 3009 39347 3043
rect 40325 3009 40359 3043
rect 41245 3009 41279 3043
rect 42717 3009 42751 3043
rect 44557 3009 44591 3043
rect 44649 3009 44683 3043
rect 44925 3009 44959 3043
rect 45201 3009 45235 3043
rect 45477 3009 45511 3043
rect 46121 3009 46155 3043
rect 46857 3009 46891 3043
rect 47777 3009 47811 3043
rect 48605 3009 48639 3043
rect 49525 3009 49559 3043
rect 50353 3009 50387 3043
rect 51181 3009 51215 3043
rect 51825 3009 51859 3043
rect 53757 3009 53791 3043
rect 54493 3009 54527 3043
rect 54677 3009 54711 3043
rect 56425 3009 56459 3043
rect 57161 3009 57195 3043
rect 57253 3009 57287 3043
rect 9873 2941 9907 2975
rect 9965 2941 9999 2975
rect 14197 2941 14231 2975
rect 16129 2941 16163 2975
rect 17509 2941 17543 2975
rect 21281 2941 21315 2975
rect 22845 2941 22879 2975
rect 26341 2941 26375 2975
rect 27353 2941 27387 2975
rect 31033 2941 31067 2975
rect 32505 2941 32539 2975
rect 33425 2941 33459 2975
rect 35265 2941 35299 2975
rect 37657 2941 37691 2975
rect 38577 2941 38611 2975
rect 39497 2941 39531 2975
rect 57437 2941 57471 2975
rect 7757 2873 7791 2907
rect 9689 2873 9723 2907
rect 10977 2873 11011 2907
rect 13553 2873 13587 2907
rect 24869 2873 24903 2907
rect 29929 2873 29963 2907
rect 44189 2873 44223 2907
rect 20453 2805 20487 2839
rect 25697 2805 25731 2839
rect 46213 2805 46247 2839
rect 51273 2805 51307 2839
rect 53113 2805 53147 2839
rect 5917 2601 5951 2635
rect 10609 2601 10643 2635
rect 17049 2601 17083 2635
rect 22109 2601 22143 2635
rect 24777 2601 24811 2635
rect 41153 2601 41187 2635
rect 44189 2601 44223 2635
rect 45753 2601 45787 2635
rect 46489 2601 46523 2635
rect 50537 2601 50571 2635
rect 51457 2601 51491 2635
rect 53113 2601 53147 2635
rect 58265 2601 58299 2635
rect 8585 2533 8619 2567
rect 10425 2533 10459 2567
rect 12265 2533 12299 2567
rect 13737 2533 13771 2567
rect 10149 2465 10183 2499
rect 22937 2465 22971 2499
rect 33425 2465 33459 2499
rect 36001 2465 36035 2499
rect 38577 2465 38611 2499
rect 40233 2465 40267 2499
rect 48973 2465 49007 2499
rect 54769 2465 54803 2499
rect 1593 2397 1627 2431
rect 1869 2397 1903 2431
rect 5089 2397 5123 2431
rect 6929 2397 6963 2431
rect 7665 2397 7699 2431
rect 9505 2397 9539 2431
rect 13553 2397 13587 2431
rect 14473 2397 14507 2431
rect 14933 2397 14967 2431
rect 15853 2397 15887 2431
rect 17509 2397 17543 2431
rect 18429 2397 18463 2431
rect 19625 2397 19659 2431
rect 20085 2397 20119 2431
rect 21005 2397 21039 2431
rect 22017 2397 22051 2431
rect 22661 2397 22695 2431
rect 23581 2397 23615 2431
rect 25237 2397 25271 2431
rect 26157 2397 26191 2431
rect 27169 2397 27203 2431
rect 28733 2397 28767 2431
rect 30205 2397 30239 2431
rect 31125 2397 31159 2431
rect 32321 2397 32355 2431
rect 33241 2397 33275 2431
rect 34897 2397 34931 2431
rect 35817 2397 35851 2431
rect 37473 2397 37507 2431
rect 38393 2397 38427 2431
rect 40049 2397 40083 2431
rect 41061 2397 41095 2431
rect 42625 2397 42659 2431
rect 43545 2397 43579 2431
rect 43693 2397 43727 2431
rect 44051 2397 44085 2431
rect 45201 2397 45235 2431
rect 45385 2397 45419 2431
rect 45574 2397 45608 2431
rect 48697 2397 48731 2431
rect 52929 2397 52963 2431
rect 56333 2397 56367 2431
rect 57069 2397 57103 2431
rect 58173 2397 58207 2431
rect 5825 2329 5859 2363
rect 8401 2329 8435 2363
rect 9689 2329 9723 2363
rect 12081 2329 12115 2363
rect 12817 2329 12851 2363
rect 15209 2329 15243 2363
rect 16129 2329 16163 2363
rect 17785 2329 17819 2363
rect 18705 2329 18739 2363
rect 20361 2329 20395 2363
rect 21281 2329 21315 2363
rect 23857 2329 23891 2363
rect 25513 2329 25547 2363
rect 26433 2329 26467 2363
rect 27445 2329 27479 2363
rect 29009 2329 29043 2363
rect 30481 2329 30515 2363
rect 31401 2329 31435 2363
rect 32597 2329 32631 2363
rect 35173 2329 35207 2363
rect 37749 2329 37783 2363
rect 42901 2329 42935 2363
rect 43821 2329 43855 2363
rect 43913 2329 43947 2363
rect 45477 2329 45511 2363
rect 46397 2329 46431 2363
rect 47869 2329 47903 2363
rect 50445 2329 50479 2363
rect 51365 2329 51399 2363
rect 54033 2329 54067 2363
rect 55597 2329 55631 2363
rect 57345 2329 57379 2363
rect 5181 2261 5215 2295
rect 7021 2261 7055 2295
rect 7757 2261 7791 2295
rect 12909 2261 12943 2295
rect 28089 2261 28123 2295
rect 47961 2261 47995 2295
rect 55689 2261 55723 2295
rect 56425 2261 56459 2295
<< metal1 >>
rect 1104 61498 58880 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 58880 61498
rect 1104 61424 58880 61446
rect 1949 61319 2007 61325
rect 1949 61285 1961 61319
rect 1995 61316 2007 61319
rect 6178 61316 6184 61328
rect 1995 61288 6184 61316
rect 1995 61285 2007 61288
rect 1949 61279 2007 61285
rect 6178 61276 6184 61288
rect 6236 61276 6242 61328
rect 9677 61319 9735 61325
rect 9677 61285 9689 61319
rect 9723 61316 9735 61319
rect 17126 61316 17132 61328
rect 9723 61288 17132 61316
rect 9723 61285 9735 61288
rect 9677 61279 9735 61285
rect 17126 61276 17132 61288
rect 17184 61276 17190 61328
rect 20717 61319 20775 61325
rect 20717 61285 20729 61319
rect 20763 61316 20775 61319
rect 21726 61316 21732 61328
rect 20763 61288 21732 61316
rect 20763 61285 20775 61288
rect 20717 61279 20775 61285
rect 21726 61276 21732 61288
rect 21784 61276 21790 61328
rect 2774 61208 2780 61260
rect 2832 61208 2838 61260
rect 44450 61208 44456 61260
rect 44508 61248 44514 61260
rect 49513 61251 49571 61257
rect 49513 61248 49525 61251
rect 44508 61220 49525 61248
rect 44508 61208 44514 61220
rect 49513 61217 49525 61220
rect 49559 61217 49571 61251
rect 49513 61211 49571 61217
rect 56778 61208 56784 61260
rect 56836 61248 56842 61260
rect 56836 61220 58112 61248
rect 56836 61208 56842 61220
rect 2501 61183 2559 61189
rect 2501 61149 2513 61183
rect 2547 61180 2559 61183
rect 2792 61180 2820 61208
rect 2547 61152 2820 61180
rect 4341 61183 4399 61189
rect 2547 61149 2559 61152
rect 2501 61143 2559 61149
rect 4341 61149 4353 61183
rect 4387 61180 4399 61183
rect 4614 61180 4620 61192
rect 4387 61152 4620 61180
rect 4387 61149 4399 61152
rect 4341 61143 4399 61149
rect 4614 61140 4620 61152
rect 4672 61140 4678 61192
rect 5074 61180 5080 61192
rect 5035 61152 5080 61180
rect 5074 61140 5080 61152
rect 5132 61140 5138 61192
rect 5810 61180 5816 61192
rect 5771 61152 5816 61180
rect 5810 61140 5816 61152
rect 5868 61140 5874 61192
rect 6730 61180 6736 61192
rect 6691 61152 6736 61180
rect 6730 61140 6736 61152
rect 6788 61140 6794 61192
rect 7558 61180 7564 61192
rect 7519 61152 7564 61180
rect 7558 61140 7564 61152
rect 7616 61140 7622 61192
rect 7834 61180 7840 61192
rect 7795 61152 7840 61180
rect 7834 61140 7840 61152
rect 7892 61140 7898 61192
rect 9493 61183 9551 61189
rect 9493 61149 9505 61183
rect 9539 61180 9551 61183
rect 9674 61180 9680 61192
rect 9539 61152 9680 61180
rect 9539 61149 9551 61152
rect 9493 61143 9551 61149
rect 9674 61140 9680 61152
rect 9732 61140 9738 61192
rect 10226 61180 10232 61192
rect 10187 61152 10232 61180
rect 10226 61140 10232 61152
rect 10284 61140 10290 61192
rect 10965 61183 11023 61189
rect 10965 61149 10977 61183
rect 11011 61180 11023 61183
rect 11146 61180 11152 61192
rect 11011 61152 11152 61180
rect 11011 61149 11023 61152
rect 10965 61143 11023 61149
rect 11146 61140 11152 61152
rect 11204 61140 11210 61192
rect 12434 61180 12440 61192
rect 12395 61152 12440 61180
rect 12434 61140 12440 61152
rect 12492 61140 12498 61192
rect 13262 61180 13268 61192
rect 13223 61152 13268 61180
rect 13262 61140 13268 61152
rect 13320 61140 13326 61192
rect 14366 61180 14372 61192
rect 14327 61152 14372 61180
rect 14366 61140 14372 61152
rect 14424 61140 14430 61192
rect 15378 61180 15384 61192
rect 15339 61152 15384 61180
rect 15378 61140 15384 61152
rect 15436 61140 15442 61192
rect 16114 61180 16120 61192
rect 16075 61152 16120 61180
rect 16114 61140 16120 61152
rect 16172 61140 16178 61192
rect 17218 61180 17224 61192
rect 17179 61152 17224 61180
rect 17218 61140 17224 61152
rect 17276 61140 17282 61192
rect 17954 61180 17960 61192
rect 17915 61152 17960 61180
rect 17954 61140 17960 61152
rect 18012 61140 18018 61192
rect 18690 61180 18696 61192
rect 18651 61152 18696 61180
rect 18690 61140 18696 61152
rect 18748 61140 18754 61192
rect 19794 61180 19800 61192
rect 19755 61152 19800 61180
rect 19794 61140 19800 61152
rect 19852 61140 19858 61192
rect 20533 61183 20591 61189
rect 20533 61149 20545 61183
rect 20579 61180 20591 61183
rect 20714 61180 20720 61192
rect 20579 61152 20720 61180
rect 20579 61149 20591 61152
rect 20533 61143 20591 61149
rect 20714 61140 20720 61152
rect 20772 61140 20778 61192
rect 21266 61180 21272 61192
rect 21227 61152 21272 61180
rect 21266 61140 21272 61152
rect 21324 61140 21330 61192
rect 22370 61180 22376 61192
rect 22331 61152 22376 61180
rect 22370 61140 22376 61152
rect 22428 61140 22434 61192
rect 23106 61180 23112 61192
rect 23067 61152 23112 61180
rect 23106 61140 23112 61152
rect 23164 61140 23170 61192
rect 23842 61180 23848 61192
rect 23803 61152 23848 61180
rect 23842 61140 23848 61152
rect 23900 61140 23906 61192
rect 25130 61140 25136 61192
rect 25188 61180 25194 61192
rect 25317 61183 25375 61189
rect 25317 61180 25329 61183
rect 25188 61152 25329 61180
rect 25188 61140 25194 61152
rect 25317 61149 25329 61152
rect 25363 61149 25375 61183
rect 26050 61180 26056 61192
rect 26011 61152 26056 61180
rect 25317 61143 25375 61149
rect 26050 61140 26056 61152
rect 26108 61140 26114 61192
rect 27522 61180 27528 61192
rect 27483 61152 27528 61180
rect 27522 61140 27528 61152
rect 27580 61140 27586 61192
rect 28350 61180 28356 61192
rect 28311 61152 28356 61180
rect 28350 61140 28356 61152
rect 28408 61140 28414 61192
rect 28994 61140 29000 61192
rect 29052 61180 29058 61192
rect 29825 61183 29883 61189
rect 29825 61180 29837 61183
rect 29052 61152 29837 61180
rect 29052 61140 29058 61152
rect 29825 61149 29837 61152
rect 29871 61149 29883 61183
rect 29825 61143 29883 61149
rect 31018 61140 31024 61192
rect 31076 61180 31082 61192
rect 31205 61183 31263 61189
rect 31205 61180 31217 61183
rect 31076 61152 31217 61180
rect 31076 61140 31082 61152
rect 31205 61149 31217 61152
rect 31251 61149 31263 61183
rect 31205 61143 31263 61149
rect 31754 61140 31760 61192
rect 31812 61180 31818 61192
rect 32401 61183 32459 61189
rect 32401 61180 32413 61183
rect 31812 61152 32413 61180
rect 31812 61140 31818 61152
rect 32401 61149 32413 61152
rect 32447 61149 32459 61183
rect 32401 61143 32459 61149
rect 32490 61140 32496 61192
rect 32548 61180 32554 61192
rect 33045 61183 33103 61189
rect 33045 61180 33057 61183
rect 32548 61152 33057 61180
rect 32548 61140 32554 61152
rect 33045 61149 33057 61152
rect 33091 61149 33103 61183
rect 33045 61143 33103 61149
rect 33226 61140 33232 61192
rect 33284 61180 33290 61192
rect 33781 61183 33839 61189
rect 33781 61180 33793 61183
rect 33284 61152 33793 61180
rect 33284 61140 33290 61152
rect 33781 61149 33793 61152
rect 33827 61149 33839 61183
rect 33781 61143 33839 61149
rect 34698 61140 34704 61192
rect 34756 61180 34762 61192
rect 34977 61183 35035 61189
rect 34977 61180 34989 61183
rect 34756 61152 34989 61180
rect 34756 61140 34762 61152
rect 34977 61149 34989 61152
rect 35023 61149 35035 61183
rect 34977 61143 35035 61149
rect 35894 61140 35900 61192
rect 35952 61180 35958 61192
rect 35952 61152 35997 61180
rect 35952 61140 35958 61152
rect 37274 61140 37280 61192
rect 37332 61180 37338 61192
rect 37553 61183 37611 61189
rect 37553 61180 37565 61183
rect 37332 61152 37565 61180
rect 37332 61140 37338 61152
rect 37553 61149 37565 61152
rect 37599 61149 37611 61183
rect 37553 61143 37611 61149
rect 37642 61140 37648 61192
rect 37700 61180 37706 61192
rect 38289 61183 38347 61189
rect 38289 61180 38301 61183
rect 37700 61152 38301 61180
rect 37700 61140 37706 61152
rect 38289 61149 38301 61152
rect 38335 61149 38347 61183
rect 38289 61143 38347 61149
rect 38378 61140 38384 61192
rect 38436 61180 38442 61192
rect 39025 61183 39083 61189
rect 39025 61180 39037 61183
rect 38436 61152 39037 61180
rect 38436 61140 38442 61152
rect 39025 61149 39037 61152
rect 39071 61149 39083 61183
rect 39025 61143 39083 61149
rect 40034 61140 40040 61192
rect 40092 61180 40098 61192
rect 40773 61183 40831 61189
rect 40773 61180 40785 61183
rect 40092 61152 40785 61180
rect 40092 61140 40098 61152
rect 40773 61149 40785 61152
rect 40819 61149 40831 61183
rect 40773 61143 40831 61149
rect 40954 61140 40960 61192
rect 41012 61180 41018 61192
rect 41601 61183 41659 61189
rect 41601 61180 41613 61183
rect 41012 61152 41613 61180
rect 41012 61140 41018 61152
rect 41601 61149 41613 61152
rect 41647 61149 41659 61183
rect 41601 61143 41659 61149
rect 42058 61140 42064 61192
rect 42116 61180 42122 61192
rect 42705 61183 42763 61189
rect 42705 61180 42717 61183
rect 42116 61152 42717 61180
rect 42116 61140 42122 61152
rect 42705 61149 42717 61152
rect 42751 61149 42763 61183
rect 42705 61143 42763 61149
rect 42794 61140 42800 61192
rect 42852 61180 42858 61192
rect 43625 61183 43683 61189
rect 43625 61180 43637 61183
rect 42852 61152 43637 61180
rect 42852 61140 42858 61152
rect 43625 61149 43637 61152
rect 43671 61149 43683 61183
rect 43625 61143 43683 61149
rect 44174 61140 44180 61192
rect 44232 61180 44238 61192
rect 44361 61183 44419 61189
rect 44361 61180 44373 61183
rect 44232 61152 44373 61180
rect 44232 61140 44238 61152
rect 44361 61149 44373 61152
rect 44407 61149 44419 61183
rect 44361 61143 44419 61149
rect 44542 61140 44548 61192
rect 44600 61180 44606 61192
rect 45281 61183 45339 61189
rect 45281 61180 45293 61183
rect 44600 61152 45293 61180
rect 44600 61140 44606 61152
rect 45281 61149 45293 61152
rect 45327 61149 45339 61183
rect 45281 61143 45339 61149
rect 45554 61140 45560 61192
rect 45612 61180 45618 61192
rect 46017 61183 46075 61189
rect 46017 61180 46029 61183
rect 45612 61152 46029 61180
rect 45612 61140 45618 61152
rect 46017 61149 46029 61152
rect 46063 61149 46075 61183
rect 46017 61143 46075 61149
rect 46106 61140 46112 61192
rect 46164 61180 46170 61192
rect 46753 61183 46811 61189
rect 46753 61180 46765 61183
rect 46164 61152 46765 61180
rect 46164 61140 46170 61152
rect 46753 61149 46765 61152
rect 46799 61149 46811 61183
rect 46753 61143 46811 61149
rect 47210 61140 47216 61192
rect 47268 61180 47274 61192
rect 47857 61183 47915 61189
rect 47857 61180 47869 61183
rect 47268 61152 47869 61180
rect 47268 61140 47274 61152
rect 47857 61149 47869 61152
rect 47903 61149 47915 61183
rect 47857 61143 47915 61149
rect 48314 61140 48320 61192
rect 48372 61180 48378 61192
rect 48593 61183 48651 61189
rect 48593 61180 48605 61183
rect 48372 61152 48605 61180
rect 48372 61140 48378 61152
rect 48593 61149 48605 61152
rect 48639 61149 48651 61183
rect 48593 61143 48651 61149
rect 48682 61140 48688 61192
rect 48740 61180 48746 61192
rect 49329 61183 49387 61189
rect 49329 61180 49341 61183
rect 48740 61152 49341 61180
rect 48740 61140 48746 61152
rect 49329 61149 49341 61152
rect 49375 61149 49387 61183
rect 51074 61180 51080 61192
rect 51035 61152 51080 61180
rect 49329 61143 49387 61149
rect 51074 61140 51080 61152
rect 51132 61140 51138 61192
rect 51994 61180 52000 61192
rect 51955 61152 52000 61180
rect 51994 61140 52000 61152
rect 52052 61140 52058 61192
rect 53190 61180 53196 61192
rect 53151 61152 53196 61180
rect 53190 61140 53196 61152
rect 53248 61140 53254 61192
rect 54202 61180 54208 61192
rect 54163 61152 54208 61180
rect 54202 61140 54208 61152
rect 54260 61140 54266 61192
rect 56134 61180 56140 61192
rect 56095 61152 56140 61180
rect 56134 61140 56140 61152
rect 56192 61140 56198 61192
rect 57149 61183 57207 61189
rect 57149 61149 57161 61183
rect 57195 61180 57207 61183
rect 57514 61180 57520 61192
rect 57195 61152 57520 61180
rect 57195 61149 57207 61152
rect 57149 61143 57207 61149
rect 57514 61140 57520 61152
rect 57572 61140 57578 61192
rect 58084 61189 58112 61220
rect 58069 61183 58127 61189
rect 58069 61149 58081 61183
rect 58115 61149 58127 61183
rect 58069 61143 58127 61149
rect 1670 61112 1676 61124
rect 1631 61084 1676 61112
rect 1670 61072 1676 61084
rect 1728 61072 1734 61124
rect 2777 61115 2835 61121
rect 2777 61081 2789 61115
rect 2823 61081 2835 61115
rect 2777 61075 2835 61081
rect 4525 61115 4583 61121
rect 4525 61081 4537 61115
rect 4571 61112 4583 61115
rect 4890 61112 4896 61124
rect 4571 61084 4896 61112
rect 4571 61081 4583 61084
rect 4525 61075 4583 61081
rect 2792 61044 2820 61075
rect 4890 61072 4896 61084
rect 4948 61072 4954 61124
rect 7650 61112 7656 61124
rect 5000 61084 7656 61112
rect 5000 61044 5028 61084
rect 7650 61072 7656 61084
rect 7708 61072 7714 61124
rect 13538 61112 13544 61124
rect 13499 61084 13544 61112
rect 13538 61072 13544 61084
rect 13596 61072 13602 61124
rect 15565 61115 15623 61121
rect 15565 61081 15577 61115
rect 15611 61112 15623 61115
rect 15654 61112 15660 61124
rect 15611 61084 15660 61112
rect 15611 61081 15623 61084
rect 15565 61075 15623 61081
rect 15654 61072 15660 61084
rect 15712 61072 15718 61124
rect 16301 61115 16359 61121
rect 16301 61081 16313 61115
rect 16347 61112 16359 61115
rect 16390 61112 16396 61124
rect 16347 61084 16396 61112
rect 16347 61081 16359 61084
rect 16301 61075 16359 61081
rect 16390 61072 16396 61084
rect 16448 61072 16454 61124
rect 18138 61112 18144 61124
rect 18099 61084 18144 61112
rect 18138 61072 18144 61084
rect 18196 61072 18202 61124
rect 19981 61115 20039 61121
rect 19981 61081 19993 61115
rect 20027 61112 20039 61115
rect 20346 61112 20352 61124
rect 20027 61084 20352 61112
rect 20027 61081 20039 61084
rect 19981 61075 20039 61081
rect 20346 61072 20352 61084
rect 20404 61072 20410 61124
rect 26421 61115 26479 61121
rect 26421 61081 26433 61115
rect 26467 61112 26479 61115
rect 31662 61112 31668 61124
rect 26467 61084 31668 61112
rect 26467 61081 26479 61084
rect 26421 61075 26479 61081
rect 31662 61072 31668 61084
rect 31720 61072 31726 61124
rect 37734 61112 37740 61124
rect 37695 61084 37740 61112
rect 37734 61072 37740 61084
rect 37792 61072 37798 61124
rect 39482 61072 39488 61124
rect 39540 61112 39546 61124
rect 40129 61115 40187 61121
rect 40129 61112 40141 61115
rect 39540 61084 40141 61112
rect 39540 61072 39546 61084
rect 40129 61081 40141 61084
rect 40175 61081 40187 61115
rect 46934 61112 46940 61124
rect 40129 61075 40187 61081
rect 42076 61084 46796 61112
rect 46895 61084 46940 61112
rect 42076 61056 42104 61084
rect 5166 61044 5172 61056
rect 2792 61016 5028 61044
rect 5127 61016 5172 61044
rect 5166 61004 5172 61016
rect 5224 61004 5230 61056
rect 5902 61044 5908 61056
rect 5863 61016 5908 61044
rect 5902 61004 5908 61016
rect 5960 61004 5966 61056
rect 6914 61004 6920 61056
rect 6972 61044 6978 61056
rect 7009 61047 7067 61053
rect 7009 61044 7021 61047
rect 6972 61016 7021 61044
rect 6972 61004 6978 61016
rect 7009 61013 7021 61016
rect 7055 61013 7067 61047
rect 10318 61044 10324 61056
rect 10279 61016 10324 61044
rect 7009 61007 7067 61013
rect 10318 61004 10324 61016
rect 10376 61004 10382 61056
rect 11057 61047 11115 61053
rect 11057 61013 11069 61047
rect 11103 61044 11115 61047
rect 11974 61044 11980 61056
rect 11103 61016 11980 61044
rect 11103 61013 11115 61016
rect 11057 61007 11115 61013
rect 11974 61004 11980 61016
rect 12032 61004 12038 61056
rect 12526 61044 12532 61056
rect 12487 61016 12532 61044
rect 12526 61004 12532 61016
rect 12584 61004 12590 61056
rect 14458 61044 14464 61056
rect 14419 61016 14464 61044
rect 14458 61004 14464 61016
rect 14516 61004 14522 61056
rect 16574 61004 16580 61056
rect 16632 61044 16638 61056
rect 17313 61047 17371 61053
rect 17313 61044 17325 61047
rect 16632 61016 17325 61044
rect 16632 61004 16638 61016
rect 17313 61013 17325 61016
rect 17359 61013 17371 61047
rect 17313 61007 17371 61013
rect 18506 61004 18512 61056
rect 18564 61044 18570 61056
rect 18785 61047 18843 61053
rect 18785 61044 18797 61047
rect 18564 61016 18797 61044
rect 18564 61004 18570 61016
rect 18785 61013 18797 61016
rect 18831 61013 18843 61047
rect 18785 61007 18843 61013
rect 20806 61004 20812 61056
rect 20864 61044 20870 61056
rect 21361 61047 21419 61053
rect 21361 61044 21373 61047
rect 20864 61016 21373 61044
rect 20864 61004 20870 61016
rect 21361 61013 21373 61016
rect 21407 61013 21419 61047
rect 21361 61007 21419 61013
rect 22278 61004 22284 61056
rect 22336 61044 22342 61056
rect 22465 61047 22523 61053
rect 22465 61044 22477 61047
rect 22336 61016 22477 61044
rect 22336 61004 22342 61016
rect 22465 61013 22477 61016
rect 22511 61013 22523 61047
rect 22465 61007 22523 61013
rect 22922 61004 22928 61056
rect 22980 61044 22986 61056
rect 23201 61047 23259 61053
rect 23201 61044 23213 61047
rect 22980 61016 23213 61044
rect 22980 61004 22986 61016
rect 23201 61013 23213 61016
rect 23247 61013 23259 61047
rect 23934 61044 23940 61056
rect 23895 61016 23940 61044
rect 23201 61007 23259 61013
rect 23934 61004 23940 61016
rect 23992 61004 23998 61056
rect 25130 61004 25136 61056
rect 25188 61044 25194 61056
rect 25409 61047 25467 61053
rect 25409 61044 25421 61047
rect 25188 61016 25421 61044
rect 25188 61004 25194 61016
rect 25409 61013 25421 61016
rect 25455 61013 25467 61047
rect 27614 61044 27620 61056
rect 27575 61016 27620 61044
rect 25409 61007 25467 61013
rect 27614 61004 27620 61016
rect 27672 61004 27678 61056
rect 28534 61044 28540 61056
rect 28495 61016 28540 61044
rect 28534 61004 28540 61016
rect 28592 61004 28598 61056
rect 29917 61047 29975 61053
rect 29917 61013 29929 61047
rect 29963 61044 29975 61047
rect 30006 61044 30012 61056
rect 29963 61016 30012 61044
rect 29963 61013 29975 61016
rect 29917 61007 29975 61013
rect 30006 61004 30012 61016
rect 30064 61004 30070 61056
rect 31018 61004 31024 61056
rect 31076 61044 31082 61056
rect 31297 61047 31355 61053
rect 31297 61044 31309 61047
rect 31076 61016 31309 61044
rect 31076 61004 31082 61016
rect 31297 61013 31309 61016
rect 31343 61013 31355 61047
rect 31297 61007 31355 61013
rect 31938 61004 31944 61056
rect 31996 61044 32002 61056
rect 32493 61047 32551 61053
rect 32493 61044 32505 61047
rect 31996 61016 32505 61044
rect 31996 61004 32002 61016
rect 32493 61013 32505 61016
rect 32539 61013 32551 61047
rect 33226 61044 33232 61056
rect 33187 61016 33232 61044
rect 32493 61007 32551 61013
rect 33226 61004 33232 61016
rect 33284 61004 33290 61056
rect 33318 61004 33324 61056
rect 33376 61044 33382 61056
rect 33965 61047 34023 61053
rect 33965 61044 33977 61047
rect 33376 61016 33977 61044
rect 33376 61004 33382 61016
rect 33965 61013 33977 61016
rect 34011 61013 34023 61047
rect 35066 61044 35072 61056
rect 35027 61016 35072 61044
rect 33965 61007 34023 61013
rect 35066 61004 35072 61016
rect 35124 61004 35130 61056
rect 35986 61044 35992 61056
rect 35947 61016 35992 61044
rect 35986 61004 35992 61016
rect 36044 61004 36050 61056
rect 37274 61004 37280 61056
rect 37332 61044 37338 61056
rect 38381 61047 38439 61053
rect 38381 61044 38393 61047
rect 37332 61016 38393 61044
rect 37332 61004 37338 61016
rect 38381 61013 38393 61016
rect 38427 61013 38439 61047
rect 38381 61007 38439 61013
rect 39117 61047 39175 61053
rect 39117 61013 39129 61047
rect 39163 61044 39175 61047
rect 39758 61044 39764 61056
rect 39163 61016 39764 61044
rect 39163 61013 39175 61016
rect 39117 61007 39175 61013
rect 39758 61004 39764 61016
rect 39816 61004 39822 61056
rect 40218 61044 40224 61056
rect 40179 61016 40224 61044
rect 40218 61004 40224 61016
rect 40276 61004 40282 61056
rect 40954 61044 40960 61056
rect 40915 61016 40960 61044
rect 40954 61004 40960 61016
rect 41012 61004 41018 61056
rect 41046 61004 41052 61056
rect 41104 61044 41110 61056
rect 41693 61047 41751 61053
rect 41693 61044 41705 61047
rect 41104 61016 41705 61044
rect 41104 61004 41110 61016
rect 41693 61013 41705 61016
rect 41739 61013 41751 61047
rect 41693 61007 41751 61013
rect 42058 61004 42064 61056
rect 42116 61004 42122 61056
rect 42794 61044 42800 61056
rect 42755 61016 42800 61044
rect 42794 61004 42800 61016
rect 42852 61004 42858 61056
rect 43714 61044 43720 61056
rect 43675 61016 43720 61044
rect 43714 61004 43720 61016
rect 43772 61004 43778 61056
rect 44266 61004 44272 61056
rect 44324 61044 44330 61056
rect 44453 61047 44511 61053
rect 44453 61044 44465 61047
rect 44324 61016 44465 61044
rect 44324 61004 44330 61016
rect 44453 61013 44465 61016
rect 44499 61013 44511 61047
rect 45370 61044 45376 61056
rect 45331 61016 45376 61044
rect 44453 61007 44511 61013
rect 45370 61004 45376 61016
rect 45428 61004 45434 61056
rect 46106 61044 46112 61056
rect 46067 61016 46112 61044
rect 46106 61004 46112 61016
rect 46164 61004 46170 61056
rect 46768 61044 46796 61084
rect 46934 61072 46940 61084
rect 46992 61072 46998 61124
rect 53469 61115 53527 61121
rect 53469 61112 53481 61115
rect 47044 61084 53481 61112
rect 47044 61044 47072 61084
rect 53469 61081 53481 61084
rect 53515 61081 53527 61115
rect 54386 61112 54392 61124
rect 54347 61084 54392 61112
rect 53469 61075 53527 61081
rect 54386 61072 54392 61084
rect 54444 61072 54450 61124
rect 56410 61112 56416 61124
rect 56371 61084 56416 61112
rect 56410 61072 56416 61084
rect 56468 61072 56474 61124
rect 47946 61044 47952 61056
rect 46768 61016 47072 61044
rect 47907 61016 47952 61044
rect 47946 61004 47952 61016
rect 48004 61004 48010 61056
rect 48682 61044 48688 61056
rect 48643 61016 48688 61044
rect 48682 61004 48688 61016
rect 48740 61004 48746 61056
rect 51166 61044 51172 61056
rect 51127 61016 51172 61044
rect 51166 61004 51172 61016
rect 51224 61004 51230 61056
rect 52086 61044 52092 61056
rect 52047 61016 52092 61044
rect 52086 61004 52092 61016
rect 52144 61004 52150 61056
rect 56870 61004 56876 61056
rect 56928 61044 56934 61056
rect 57241 61047 57299 61053
rect 57241 61044 57253 61047
rect 56928 61016 57253 61044
rect 56928 61004 56934 61016
rect 57241 61013 57253 61016
rect 57287 61013 57299 61047
rect 57241 61007 57299 61013
rect 58158 61004 58164 61056
rect 58216 61044 58222 61056
rect 58253 61047 58311 61053
rect 58253 61044 58265 61047
rect 58216 61016 58265 61044
rect 58216 61004 58222 61016
rect 58253 61013 58265 61016
rect 58299 61013 58311 61047
rect 58253 61007 58311 61013
rect 1104 60954 58880 60976
rect 1104 60902 19574 60954
rect 19626 60902 19638 60954
rect 19690 60902 19702 60954
rect 19754 60902 19766 60954
rect 19818 60902 19830 60954
rect 19882 60902 50294 60954
rect 50346 60902 50358 60954
rect 50410 60902 50422 60954
rect 50474 60902 50486 60954
rect 50538 60902 50550 60954
rect 50602 60902 58880 60954
rect 1104 60880 58880 60902
rect 5902 60800 5908 60852
rect 5960 60840 5966 60852
rect 23474 60840 23480 60852
rect 5960 60812 23480 60840
rect 5960 60800 5966 60812
rect 23474 60800 23480 60812
rect 23532 60800 23538 60852
rect 26878 60800 26884 60852
rect 26936 60840 26942 60852
rect 40954 60840 40960 60852
rect 26936 60812 40960 60840
rect 26936 60800 26942 60812
rect 40954 60800 40960 60812
rect 41012 60800 41018 60852
rect 58250 60840 58256 60852
rect 57164 60812 58256 60840
rect 1670 60772 1676 60784
rect 1631 60744 1676 60772
rect 1670 60732 1676 60744
rect 1728 60732 1734 60784
rect 3234 60772 3240 60784
rect 3195 60744 3240 60772
rect 3234 60732 3240 60744
rect 3292 60732 3298 60784
rect 3970 60772 3976 60784
rect 3931 60744 3976 60772
rect 3970 60732 3976 60744
rect 4028 60732 4034 60784
rect 8294 60732 8300 60784
rect 8352 60772 8358 60784
rect 8389 60775 8447 60781
rect 8389 60772 8401 60775
rect 8352 60744 8401 60772
rect 8352 60732 8358 60744
rect 8389 60741 8401 60744
rect 8435 60741 8447 60775
rect 9122 60772 9128 60784
rect 9083 60744 9128 60772
rect 8389 60735 8447 60741
rect 9122 60732 9128 60744
rect 9180 60732 9186 60784
rect 12066 60772 12072 60784
rect 12027 60744 12072 60772
rect 12066 60732 12072 60744
rect 12124 60732 12130 60784
rect 14826 60732 14832 60784
rect 14884 60772 14890 60784
rect 15013 60775 15071 60781
rect 15013 60772 15025 60775
rect 14884 60744 15025 60772
rect 14884 60732 14890 60744
rect 15013 60741 15025 60744
rect 15059 60741 15071 60775
rect 15013 60735 15071 60741
rect 19334 60732 19340 60784
rect 19392 60772 19398 60784
rect 19429 60775 19487 60781
rect 19429 60772 19441 60775
rect 19392 60744 19441 60772
rect 19392 60732 19398 60744
rect 19429 60741 19441 60744
rect 19475 60741 19487 60775
rect 24578 60772 24584 60784
rect 24539 60744 24584 60772
rect 19429 60735 19487 60741
rect 24578 60732 24584 60744
rect 24636 60732 24642 60784
rect 33962 60732 33968 60784
rect 34020 60772 34026 60784
rect 34149 60775 34207 60781
rect 34149 60772 34161 60775
rect 34020 60744 34161 60772
rect 34020 60732 34026 60744
rect 34149 60741 34161 60744
rect 34195 60741 34207 60775
rect 36354 60772 36360 60784
rect 36315 60744 36360 60772
rect 34149 60735 34207 60741
rect 36354 60732 36360 60744
rect 36412 60732 36418 60784
rect 46658 60772 46664 60784
rect 46619 60744 46664 60772
rect 46658 60732 46664 60744
rect 46716 60732 46722 60784
rect 50154 60732 50160 60784
rect 50212 60772 50218 60784
rect 50341 60775 50399 60781
rect 50341 60772 50353 60775
rect 50212 60744 50353 60772
rect 50212 60732 50218 60744
rect 50341 60741 50353 60744
rect 50387 60741 50399 60775
rect 50341 60735 50399 60741
rect 52454 60732 52460 60784
rect 52512 60772 52518 60784
rect 53009 60775 53067 60781
rect 53009 60772 53021 60775
rect 52512 60744 53021 60772
rect 52512 60732 52518 60744
rect 53009 60741 53021 60744
rect 53055 60741 53067 60775
rect 54754 60772 54760 60784
rect 54715 60744 54760 60772
rect 53009 60735 53067 60741
rect 54754 60732 54760 60744
rect 54812 60732 54818 60784
rect 55490 60772 55496 60784
rect 55451 60744 55496 60772
rect 55490 60732 55496 60744
rect 55548 60732 55554 60784
rect 57164 60781 57192 60812
rect 58250 60800 58256 60812
rect 58308 60800 58314 60852
rect 57149 60775 57207 60781
rect 57149 60741 57161 60775
rect 57195 60741 57207 60775
rect 57149 60735 57207 60741
rect 57790 60732 57796 60784
rect 57848 60772 57854 60784
rect 58161 60775 58219 60781
rect 58161 60772 58173 60775
rect 57848 60744 58173 60772
rect 57848 60732 57854 60744
rect 58161 60741 58173 60744
rect 58207 60741 58219 60775
rect 58161 60735 58219 60741
rect 26602 60664 26608 60716
rect 26660 60704 26666 60716
rect 27157 60707 27215 60713
rect 27157 60704 27169 60707
rect 26660 60676 27169 60704
rect 26660 60664 26666 60676
rect 27157 60673 27169 60676
rect 27203 60673 27215 60707
rect 29638 60704 29644 60716
rect 29599 60676 29644 60704
rect 27157 60667 27215 60673
rect 29638 60664 29644 60676
rect 29696 60664 29702 60716
rect 30282 60664 30288 60716
rect 30340 60704 30346 60716
rect 30377 60707 30435 60713
rect 30377 60704 30389 60707
rect 30340 60676 30389 60704
rect 30340 60664 30346 60676
rect 30377 60673 30389 60676
rect 30423 60673 30435 60707
rect 30377 60667 30435 60673
rect 41322 60664 41328 60716
rect 41380 60704 41386 60716
rect 41417 60707 41475 60713
rect 41417 60704 41429 60707
rect 41380 60676 41429 60704
rect 41380 60664 41386 60676
rect 41417 60673 41429 60676
rect 41463 60673 41475 60707
rect 49510 60704 49516 60716
rect 49471 60676 49516 60704
rect 41417 60667 41475 60673
rect 49510 60664 49516 60676
rect 49568 60664 49574 60716
rect 56134 60704 56140 60716
rect 56095 60676 56140 60704
rect 56134 60664 56140 60676
rect 56192 60664 56198 60716
rect 9309 60639 9367 60645
rect 9309 60605 9321 60639
rect 9355 60636 9367 60639
rect 15102 60636 15108 60648
rect 9355 60608 15108 60636
rect 9355 60605 9367 60608
rect 9309 60599 9367 60605
rect 15102 60596 15108 60608
rect 15160 60596 15166 60648
rect 56318 60636 56324 60648
rect 56279 60608 56324 60636
rect 56318 60596 56324 60608
rect 56376 60596 56382 60648
rect 4157 60571 4215 60577
rect 4157 60537 4169 60571
rect 4203 60568 4215 60571
rect 4798 60568 4804 60580
rect 4203 60540 4804 60568
rect 4203 60537 4215 60540
rect 4157 60531 4215 60537
rect 4798 60528 4804 60540
rect 4856 60528 4862 60580
rect 8570 60568 8576 60580
rect 8531 60540 8576 60568
rect 8570 60528 8576 60540
rect 8628 60528 8634 60580
rect 15197 60571 15255 60577
rect 15197 60537 15209 60571
rect 15243 60568 15255 60571
rect 16022 60568 16028 60580
rect 15243 60540 16028 60568
rect 15243 60537 15255 60540
rect 15197 60531 15255 60537
rect 16022 60528 16028 60540
rect 16080 60528 16086 60580
rect 19613 60571 19671 60577
rect 19613 60537 19625 60571
rect 19659 60568 19671 60571
rect 20438 60568 20444 60580
rect 19659 60540 20444 60568
rect 19659 60537 19671 60540
rect 19613 60531 19671 60537
rect 20438 60528 20444 60540
rect 20496 60528 20502 60580
rect 24765 60571 24823 60577
rect 24765 60537 24777 60571
rect 24811 60568 24823 60571
rect 25314 60568 25320 60580
rect 24811 60540 25320 60568
rect 24811 60537 24823 60540
rect 24765 60531 24823 60537
rect 25314 60528 25320 60540
rect 25372 60528 25378 60580
rect 1946 60500 1952 60512
rect 1907 60472 1952 60500
rect 1946 60460 1952 60472
rect 2004 60460 2010 60512
rect 3326 60500 3332 60512
rect 3287 60472 3332 60500
rect 3326 60460 3332 60472
rect 3384 60460 3390 60512
rect 12158 60500 12164 60512
rect 12119 60472 12164 60500
rect 12158 60460 12164 60472
rect 12216 60460 12222 60512
rect 27338 60500 27344 60512
rect 27299 60472 27344 60500
rect 27338 60460 27344 60472
rect 27396 60460 27402 60512
rect 29822 60500 29828 60512
rect 29783 60472 29828 60500
rect 29822 60460 29828 60472
rect 29880 60460 29886 60512
rect 30558 60500 30564 60512
rect 30519 60472 30564 60500
rect 30558 60460 30564 60472
rect 30616 60460 30622 60512
rect 34238 60500 34244 60512
rect 34199 60472 34244 60500
rect 34238 60460 34244 60472
rect 34296 60460 34302 60512
rect 36446 60500 36452 60512
rect 36407 60472 36452 60500
rect 36446 60460 36452 60472
rect 36504 60460 36510 60512
rect 41598 60500 41604 60512
rect 41559 60472 41604 60500
rect 41598 60460 41604 60472
rect 41656 60460 41662 60512
rect 46750 60500 46756 60512
rect 46711 60472 46756 60500
rect 46750 60460 46756 60472
rect 46808 60460 46814 60512
rect 49694 60500 49700 60512
rect 49655 60472 49700 60500
rect 49694 60460 49700 60472
rect 49752 60460 49758 60512
rect 49786 60460 49792 60512
rect 49844 60500 49850 60512
rect 50433 60503 50491 60509
rect 50433 60500 50445 60503
rect 49844 60472 50445 60500
rect 49844 60460 49850 60472
rect 50433 60469 50445 60472
rect 50479 60469 50491 60503
rect 53098 60500 53104 60512
rect 53059 60472 53104 60500
rect 50433 60463 50491 60469
rect 53098 60460 53104 60472
rect 53156 60460 53162 60512
rect 54846 60500 54852 60512
rect 54807 60472 54852 60500
rect 54846 60460 54852 60472
rect 54904 60460 54910 60512
rect 55582 60500 55588 60512
rect 55543 60472 55588 60500
rect 55582 60460 55588 60472
rect 55640 60460 55646 60512
rect 57054 60460 57060 60512
rect 57112 60500 57118 60512
rect 57241 60503 57299 60509
rect 57241 60500 57253 60503
rect 57112 60472 57253 60500
rect 57112 60460 57118 60472
rect 57241 60469 57253 60472
rect 57287 60469 57299 60503
rect 58250 60500 58256 60512
rect 58211 60472 58256 60500
rect 57241 60463 57299 60469
rect 58250 60460 58256 60472
rect 58308 60460 58314 60512
rect 1104 60410 58880 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 58880 60410
rect 1104 60336 58880 60358
rect 12158 60256 12164 60308
rect 12216 60296 12222 60308
rect 21818 60296 21824 60308
rect 12216 60268 21824 60296
rect 12216 60256 12222 60268
rect 21818 60256 21824 60268
rect 21876 60256 21882 60308
rect 28258 60256 28264 60308
rect 28316 60296 28322 60308
rect 41598 60296 41604 60308
rect 28316 60268 41604 60296
rect 28316 60256 28322 60268
rect 41598 60256 41604 60268
rect 41656 60256 41662 60308
rect 49602 60256 49608 60308
rect 49660 60296 49666 60308
rect 58250 60296 58256 60308
rect 49660 60268 58256 60296
rect 49660 60256 49666 60268
rect 58250 60256 58256 60268
rect 58308 60256 58314 60308
rect 54478 60188 54484 60240
rect 54536 60228 54542 60240
rect 57241 60231 57299 60237
rect 57241 60228 57253 60231
rect 54536 60200 57253 60228
rect 54536 60188 54542 60200
rect 57241 60197 57253 60200
rect 57287 60197 57299 60231
rect 57241 60191 57299 60197
rect 1578 60052 1584 60104
rect 1636 60092 1642 60104
rect 1765 60095 1823 60101
rect 1765 60092 1777 60095
rect 1636 60064 1777 60092
rect 1636 60052 1642 60064
rect 1765 60061 1777 60064
rect 1811 60061 1823 60095
rect 2498 60092 2504 60104
rect 2459 60064 2504 60092
rect 1765 60055 1823 60061
rect 2498 60052 2504 60064
rect 2556 60052 2562 60104
rect 56226 60092 56232 60104
rect 56187 60064 56232 60092
rect 56226 60052 56232 60064
rect 56284 60052 56290 60104
rect 1949 60027 2007 60033
rect 1949 59993 1961 60027
rect 1995 60024 2007 60027
rect 2038 60024 2044 60036
rect 1995 59996 2044 60024
rect 1995 59993 2007 59996
rect 1949 59987 2007 59993
rect 2038 59984 2044 59996
rect 2096 59984 2102 60036
rect 56042 59984 56048 60036
rect 56100 60024 56106 60036
rect 57057 60027 57115 60033
rect 57057 60024 57069 60027
rect 56100 59996 57069 60024
rect 56100 59984 56106 59996
rect 57057 59993 57069 59996
rect 57103 59993 57115 60027
rect 57974 60024 57980 60036
rect 57935 59996 57980 60024
rect 57057 59987 57115 59993
rect 57974 59984 57980 59996
rect 58032 59984 58038 60036
rect 58345 60027 58403 60033
rect 58345 59993 58357 60027
rect 58391 60024 58403 60027
rect 58986 60024 58992 60036
rect 58391 59996 58992 60024
rect 58391 59993 58403 59996
rect 58345 59987 58403 59993
rect 58986 59984 58992 59996
rect 59044 59984 59050 60036
rect 2406 59916 2412 59968
rect 2464 59956 2470 59968
rect 2593 59959 2651 59965
rect 2593 59956 2605 59959
rect 2464 59928 2605 59956
rect 2464 59916 2470 59928
rect 2593 59925 2605 59928
rect 2639 59925 2651 59959
rect 2593 59919 2651 59925
rect 54754 59916 54760 59968
rect 54812 59956 54818 59968
rect 56321 59959 56379 59965
rect 56321 59956 56333 59959
rect 54812 59928 56333 59956
rect 54812 59916 54818 59928
rect 56321 59925 56333 59928
rect 56367 59925 56379 59959
rect 56321 59919 56379 59925
rect 1104 59866 58880 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 58880 59866
rect 1104 59792 58880 59814
rect 842 59644 848 59696
rect 900 59684 906 59696
rect 2409 59687 2467 59693
rect 2409 59684 2421 59687
rect 900 59656 2421 59684
rect 900 59644 906 59656
rect 2409 59653 2421 59656
rect 2455 59653 2467 59687
rect 58710 59684 58716 59696
rect 2409 59647 2467 59653
rect 57072 59656 58716 59684
rect 1578 59616 1584 59628
rect 1539 59588 1584 59616
rect 1578 59576 1584 59588
rect 1636 59576 1642 59628
rect 57072 59625 57100 59656
rect 58710 59644 58716 59656
rect 58768 59644 58774 59696
rect 57057 59619 57115 59625
rect 57057 59585 57069 59619
rect 57103 59585 57115 59619
rect 57057 59579 57115 59585
rect 57882 59576 57888 59628
rect 57940 59616 57946 59628
rect 58069 59619 58127 59625
rect 58069 59616 58081 59619
rect 57940 59588 58081 59616
rect 57940 59576 57946 59588
rect 58069 59585 58081 59588
rect 58115 59585 58127 59619
rect 58069 59579 58127 59585
rect 57238 59548 57244 59560
rect 57199 59520 57244 59548
rect 57238 59508 57244 59520
rect 57296 59508 57302 59560
rect 2590 59480 2596 59492
rect 2551 59452 2596 59480
rect 2590 59440 2596 59452
rect 2648 59440 2654 59492
rect 1765 59415 1823 59421
rect 1765 59381 1777 59415
rect 1811 59412 1823 59415
rect 2682 59412 2688 59424
rect 1811 59384 2688 59412
rect 1811 59381 1823 59384
rect 1765 59375 1823 59381
rect 2682 59372 2688 59384
rect 2740 59372 2746 59424
rect 31662 59372 31668 59424
rect 31720 59412 31726 59424
rect 33686 59412 33692 59424
rect 31720 59384 33692 59412
rect 31720 59372 31726 59384
rect 33686 59372 33692 59384
rect 33744 59372 33750 59424
rect 58253 59415 58311 59421
rect 58253 59381 58265 59415
rect 58299 59412 58311 59415
rect 59170 59412 59176 59424
rect 58299 59384 59176 59412
rect 58299 59381 58311 59384
rect 58253 59375 58311 59381
rect 59170 59372 59176 59384
rect 59228 59372 59234 59424
rect 1104 59322 58880 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 58880 59322
rect 1104 59248 58880 59270
rect 1946 59032 1952 59084
rect 2004 59072 2010 59084
rect 43901 59075 43959 59081
rect 43901 59072 43913 59075
rect 2004 59044 43913 59072
rect 2004 59032 2010 59044
rect 43901 59041 43913 59044
rect 43947 59041 43959 59075
rect 44361 59075 44419 59081
rect 44361 59072 44373 59075
rect 43901 59035 43959 59041
rect 44008 59044 44373 59072
rect 1578 59004 1584 59016
rect 1539 58976 1584 59004
rect 1578 58964 1584 58976
rect 1636 58964 1642 59016
rect 40126 58964 40132 59016
rect 40184 59004 40190 59016
rect 44008 59004 44036 59044
rect 44361 59041 44373 59044
rect 44407 59041 44419 59075
rect 53098 59072 53104 59084
rect 44361 59035 44419 59041
rect 44468 59044 53104 59072
rect 40184 58976 44036 59004
rect 40184 58964 40190 58976
rect 44082 58964 44088 59016
rect 44140 59004 44146 59016
rect 44468 59013 44496 59044
rect 53098 59032 53104 59044
rect 53156 59032 53162 59084
rect 44453 59007 44511 59013
rect 44140 58976 44185 59004
rect 44140 58964 44146 58976
rect 44453 58973 44465 59007
rect 44499 58973 44511 59007
rect 44453 58967 44511 58973
rect 57241 59007 57299 59013
rect 57241 58973 57253 59007
rect 57287 59004 57299 59007
rect 57330 59004 57336 59016
rect 57287 58976 57336 59004
rect 57287 58973 57299 58976
rect 57241 58967 57299 58973
rect 57330 58964 57336 58976
rect 57388 58964 57394 59016
rect 56502 58896 56508 58948
rect 56560 58936 56566 58948
rect 57977 58939 58035 58945
rect 57977 58936 57989 58939
rect 56560 58908 57989 58936
rect 56560 58896 56566 58908
rect 57977 58905 57989 58908
rect 58023 58905 58035 58939
rect 57977 58899 58035 58905
rect 1762 58868 1768 58880
rect 1723 58840 1768 58868
rect 1762 58828 1768 58840
rect 1820 58828 1826 58880
rect 43717 58871 43775 58877
rect 43717 58837 43729 58871
rect 43763 58868 43775 58871
rect 44818 58868 44824 58880
rect 43763 58840 44824 58868
rect 43763 58837 43775 58840
rect 43717 58831 43775 58837
rect 44818 58828 44824 58840
rect 44876 58828 44882 58880
rect 57330 58868 57336 58880
rect 57291 58840 57336 58868
rect 57330 58828 57336 58840
rect 57388 58828 57394 58880
rect 58066 58868 58072 58880
rect 58027 58840 58072 58868
rect 58066 58828 58072 58840
rect 58124 58828 58130 58880
rect 1104 58778 58880 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 58880 58778
rect 1104 58704 58880 58726
rect 23106 58664 23112 58676
rect 14936 58636 23112 58664
rect 1670 58528 1676 58540
rect 1631 58500 1676 58528
rect 1670 58488 1676 58500
rect 1728 58488 1734 58540
rect 14829 58531 14887 58537
rect 14829 58497 14841 58531
rect 14875 58497 14887 58531
rect 14936 58528 14964 58636
rect 23106 58624 23112 58636
rect 23164 58624 23170 58676
rect 58158 58664 58164 58676
rect 45526 58636 58164 58664
rect 15102 58596 15108 58608
rect 15063 58568 15108 58596
rect 15102 58556 15108 58568
rect 15160 58556 15166 58608
rect 16666 58556 16672 58608
rect 16724 58596 16730 58608
rect 17129 58599 17187 58605
rect 17129 58596 17141 58599
rect 16724 58568 17141 58596
rect 16724 58556 16730 58568
rect 17129 58565 17141 58568
rect 17175 58565 17187 58599
rect 17129 58559 17187 58565
rect 17218 58556 17224 58608
rect 17276 58596 17282 58608
rect 45526 58596 45554 58636
rect 58158 58624 58164 58636
rect 58216 58624 58222 58676
rect 17276 58568 17321 58596
rect 22066 58568 45554 58596
rect 17276 58556 17282 58568
rect 15013 58531 15071 58537
rect 15013 58528 15025 58531
rect 14936 58500 15025 58528
rect 14829 58491 14887 58497
rect 15013 58497 15025 58500
rect 15059 58497 15071 58531
rect 15013 58491 15071 58497
rect 15249 58531 15307 58537
rect 15249 58497 15261 58531
rect 15295 58528 15307 58531
rect 16758 58528 16764 58540
rect 15295 58500 16764 58528
rect 15295 58497 15307 58500
rect 15249 58491 15307 58497
rect 14553 58463 14611 58469
rect 14553 58429 14565 58463
rect 14599 58460 14611 58463
rect 14844 58460 14872 58491
rect 16758 58488 16764 58500
rect 16816 58488 16822 58540
rect 17402 58537 17408 58540
rect 16945 58531 17003 58537
rect 16945 58497 16957 58531
rect 16991 58497 17003 58531
rect 16945 58491 17003 58497
rect 17365 58531 17408 58537
rect 17365 58497 17377 58531
rect 17460 58528 17466 58540
rect 21910 58528 21916 58540
rect 17460 58500 21916 58528
rect 17365 58491 17408 58497
rect 16850 58460 16856 58472
rect 14599 58432 16856 58460
rect 14599 58429 14611 58432
rect 14553 58423 14611 58429
rect 16850 58420 16856 58432
rect 16908 58420 16914 58472
rect 16960 58460 16988 58491
rect 17402 58488 17408 58491
rect 17460 58488 17466 58500
rect 21910 58488 21916 58500
rect 21968 58488 21974 58540
rect 16960 58432 17080 58460
rect 1949 58395 2007 58401
rect 1949 58361 1961 58395
rect 1995 58392 2007 58395
rect 1995 58364 15516 58392
rect 1995 58361 2007 58364
rect 1949 58355 2007 58361
rect 15378 58324 15384 58336
rect 15339 58296 15384 58324
rect 15378 58284 15384 58296
rect 15436 58284 15442 58336
rect 15488 58324 15516 58364
rect 16574 58352 16580 58404
rect 16632 58392 16638 58404
rect 17052 58392 17080 58432
rect 17218 58420 17224 58472
rect 17276 58460 17282 58472
rect 22066 58460 22094 58568
rect 39485 58531 39543 58537
rect 39485 58497 39497 58531
rect 39531 58497 39543 58531
rect 39666 58528 39672 58540
rect 39627 58500 39672 58528
rect 39485 58491 39543 58497
rect 17276 58432 22094 58460
rect 39500 58460 39528 58491
rect 39666 58488 39672 58500
rect 39724 58488 39730 58540
rect 39758 58488 39764 58540
rect 39816 58528 39822 58540
rect 39905 58531 39963 58537
rect 39816 58500 39861 58528
rect 39816 58488 39822 58500
rect 39905 58497 39917 58531
rect 39951 58528 39963 58531
rect 43990 58528 43996 58540
rect 39951 58500 43996 58528
rect 39951 58497 39963 58500
rect 39905 58491 39963 58497
rect 43990 58488 43996 58500
rect 44048 58488 44054 58540
rect 58158 58528 58164 58540
rect 58119 58500 58164 58528
rect 58158 58488 58164 58500
rect 58216 58488 58222 58540
rect 57330 58460 57336 58472
rect 39500 58432 57336 58460
rect 17276 58420 17282 58432
rect 57330 58420 57336 58432
rect 57388 58420 57394 58472
rect 43898 58392 43904 58404
rect 16632 58364 17080 58392
rect 17236 58364 43904 58392
rect 16632 58352 16638 58364
rect 17236 58324 17264 58364
rect 43898 58352 43904 58364
rect 43956 58352 43962 58404
rect 17494 58324 17500 58336
rect 15488 58296 17264 58324
rect 17455 58296 17500 58324
rect 17494 58284 17500 58296
rect 17552 58284 17558 58336
rect 40034 58324 40040 58336
rect 39995 58296 40040 58324
rect 40034 58284 40040 58296
rect 40092 58284 40098 58336
rect 55214 58284 55220 58336
rect 55272 58324 55278 58336
rect 58253 58327 58311 58333
rect 58253 58324 58265 58327
rect 55272 58296 58265 58324
rect 55272 58284 55278 58296
rect 58253 58293 58265 58296
rect 58299 58293 58311 58327
rect 58253 58287 58311 58293
rect 1104 58234 58880 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 58880 58234
rect 1104 58160 58880 58182
rect 16666 58080 16672 58132
rect 16724 58120 16730 58132
rect 17126 58120 17132 58132
rect 16724 58092 17132 58120
rect 16724 58080 16730 58092
rect 17126 58080 17132 58092
rect 17184 58080 17190 58132
rect 23124 58024 25084 58052
rect 1578 57916 1584 57928
rect 1539 57888 1584 57916
rect 1578 57876 1584 57888
rect 1636 57876 1642 57928
rect 21266 57916 21272 57928
rect 21227 57888 21272 57916
rect 21266 57876 21272 57888
rect 21324 57876 21330 57928
rect 21358 57876 21364 57928
rect 21416 57916 21422 57928
rect 21634 57916 21640 57928
rect 21416 57888 21461 57916
rect 21595 57888 21640 57916
rect 21416 57876 21422 57888
rect 21634 57876 21640 57888
rect 21692 57876 21698 57928
rect 21913 57919 21971 57925
rect 21913 57885 21925 57919
rect 21959 57916 21971 57919
rect 22002 57916 22008 57928
rect 21959 57888 22008 57916
rect 21959 57885 21971 57888
rect 21913 57879 21971 57885
rect 22002 57876 22008 57888
rect 22060 57876 22066 57928
rect 22097 57919 22155 57925
rect 22097 57885 22109 57919
rect 22143 57885 22155 57919
rect 22097 57879 22155 57885
rect 18138 57808 18144 57860
rect 18196 57848 18202 57860
rect 18196 57820 21036 57848
rect 18196 57808 18202 57820
rect 1765 57783 1823 57789
rect 1765 57749 1777 57783
rect 1811 57780 1823 57783
rect 1946 57780 1952 57792
rect 1811 57752 1952 57780
rect 1811 57749 1823 57752
rect 1765 57743 1823 57749
rect 1946 57740 1952 57752
rect 2004 57740 2010 57792
rect 20898 57780 20904 57792
rect 20859 57752 20904 57780
rect 20898 57740 20904 57752
rect 20956 57740 20962 57792
rect 21008 57780 21036 57820
rect 21818 57808 21824 57860
rect 21876 57848 21882 57860
rect 22112 57848 22140 57879
rect 22462 57876 22468 57928
rect 22520 57916 22526 57928
rect 22741 57919 22799 57925
rect 22741 57916 22753 57919
rect 22520 57888 22753 57916
rect 22520 57876 22526 57888
rect 22741 57885 22753 57888
rect 22787 57885 22799 57919
rect 22741 57879 22799 57885
rect 22834 57919 22892 57925
rect 22834 57885 22846 57919
rect 22880 57885 22892 57919
rect 22834 57879 22892 57885
rect 21876 57820 22140 57848
rect 21876 57808 21882 57820
rect 22848 57780 22876 57879
rect 23014 57876 23020 57928
rect 23072 57916 23078 57928
rect 23124 57916 23152 58024
rect 23400 57956 24716 57984
rect 23072 57888 23165 57916
rect 23072 57876 23078 57888
rect 23198 57876 23204 57928
rect 23256 57925 23262 57928
rect 23256 57916 23264 57925
rect 23400 57916 23428 57956
rect 23256 57888 23428 57916
rect 23256 57879 23264 57888
rect 23256 57876 23262 57879
rect 23474 57876 23480 57928
rect 23532 57916 23538 57928
rect 24581 57919 24639 57925
rect 24581 57916 24593 57919
rect 23532 57888 24593 57916
rect 23532 57876 23538 57888
rect 24581 57885 24593 57888
rect 24627 57885 24639 57919
rect 24688 57916 24716 57956
rect 24954 57919 25012 57925
rect 24954 57916 24966 57919
rect 24688 57888 24966 57916
rect 24581 57879 24639 57885
rect 24954 57885 24966 57888
rect 25000 57885 25012 57919
rect 25056 57916 25084 58024
rect 31864 58024 32996 58052
rect 31864 57984 31892 58024
rect 31680 57956 31892 57984
rect 32508 57956 32904 57984
rect 30742 57916 30748 57928
rect 25056 57888 30748 57916
rect 24954 57879 25012 57885
rect 30742 57876 30748 57888
rect 30800 57876 30806 57928
rect 31680 57916 31708 57956
rect 32508 57928 32536 57956
rect 31846 57916 31852 57928
rect 30944 57888 31708 57916
rect 31807 57888 31852 57916
rect 23109 57851 23167 57857
rect 23109 57817 23121 57851
rect 23155 57848 23167 57851
rect 24762 57848 24768 57860
rect 23155 57820 24624 57848
rect 24723 57820 24768 57848
rect 23155 57817 23167 57820
rect 23109 57811 23167 57817
rect 23382 57780 23388 57792
rect 21008 57752 22876 57780
rect 23343 57752 23388 57780
rect 23382 57740 23388 57752
rect 23440 57740 23446 57792
rect 24596 57780 24624 57820
rect 24762 57808 24768 57820
rect 24820 57808 24826 57860
rect 24854 57808 24860 57860
rect 24912 57848 24918 57860
rect 30944 57848 30972 57888
rect 31846 57876 31852 57888
rect 31904 57876 31910 57928
rect 31938 57876 31944 57928
rect 31996 57916 32002 57928
rect 32214 57916 32220 57928
rect 31996 57888 32041 57916
rect 32175 57888 32220 57916
rect 31996 57876 32002 57888
rect 32214 57876 32220 57888
rect 32272 57876 32278 57928
rect 32490 57916 32496 57928
rect 32451 57888 32496 57916
rect 32490 57876 32496 57888
rect 32548 57876 32554 57928
rect 32674 57916 32680 57928
rect 32635 57888 32680 57916
rect 32674 57876 32680 57888
rect 32732 57876 32738 57928
rect 32876 57848 32904 57956
rect 32968 57916 32996 58024
rect 43898 57984 43904 57996
rect 38304 57956 40356 57984
rect 43859 57956 43904 57984
rect 37274 57916 37280 57928
rect 32968 57888 37280 57916
rect 37274 57876 37280 57888
rect 37332 57876 37338 57928
rect 38304 57848 38332 57956
rect 38654 57916 38660 57928
rect 38615 57888 38660 57916
rect 38654 57876 38660 57888
rect 38712 57876 38718 57928
rect 40218 57916 40224 57928
rect 38764 57888 40224 57916
rect 38470 57848 38476 57860
rect 24912 57820 24957 57848
rect 25056 57820 30972 57848
rect 31036 57820 31616 57848
rect 32876 57820 38332 57848
rect 38431 57820 38476 57848
rect 24912 57808 24918 57820
rect 25056 57780 25084 57820
rect 24596 57752 25084 57780
rect 25150 57783 25208 57789
rect 25150 57749 25162 57783
rect 25196 57780 25208 57783
rect 25406 57780 25412 57792
rect 25196 57752 25412 57780
rect 25196 57749 25208 57752
rect 25150 57743 25208 57749
rect 25406 57740 25412 57752
rect 25464 57740 25470 57792
rect 25498 57740 25504 57792
rect 25556 57780 25562 57792
rect 31036 57780 31064 57820
rect 31478 57780 31484 57792
rect 25556 57752 31064 57780
rect 31439 57752 31484 57780
rect 25556 57740 25562 57752
rect 31478 57740 31484 57752
rect 31536 57740 31542 57792
rect 31588 57780 31616 57820
rect 38470 57808 38476 57820
rect 38528 57808 38534 57860
rect 38764 57848 38792 57888
rect 40218 57876 40224 57888
rect 40276 57876 40282 57928
rect 40328 57916 40356 57956
rect 43898 57944 43904 57956
rect 43956 57944 43962 57996
rect 43990 57944 43996 57996
rect 44048 57984 44054 57996
rect 44361 57987 44419 57993
rect 44361 57984 44373 57987
rect 44048 57956 44373 57984
rect 44048 57944 44054 57956
rect 44361 57953 44373 57956
rect 44407 57953 44419 57987
rect 44361 57947 44419 57953
rect 54404 57956 54708 57984
rect 43806 57916 43812 57928
rect 40328 57888 43812 57916
rect 43806 57876 43812 57888
rect 43864 57916 43870 57928
rect 44082 57916 44088 57928
rect 43864 57888 44088 57916
rect 43864 57876 43870 57888
rect 44082 57876 44088 57888
rect 44140 57876 44146 57928
rect 44453 57919 44511 57925
rect 44453 57885 44465 57919
rect 44499 57885 44511 57919
rect 44453 57879 44511 57885
rect 38930 57848 38936 57860
rect 38580 57820 38792 57848
rect 38891 57820 38936 57848
rect 38580 57780 38608 57820
rect 38930 57808 38936 57820
rect 38988 57848 38994 57860
rect 39666 57848 39672 57860
rect 38988 57820 39672 57848
rect 38988 57808 38994 57820
rect 39666 57808 39672 57820
rect 39724 57808 39730 57860
rect 44468 57848 44496 57879
rect 50062 57876 50068 57928
rect 50120 57916 50126 57928
rect 54113 57919 54171 57925
rect 50120 57888 51074 57916
rect 50120 57876 50126 57888
rect 49786 57848 49792 57860
rect 44468 57820 49792 57848
rect 49786 57808 49792 57820
rect 49844 57808 49850 57860
rect 38838 57780 38844 57792
rect 31588 57752 38608 57780
rect 38799 57752 38844 57780
rect 38838 57740 38844 57752
rect 38896 57740 38902 57792
rect 43717 57783 43775 57789
rect 43717 57749 43729 57783
rect 43763 57780 43775 57783
rect 44082 57780 44088 57792
rect 43763 57752 44088 57780
rect 43763 57749 43775 57752
rect 43717 57743 43775 57749
rect 44082 57740 44088 57752
rect 44140 57740 44146 57792
rect 51046 57780 51074 57888
rect 54113 57885 54125 57919
rect 54159 57916 54171 57919
rect 54404 57916 54432 57956
rect 54570 57925 54576 57928
rect 54159 57888 54432 57916
rect 54533 57919 54576 57925
rect 54159 57885 54171 57888
rect 54113 57879 54171 57885
rect 54533 57885 54545 57919
rect 54533 57879 54576 57885
rect 54570 57876 54576 57879
rect 54628 57876 54634 57928
rect 54680 57916 54708 57956
rect 55214 57916 55220 57928
rect 54680 57888 55220 57916
rect 55214 57876 55220 57888
rect 55272 57876 55278 57928
rect 54018 57808 54024 57860
rect 54076 57848 54082 57860
rect 54297 57851 54355 57857
rect 54297 57848 54309 57851
rect 54076 57820 54309 57848
rect 54076 57808 54082 57820
rect 54297 57817 54309 57820
rect 54343 57817 54355 57851
rect 54297 57811 54355 57817
rect 54389 57851 54447 57857
rect 54389 57817 54401 57851
rect 54435 57848 54447 57851
rect 54754 57848 54760 57860
rect 54435 57820 54760 57848
rect 54435 57817 54447 57820
rect 54389 57811 54447 57817
rect 54754 57808 54760 57820
rect 54812 57808 54818 57860
rect 58158 57848 58164 57860
rect 58119 57820 58164 57848
rect 58158 57808 58164 57820
rect 58216 57808 58222 57860
rect 54673 57783 54731 57789
rect 54673 57780 54685 57783
rect 51046 57752 54685 57780
rect 54673 57749 54685 57752
rect 54719 57749 54731 57783
rect 58250 57780 58256 57792
rect 58211 57752 58256 57780
rect 54673 57743 54731 57749
rect 58250 57740 58256 57752
rect 58308 57740 58314 57792
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 20717 57579 20775 57585
rect 20717 57545 20729 57579
rect 20763 57576 20775 57579
rect 21634 57576 21640 57588
rect 20763 57548 21640 57576
rect 20763 57545 20775 57548
rect 20717 57539 20775 57545
rect 21634 57536 21640 57548
rect 21692 57536 21698 57588
rect 25498 57576 25504 57588
rect 21744 57548 25504 57576
rect 20438 57508 20444 57520
rect 20399 57480 20444 57508
rect 20438 57468 20444 57480
rect 20496 57468 20502 57520
rect 21358 57468 21364 57520
rect 21416 57508 21422 57520
rect 21744 57508 21772 57548
rect 25498 57536 25504 57548
rect 25556 57536 25562 57588
rect 34514 57576 34520 57588
rect 25608 57548 34520 57576
rect 21416 57480 21772 57508
rect 21416 57468 21422 57480
rect 21818 57468 21824 57520
rect 21876 57508 21882 57520
rect 23382 57508 23388 57520
rect 21876 57480 23388 57508
rect 21876 57468 21882 57480
rect 23382 57468 23388 57480
rect 23440 57468 23446 57520
rect 19889 57443 19947 57449
rect 19889 57409 19901 57443
rect 19935 57440 19947 57443
rect 20162 57440 20168 57452
rect 19935 57412 20168 57440
rect 19935 57409 19947 57412
rect 19889 57403 19947 57409
rect 20162 57400 20168 57412
rect 20220 57400 20226 57452
rect 20349 57443 20407 57449
rect 20349 57409 20361 57443
rect 20395 57409 20407 57443
rect 20349 57403 20407 57409
rect 20533 57443 20591 57449
rect 20533 57409 20545 57443
rect 20579 57440 20591 57443
rect 20622 57440 20628 57452
rect 20579 57412 20628 57440
rect 20579 57409 20591 57412
rect 20533 57403 20591 57409
rect 20364 57372 20392 57403
rect 20622 57400 20628 57412
rect 20680 57400 20686 57452
rect 21266 57400 21272 57452
rect 21324 57440 21330 57452
rect 22186 57440 22192 57452
rect 21324 57412 22192 57440
rect 21324 57400 21330 57412
rect 22186 57400 22192 57412
rect 22244 57400 22250 57452
rect 22462 57400 22468 57452
rect 22520 57440 22526 57452
rect 25608 57440 25636 57548
rect 34514 57536 34520 57548
rect 34572 57536 34578 57588
rect 38654 57576 38660 57588
rect 36004 57548 38516 57576
rect 38615 57548 38660 57576
rect 32214 57508 32220 57520
rect 31128 57480 32220 57508
rect 31128 57452 31156 57480
rect 32214 57468 32220 57480
rect 32272 57468 32278 57520
rect 29914 57440 29920 57452
rect 22520 57412 25636 57440
rect 25700 57412 29920 57440
rect 22520 57400 22526 57412
rect 22204 57372 22232 57400
rect 23198 57372 23204 57384
rect 20364 57344 21588 57372
rect 22204 57344 23204 57372
rect 21560 57316 21588 57344
rect 23198 57332 23204 57344
rect 23256 57372 23262 57384
rect 25700 57372 25728 57412
rect 29914 57400 29920 57412
rect 29972 57400 29978 57452
rect 30742 57440 30748 57452
rect 30703 57412 30748 57440
rect 30742 57400 30748 57412
rect 30800 57400 30806 57452
rect 31018 57440 31024 57452
rect 30979 57412 31024 57440
rect 31018 57400 31024 57412
rect 31076 57400 31082 57452
rect 31110 57400 31116 57452
rect 31168 57440 31174 57452
rect 31386 57440 31392 57452
rect 31168 57412 31213 57440
rect 31347 57412 31392 57440
rect 31168 57400 31174 57412
rect 31386 57400 31392 57412
rect 31444 57400 31450 57452
rect 31570 57440 31576 57452
rect 31531 57412 31576 57440
rect 31570 57400 31576 57412
rect 31628 57400 31634 57452
rect 36004 57449 36032 57548
rect 37734 57468 37740 57520
rect 37792 57508 37798 57520
rect 38381 57511 38439 57517
rect 38381 57508 38393 57511
rect 37792 57480 38393 57508
rect 37792 57468 37798 57480
rect 38381 57477 38393 57480
rect 38427 57477 38439 57511
rect 38488 57508 38516 57548
rect 38654 57536 38660 57548
rect 38712 57536 38718 57588
rect 38838 57536 38844 57588
rect 38896 57576 38902 57588
rect 49602 57576 49608 57588
rect 38896 57548 49608 57576
rect 38896 57536 38902 57548
rect 49602 57536 49608 57548
rect 49660 57536 49666 57588
rect 54570 57576 54576 57588
rect 53944 57548 54576 57576
rect 51074 57508 51080 57520
rect 38488 57480 51080 57508
rect 38381 57471 38439 57477
rect 51074 57468 51080 57480
rect 51132 57468 51138 57520
rect 35713 57443 35771 57449
rect 35713 57409 35725 57443
rect 35759 57440 35771 57443
rect 35989 57443 36047 57449
rect 35759 57412 35793 57440
rect 35759 57409 35771 57412
rect 35713 57403 35771 57409
rect 35989 57409 36001 57443
rect 36035 57409 36047 57443
rect 35989 57403 36047 57409
rect 23256 57344 25728 57372
rect 23256 57332 23262 57344
rect 25774 57332 25780 57384
rect 25832 57372 25838 57384
rect 35728 57372 35756 57403
rect 36078 57400 36084 57452
rect 36136 57440 36142 57452
rect 36354 57440 36360 57452
rect 36136 57412 36181 57440
rect 36315 57412 36360 57440
rect 36136 57400 36142 57412
rect 36354 57400 36360 57412
rect 36412 57400 36418 57452
rect 36630 57440 36636 57452
rect 36591 57412 36636 57440
rect 36630 57400 36636 57412
rect 36688 57400 36694 57452
rect 38102 57440 38108 57452
rect 38063 57412 38108 57440
rect 38102 57400 38108 57412
rect 38160 57400 38166 57452
rect 38194 57400 38200 57452
rect 38252 57440 38258 57452
rect 38289 57443 38347 57449
rect 38289 57440 38301 57443
rect 38252 57412 38301 57440
rect 38252 57400 38258 57412
rect 38289 57409 38301 57412
rect 38335 57409 38347 57443
rect 38289 57403 38347 57409
rect 38473 57443 38531 57449
rect 38473 57409 38485 57443
rect 38519 57440 38531 57443
rect 38562 57440 38568 57452
rect 38519 57412 38568 57440
rect 38519 57409 38531 57412
rect 38473 57403 38531 57409
rect 38562 57400 38568 57412
rect 38620 57440 38626 57452
rect 40126 57440 40132 57452
rect 38620 57412 40132 57440
rect 38620 57400 38626 57412
rect 40126 57400 40132 57412
rect 40184 57400 40190 57452
rect 53944 57440 53972 57548
rect 54570 57536 54576 57548
rect 54628 57576 54634 57588
rect 54628 57548 55076 57576
rect 54628 57536 54634 57548
rect 45526 57412 53972 57440
rect 45526 57372 45554 57412
rect 54018 57400 54024 57452
rect 54076 57440 54082 57452
rect 54433 57443 54491 57449
rect 54433 57440 54445 57443
rect 54076 57412 54445 57440
rect 54076 57400 54082 57412
rect 54433 57409 54445 57412
rect 54479 57409 54491 57443
rect 54846 57440 54852 57452
rect 54807 57412 54852 57440
rect 54433 57403 54491 57409
rect 54846 57400 54852 57412
rect 54904 57400 54910 57452
rect 55048 57449 55076 57548
rect 55033 57443 55091 57449
rect 55033 57409 55045 57443
rect 55079 57409 55091 57443
rect 58158 57440 58164 57452
rect 58119 57412 58164 57440
rect 55033 57403 55091 57409
rect 58158 57400 58164 57412
rect 58216 57400 58222 57452
rect 53926 57372 53932 57384
rect 25832 57344 38148 57372
rect 25832 57332 25838 57344
rect 21542 57264 21548 57316
rect 21600 57304 21606 57316
rect 38010 57304 38016 57316
rect 21600 57276 25912 57304
rect 21600 57264 21606 57276
rect 20622 57196 20628 57248
rect 20680 57236 20686 57248
rect 21910 57236 21916 57248
rect 20680 57208 21916 57236
rect 20680 57196 20686 57208
rect 21910 57196 21916 57208
rect 21968 57236 21974 57248
rect 23014 57236 23020 57248
rect 21968 57208 23020 57236
rect 21968 57196 21974 57208
rect 23014 57196 23020 57208
rect 23072 57196 23078 57248
rect 23106 57196 23112 57248
rect 23164 57236 23170 57248
rect 25590 57236 25596 57248
rect 23164 57208 25596 57236
rect 23164 57196 23170 57208
rect 25590 57196 25596 57208
rect 25648 57196 25654 57248
rect 25884 57236 25912 57276
rect 26206 57276 38016 57304
rect 26206 57236 26234 57276
rect 38010 57264 38016 57276
rect 38068 57264 38074 57316
rect 38120 57304 38148 57344
rect 38672 57344 45554 57372
rect 53887 57344 53932 57372
rect 38672 57304 38700 57344
rect 53926 57332 53932 57344
rect 53984 57332 53990 57384
rect 54297 57375 54355 57381
rect 54297 57341 54309 57375
rect 54343 57341 54355 57375
rect 54297 57335 54355 57341
rect 38120 57276 38700 57304
rect 40586 57264 40592 57316
rect 40644 57304 40650 57316
rect 45370 57304 45376 57316
rect 40644 57276 45376 57304
rect 40644 57264 40650 57276
rect 45370 57264 45376 57276
rect 45428 57264 45434 57316
rect 51074 57264 51080 57316
rect 51132 57304 51138 57316
rect 54312 57304 54340 57335
rect 58345 57307 58403 57313
rect 58345 57304 58357 57307
rect 51132 57276 54156 57304
rect 54312 57276 58357 57304
rect 51132 57264 51138 57276
rect 30374 57236 30380 57248
rect 25884 57208 26234 57236
rect 30335 57208 30380 57236
rect 30374 57196 30380 57208
rect 30432 57196 30438 57248
rect 31386 57196 31392 57248
rect 31444 57236 31450 57248
rect 32490 57236 32496 57248
rect 31444 57208 32496 57236
rect 31444 57196 31450 57208
rect 32490 57196 32496 57208
rect 32548 57196 32554 57248
rect 35342 57236 35348 57248
rect 35303 57208 35348 57236
rect 35342 57196 35348 57208
rect 35400 57196 35406 57248
rect 36354 57196 36360 57248
rect 36412 57236 36418 57248
rect 54018 57236 54024 57248
rect 36412 57208 54024 57236
rect 36412 57196 36418 57208
rect 54018 57196 54024 57208
rect 54076 57196 54082 57248
rect 54128 57236 54156 57276
rect 58345 57273 58357 57276
rect 58391 57273 58403 57307
rect 58345 57267 58403 57273
rect 55582 57236 55588 57248
rect 54128 57208 55588 57236
rect 55582 57196 55588 57208
rect 55640 57196 55646 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 1762 56992 1768 57044
rect 1820 57032 1826 57044
rect 31570 57032 31576 57044
rect 1820 57004 31576 57032
rect 1820 56992 1826 57004
rect 31570 56992 31576 57004
rect 31628 56992 31634 57044
rect 34514 56992 34520 57044
rect 34572 57032 34578 57044
rect 34974 57032 34980 57044
rect 34572 57004 34980 57032
rect 34572 56992 34578 57004
rect 34974 56992 34980 57004
rect 35032 57032 35038 57044
rect 36078 57032 36084 57044
rect 35032 57004 36084 57032
rect 35032 56992 35038 57004
rect 36078 56992 36084 57004
rect 36136 56992 36142 57044
rect 36630 56992 36636 57044
rect 36688 57032 36694 57044
rect 58250 57032 58256 57044
rect 36688 57004 58256 57032
rect 36688 56992 36694 57004
rect 58250 56992 58256 57004
rect 58308 56992 58314 57044
rect 22094 56924 22100 56976
rect 22152 56964 22158 56976
rect 22281 56967 22339 56973
rect 22281 56964 22293 56967
rect 22152 56936 22293 56964
rect 22152 56924 22158 56936
rect 22281 56933 22293 56936
rect 22327 56933 22339 56967
rect 22281 56927 22339 56933
rect 24854 56924 24860 56976
rect 24912 56964 24918 56976
rect 40586 56964 40592 56976
rect 24912 56936 40592 56964
rect 24912 56924 24918 56936
rect 40586 56924 40592 56936
rect 40644 56924 40650 56976
rect 43806 56924 43812 56976
rect 43864 56964 43870 56976
rect 43864 56936 44128 56964
rect 43864 56924 43870 56936
rect 2682 56856 2688 56908
rect 2740 56896 2746 56908
rect 32674 56896 32680 56908
rect 2740 56868 32680 56896
rect 2740 56856 2746 56868
rect 32674 56856 32680 56868
rect 32732 56856 32738 56908
rect 1670 56828 1676 56840
rect 1631 56800 1676 56828
rect 1670 56788 1676 56800
rect 1728 56788 1734 56840
rect 21634 56828 21640 56840
rect 21595 56800 21640 56828
rect 21634 56788 21640 56800
rect 21692 56788 21698 56840
rect 21726 56788 21732 56840
rect 21784 56828 21790 56840
rect 21784 56800 21829 56828
rect 21784 56788 21790 56800
rect 21910 56788 21916 56840
rect 21968 56828 21974 56840
rect 22186 56837 22192 56840
rect 22143 56831 22192 56837
rect 21968 56800 22013 56828
rect 21968 56788 21974 56800
rect 22143 56797 22155 56831
rect 22189 56797 22192 56831
rect 22143 56791 22192 56797
rect 22186 56788 22192 56791
rect 22244 56788 22250 56840
rect 29914 56788 29920 56840
rect 29972 56828 29978 56840
rect 38562 56828 38568 56840
rect 29972 56800 38568 56828
rect 29972 56788 29978 56800
rect 38562 56788 38568 56800
rect 38620 56788 38626 56840
rect 41046 56828 41052 56840
rect 38764 56800 41052 56828
rect 15746 56720 15752 56772
rect 15804 56760 15810 56772
rect 17126 56760 17132 56772
rect 15804 56732 17132 56760
rect 15804 56720 15810 56732
rect 17126 56720 17132 56732
rect 17184 56760 17190 56772
rect 20622 56760 20628 56772
rect 17184 56732 20628 56760
rect 17184 56720 17190 56732
rect 20622 56720 20628 56732
rect 20680 56720 20686 56772
rect 21358 56720 21364 56772
rect 21416 56760 21422 56772
rect 21818 56760 21824 56772
rect 21416 56732 21824 56760
rect 21416 56720 21422 56732
rect 21818 56720 21824 56732
rect 21876 56720 21882 56772
rect 22005 56763 22063 56769
rect 22005 56729 22017 56763
rect 22051 56760 22063 56763
rect 38764 56760 38792 56800
rect 41046 56788 41052 56800
rect 41104 56788 41110 56840
rect 43901 56831 43959 56837
rect 43901 56797 43913 56831
rect 43947 56797 43959 56831
rect 43901 56791 43959 56797
rect 43916 56760 43944 56791
rect 43990 56788 43996 56840
rect 44048 56788 44054 56840
rect 44100 56837 44128 56936
rect 54113 56899 54171 56905
rect 54113 56865 54125 56899
rect 54159 56896 54171 56899
rect 58345 56899 58403 56905
rect 58345 56896 58357 56899
rect 54159 56868 58357 56896
rect 54159 56865 54171 56868
rect 54113 56859 54171 56865
rect 58345 56865 58357 56868
rect 58391 56865 58403 56899
rect 58345 56859 58403 56865
rect 44085 56831 44143 56837
rect 44085 56797 44097 56831
rect 44131 56797 44143 56831
rect 44450 56828 44456 56840
rect 44411 56800 44456 56828
rect 44085 56791 44143 56797
rect 44450 56788 44456 56800
rect 44508 56788 44514 56840
rect 44545 56831 44603 56837
rect 44545 56797 44557 56831
rect 44591 56797 44603 56831
rect 54018 56828 54024 56840
rect 53979 56800 54024 56828
rect 44545 56791 44603 56797
rect 22051 56732 38792 56760
rect 39868 56732 43944 56760
rect 44008 56760 44036 56788
rect 44560 56760 44588 56791
rect 54018 56788 54024 56800
rect 54076 56788 54082 56840
rect 54386 56828 54392 56840
rect 54347 56800 54392 56828
rect 54386 56788 54392 56800
rect 54444 56788 54450 56840
rect 54570 56828 54576 56840
rect 54531 56800 54576 56828
rect 54570 56788 54576 56800
rect 54628 56788 54634 56840
rect 58158 56760 58164 56772
rect 44008 56732 44588 56760
rect 58119 56732 58164 56760
rect 22051 56729 22063 56732
rect 22005 56723 22063 56729
rect 1949 56695 2007 56701
rect 1949 56661 1961 56695
rect 1995 56692 2007 56695
rect 39868 56692 39896 56732
rect 58158 56720 58164 56732
rect 58216 56720 58222 56772
rect 1995 56664 39896 56692
rect 43717 56695 43775 56701
rect 1995 56661 2007 56664
rect 1949 56655 2007 56661
rect 43717 56661 43729 56695
rect 43763 56692 43775 56695
rect 43990 56692 43996 56704
rect 43763 56664 43996 56692
rect 43763 56661 43775 56664
rect 43717 56655 43775 56661
rect 43990 56652 43996 56664
rect 44048 56652 44054 56704
rect 53466 56692 53472 56704
rect 53427 56664 53472 56692
rect 53466 56652 53472 56664
rect 53524 56652 53530 56704
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 8570 56448 8576 56500
rect 8628 56488 8634 56500
rect 8628 56460 22094 56488
rect 8628 56448 8634 56460
rect 15654 56420 15660 56432
rect 15615 56392 15660 56420
rect 15654 56380 15660 56392
rect 15712 56380 15718 56432
rect 22066 56420 22094 56460
rect 29546 56448 29552 56500
rect 29604 56488 29610 56500
rect 48682 56488 48688 56500
rect 29604 56460 34100 56488
rect 29604 56448 29610 56460
rect 22066 56392 33732 56420
rect 1670 56352 1676 56364
rect 1631 56324 1676 56352
rect 1670 56312 1676 56324
rect 1728 56312 1734 56364
rect 9030 56312 9036 56364
rect 9088 56352 9094 56364
rect 15381 56355 15439 56361
rect 15381 56352 15393 56355
rect 9088 56324 15393 56352
rect 9088 56312 9094 56324
rect 15381 56321 15393 56324
rect 15427 56321 15439 56355
rect 15562 56352 15568 56364
rect 15523 56324 15568 56352
rect 15381 56315 15439 56321
rect 15562 56312 15568 56324
rect 15620 56312 15626 56364
rect 15746 56352 15752 56364
rect 15707 56324 15752 56352
rect 15746 56312 15752 56324
rect 15804 56312 15810 56364
rect 29454 56352 29460 56364
rect 29415 56324 29460 56352
rect 29454 56312 29460 56324
rect 29512 56312 29518 56364
rect 29638 56352 29644 56364
rect 29599 56324 29644 56352
rect 29638 56312 29644 56324
rect 29696 56312 29702 56364
rect 29914 56361 29920 56364
rect 29733 56355 29791 56361
rect 29733 56321 29745 56355
rect 29779 56321 29791 56355
rect 29733 56315 29791 56321
rect 29877 56355 29920 56361
rect 29877 56321 29889 56355
rect 29877 56315 29920 56321
rect 20990 56244 20996 56296
rect 21048 56284 21054 56296
rect 22002 56284 22008 56296
rect 21048 56256 22008 56284
rect 21048 56244 21054 56256
rect 22002 56244 22008 56256
rect 22060 56284 22066 56296
rect 29748 56284 29776 56315
rect 29914 56312 29920 56315
rect 29972 56312 29978 56364
rect 33594 56352 33600 56364
rect 33555 56324 33600 56352
rect 33594 56312 33600 56324
rect 33652 56312 33658 56364
rect 33704 56352 33732 56392
rect 33778 56380 33784 56432
rect 33836 56420 33842 56432
rect 34072 56420 34100 56460
rect 34716 56460 48688 56488
rect 34609 56423 34667 56429
rect 34609 56420 34621 56423
rect 33836 56392 33881 56420
rect 34072 56392 34621 56420
rect 33836 56380 33842 56392
rect 34609 56389 34621 56392
rect 34655 56389 34667 56423
rect 34609 56383 34667 56389
rect 33873 56355 33931 56361
rect 33873 56352 33885 56355
rect 33704 56324 33885 56352
rect 33873 56321 33885 56324
rect 33919 56321 33931 56355
rect 33873 56315 33931 56321
rect 33962 56312 33968 56364
rect 34020 56352 34026 56364
rect 34020 56324 34065 56352
rect 34020 56312 34026 56324
rect 34716 56284 34744 56460
rect 48682 56448 48688 56460
rect 48740 56448 48746 56500
rect 34974 56284 34980 56296
rect 22060 56256 29684 56284
rect 29748 56256 34744 56284
rect 34935 56256 34980 56284
rect 22060 56244 22066 56256
rect 15933 56219 15991 56225
rect 15933 56185 15945 56219
rect 15979 56216 15991 56219
rect 29546 56216 29552 56228
rect 15979 56188 29552 56216
rect 15979 56185 15991 56188
rect 15933 56179 15991 56185
rect 29546 56176 29552 56188
rect 29604 56176 29610 56228
rect 29656 56216 29684 56256
rect 34974 56244 34980 56256
rect 35032 56244 35038 56296
rect 33962 56216 33968 56228
rect 29656 56188 33968 56216
rect 33962 56176 33968 56188
rect 34020 56176 34026 56228
rect 34885 56219 34943 56225
rect 34885 56185 34897 56219
rect 34931 56216 34943 56219
rect 34931 56188 35894 56216
rect 34931 56185 34943 56188
rect 34885 56179 34943 56185
rect 1762 56148 1768 56160
rect 1723 56120 1768 56148
rect 1762 56108 1768 56120
rect 1820 56108 1826 56160
rect 28350 56108 28356 56160
rect 28408 56148 28414 56160
rect 29638 56148 29644 56160
rect 28408 56120 29644 56148
rect 28408 56108 28414 56120
rect 29638 56108 29644 56120
rect 29696 56108 29702 56160
rect 30009 56151 30067 56157
rect 30009 56117 30021 56151
rect 30055 56148 30067 56151
rect 30466 56148 30472 56160
rect 30055 56120 30472 56148
rect 30055 56117 30067 56120
rect 30009 56111 30067 56117
rect 30466 56108 30472 56120
rect 30524 56108 30530 56160
rect 34149 56151 34207 56157
rect 34149 56117 34161 56151
rect 34195 56148 34207 56151
rect 34747 56151 34805 56157
rect 34747 56148 34759 56151
rect 34195 56120 34759 56148
rect 34195 56117 34207 56120
rect 34149 56111 34207 56117
rect 34747 56117 34759 56120
rect 34793 56117 34805 56151
rect 34747 56111 34805 56117
rect 35253 56151 35311 56157
rect 35253 56117 35265 56151
rect 35299 56148 35311 56151
rect 35526 56148 35532 56160
rect 35299 56120 35532 56148
rect 35299 56117 35311 56120
rect 35253 56111 35311 56117
rect 35526 56108 35532 56120
rect 35584 56108 35590 56160
rect 35866 56148 35894 56188
rect 50062 56148 50068 56160
rect 35866 56120 50068 56148
rect 50062 56108 50068 56120
rect 50120 56108 50126 56160
rect 58342 56148 58348 56160
rect 58303 56120 58348 56148
rect 58342 56108 58348 56120
rect 58400 56108 58406 56160
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 1762 55904 1768 55956
rect 1820 55944 1826 55956
rect 29454 55944 29460 55956
rect 1820 55916 29460 55944
rect 1820 55904 1826 55916
rect 29454 55904 29460 55916
rect 29512 55904 29518 55956
rect 29638 55904 29644 55956
rect 29696 55944 29702 55956
rect 31386 55944 31392 55956
rect 29696 55916 31392 55944
rect 29696 55904 29702 55916
rect 31386 55904 31392 55916
rect 31444 55904 31450 55956
rect 43990 55904 43996 55956
rect 44048 55944 44054 55956
rect 44910 55944 44916 55956
rect 44048 55916 44916 55944
rect 44048 55904 44054 55916
rect 44910 55904 44916 55916
rect 44968 55904 44974 55956
rect 33594 55836 33600 55888
rect 33652 55876 33658 55888
rect 39390 55876 39396 55888
rect 33652 55848 39396 55876
rect 33652 55836 33658 55848
rect 39390 55836 39396 55848
rect 39448 55836 39454 55888
rect 1670 55672 1676 55684
rect 1631 55644 1676 55672
rect 1670 55632 1676 55644
rect 1728 55632 1734 55684
rect 1949 55607 2007 55613
rect 1949 55573 1961 55607
rect 1995 55604 2007 55607
rect 43438 55604 43444 55616
rect 1995 55576 43444 55604
rect 1995 55573 2007 55576
rect 1949 55567 2007 55573
rect 43438 55564 43444 55576
rect 43496 55564 43502 55616
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 1765 55403 1823 55409
rect 1765 55369 1777 55403
rect 1811 55400 1823 55403
rect 9122 55400 9128 55412
rect 1811 55372 9128 55400
rect 1811 55369 1823 55372
rect 1765 55363 1823 55369
rect 9122 55360 9128 55372
rect 9180 55360 9186 55412
rect 43257 55403 43315 55409
rect 43257 55369 43269 55403
rect 43303 55400 43315 55403
rect 43530 55400 43536 55412
rect 43303 55372 43536 55400
rect 43303 55369 43315 55372
rect 43257 55363 43315 55369
rect 43530 55360 43536 55372
rect 43588 55360 43594 55412
rect 1578 55264 1584 55276
rect 1539 55236 1584 55264
rect 1578 55224 1584 55236
rect 1636 55224 1642 55276
rect 43438 55264 43444 55276
rect 43399 55236 43444 55264
rect 43438 55224 43444 55236
rect 43496 55224 43502 55276
rect 43625 55267 43683 55273
rect 43625 55233 43637 55267
rect 43671 55264 43683 55267
rect 43806 55264 43812 55276
rect 43671 55236 43812 55264
rect 43671 55233 43683 55236
rect 43625 55227 43683 55233
rect 43806 55224 43812 55236
rect 43864 55224 43870 55276
rect 43993 55267 44051 55273
rect 43993 55233 44005 55267
rect 44039 55264 44051 55267
rect 47946 55264 47952 55276
rect 44039 55236 47952 55264
rect 44039 55233 44051 55236
rect 43993 55227 44051 55233
rect 47946 55224 47952 55236
rect 48004 55224 48010 55276
rect 43898 55196 43904 55208
rect 43859 55168 43904 55196
rect 43898 55156 43904 55168
rect 43956 55156 43962 55208
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 58342 54652 58348 54664
rect 58303 54624 58348 54652
rect 58342 54612 58348 54624
rect 58400 54612 58406 54664
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 1670 54176 1676 54188
rect 1631 54148 1676 54176
rect 1670 54136 1676 54148
rect 1728 54136 1734 54188
rect 43254 54176 43260 54188
rect 43215 54148 43260 54176
rect 43254 54136 43260 54148
rect 43312 54136 43318 54188
rect 43625 54179 43683 54185
rect 43625 54145 43637 54179
rect 43671 54176 43683 54179
rect 46934 54176 46940 54188
rect 43671 54148 46940 54176
rect 43671 54145 43683 54148
rect 43625 54139 43683 54145
rect 46934 54136 46940 54148
rect 46992 54136 46998 54188
rect 42702 54108 42708 54120
rect 42663 54080 42708 54108
rect 42702 54068 42708 54080
rect 42760 54068 42766 54120
rect 43073 54111 43131 54117
rect 43073 54077 43085 54111
rect 43119 54077 43131 54111
rect 43073 54071 43131 54077
rect 43533 54111 43591 54117
rect 43533 54077 43545 54111
rect 43579 54108 43591 54111
rect 43898 54108 43904 54120
rect 43579 54080 43904 54108
rect 43579 54077 43591 54080
rect 43533 54071 43591 54077
rect 1949 53975 2007 53981
rect 1949 53941 1961 53975
rect 1995 53972 2007 53975
rect 43088 53972 43116 54071
rect 43898 54068 43904 54080
rect 43956 54068 43962 54120
rect 1995 53944 43116 53972
rect 1995 53941 2007 53944
rect 1949 53935 2007 53941
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1578 53564 1584 53576
rect 1539 53536 1584 53564
rect 1578 53524 1584 53536
rect 1636 53524 1642 53576
rect 1765 53431 1823 53437
rect 1765 53397 1777 53431
rect 1811 53428 1823 53431
rect 18598 53428 18604 53440
rect 1811 53400 18604 53428
rect 1811 53397 1823 53400
rect 1765 53391 1823 53397
rect 18598 53388 18604 53400
rect 18656 53388 18662 53440
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 1946 53116 1952 53168
rect 2004 53156 2010 53168
rect 19334 53156 19340 53168
rect 2004 53128 19340 53156
rect 2004 53116 2010 53128
rect 19334 53116 19340 53128
rect 19392 53116 19398 53168
rect 1578 53088 1584 53100
rect 1539 53060 1584 53088
rect 1578 53048 1584 53060
rect 1636 53048 1642 53100
rect 1765 52887 1823 52893
rect 1765 52853 1777 52887
rect 1811 52884 1823 52887
rect 1854 52884 1860 52896
rect 1811 52856 1860 52884
rect 1811 52853 1823 52856
rect 1765 52847 1823 52853
rect 1854 52844 1860 52856
rect 1912 52844 1918 52896
rect 58342 52884 58348 52896
rect 58303 52856 58348 52884
rect 58342 52844 58348 52856
rect 58400 52844 58406 52896
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 44082 52640 44088 52692
rect 44140 52680 44146 52692
rect 46014 52680 46020 52692
rect 44140 52652 46020 52680
rect 44140 52640 44146 52652
rect 46014 52640 46020 52652
rect 46072 52640 46078 52692
rect 1857 52479 1915 52485
rect 1857 52445 1869 52479
rect 1903 52476 1915 52479
rect 5442 52476 5448 52488
rect 1903 52448 5448 52476
rect 1903 52445 1915 52448
rect 1857 52439 1915 52445
rect 5442 52436 5448 52448
rect 5500 52436 5506 52488
rect 1670 52408 1676 52420
rect 1631 52380 1676 52408
rect 1670 52368 1676 52380
rect 1728 52368 1734 52420
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 5442 52068 5448 52080
rect 5403 52040 5448 52068
rect 5442 52028 5448 52040
rect 5500 52028 5506 52080
rect 5166 52000 5172 52012
rect 5127 51972 5172 52000
rect 5166 51960 5172 51972
rect 5224 51960 5230 52012
rect 5353 52003 5411 52009
rect 5353 51969 5365 52003
rect 5399 51969 5411 52003
rect 5353 51963 5411 51969
rect 5589 52003 5647 52009
rect 5589 51969 5601 52003
rect 5635 52000 5647 52003
rect 15562 52000 15568 52012
rect 5635 51972 15568 52000
rect 5635 51969 5647 51972
rect 5589 51963 5647 51969
rect 4614 51892 4620 51944
rect 4672 51932 4678 51944
rect 5368 51932 5396 51963
rect 15562 51960 15568 51972
rect 15620 52000 15626 52012
rect 20438 52000 20444 52012
rect 15620 51972 20444 52000
rect 15620 51960 15626 51972
rect 20438 51960 20444 51972
rect 20496 51960 20502 52012
rect 4672 51904 5396 51932
rect 4672 51892 4678 51904
rect 5718 51796 5724 51808
rect 5679 51768 5724 51796
rect 5718 51756 5724 51768
rect 5776 51756 5782 51808
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 22186 51484 22192 51536
rect 22244 51524 22250 51536
rect 22244 51496 22692 51524
rect 22244 51484 22250 51496
rect 6886 51428 22600 51456
rect 1670 51320 1676 51332
rect 1631 51292 1676 51320
rect 1670 51280 1676 51292
rect 1728 51280 1734 51332
rect 1765 51255 1823 51261
rect 1765 51221 1777 51255
rect 1811 51252 1823 51255
rect 6886 51252 6914 51428
rect 22186 51348 22192 51400
rect 22244 51388 22250 51400
rect 22462 51388 22468 51400
rect 22244 51360 22468 51388
rect 22244 51348 22250 51360
rect 22462 51348 22468 51360
rect 22520 51348 22526 51400
rect 22572 51397 22600 51428
rect 22558 51391 22616 51397
rect 22558 51357 22570 51391
rect 22604 51357 22616 51391
rect 22664 51388 22692 51496
rect 23014 51397 23020 51400
rect 22971 51391 23020 51397
rect 22971 51388 22983 51391
rect 22664 51360 22983 51388
rect 22558 51351 22616 51357
rect 22971 51357 22983 51360
rect 23017 51357 23020 51391
rect 22971 51351 23020 51357
rect 23014 51348 23020 51351
rect 23072 51348 23078 51400
rect 58342 51388 58348 51400
rect 58303 51360 58348 51388
rect 58342 51348 58348 51360
rect 58400 51348 58406 51400
rect 20438 51280 20444 51332
rect 20496 51320 20502 51332
rect 22741 51323 22799 51329
rect 22741 51320 22753 51323
rect 20496 51292 22753 51320
rect 20496 51280 20502 51292
rect 22741 51289 22753 51292
rect 22787 51289 22799 51323
rect 22741 51283 22799 51289
rect 22833 51323 22891 51329
rect 22833 51289 22845 51323
rect 22879 51320 22891 51323
rect 43714 51320 43720 51332
rect 22879 51292 43720 51320
rect 22879 51289 22891 51292
rect 22833 51283 22891 51289
rect 43714 51280 43720 51292
rect 43772 51280 43778 51332
rect 23106 51252 23112 51264
rect 1811 51224 6914 51252
rect 23067 51224 23112 51252
rect 1811 51221 1823 51224
rect 1765 51215 1823 51221
rect 23106 51212 23112 51224
rect 23164 51212 23170 51264
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1670 50912 1676 50924
rect 1631 50884 1676 50912
rect 1670 50872 1676 50884
rect 1728 50872 1734 50924
rect 1857 50779 1915 50785
rect 1857 50745 1869 50779
rect 1903 50776 1915 50779
rect 8938 50776 8944 50788
rect 1903 50748 8944 50776
rect 1903 50745 1915 50748
rect 1857 50739 1915 50745
rect 8938 50736 8944 50748
rect 8996 50736 9002 50788
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 57790 50260 57796 50312
rect 57848 50300 57854 50312
rect 57885 50303 57943 50309
rect 57885 50300 57897 50303
rect 57848 50272 57897 50300
rect 57848 50260 57854 50272
rect 57885 50269 57897 50272
rect 57931 50269 57943 50303
rect 57885 50263 57943 50269
rect 1670 50232 1676 50244
rect 1631 50204 1676 50232
rect 1670 50192 1676 50204
rect 1728 50192 1734 50244
rect 58161 50235 58219 50241
rect 58161 50232 58173 50235
rect 57900 50204 58173 50232
rect 57900 50176 57928 50204
rect 58161 50201 58173 50204
rect 58207 50201 58219 50235
rect 58161 50195 58219 50201
rect 1765 50167 1823 50173
rect 1765 50133 1777 50167
rect 1811 50164 1823 50167
rect 20530 50164 20536 50176
rect 1811 50136 20536 50164
rect 1811 50133 1823 50136
rect 1765 50127 1823 50133
rect 20530 50124 20536 50136
rect 20588 50124 20594 50176
rect 57882 50124 57888 50176
rect 57940 50124 57946 50176
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 20438 49852 20444 49904
rect 20496 49892 20502 49904
rect 20806 49892 20812 49904
rect 20496 49864 20668 49892
rect 20767 49864 20812 49892
rect 20496 49852 20502 49864
rect 1670 49824 1676 49836
rect 1631 49796 1676 49824
rect 1670 49784 1676 49796
rect 1728 49784 1734 49836
rect 20530 49824 20536 49836
rect 20491 49796 20536 49824
rect 20530 49784 20536 49796
rect 20588 49784 20594 49836
rect 20640 49824 20668 49864
rect 20806 49852 20812 49864
rect 20864 49852 20870 49904
rect 20717 49827 20775 49833
rect 20717 49824 20729 49827
rect 20640 49796 20729 49824
rect 20717 49793 20729 49796
rect 20763 49793 20775 49827
rect 20717 49787 20775 49793
rect 20901 49827 20959 49833
rect 20901 49793 20913 49827
rect 20947 49793 20959 49827
rect 20901 49787 20959 49793
rect 1857 49759 1915 49765
rect 1857 49725 1869 49759
rect 1903 49756 1915 49759
rect 17862 49756 17868 49768
rect 1903 49728 17868 49756
rect 1903 49725 1915 49728
rect 1857 49719 1915 49725
rect 17862 49716 17868 49728
rect 17920 49716 17926 49768
rect 20622 49716 20628 49768
rect 20680 49756 20686 49768
rect 20916 49756 20944 49787
rect 20680 49728 20944 49756
rect 20680 49716 20686 49728
rect 21085 49623 21143 49629
rect 21085 49589 21097 49623
rect 21131 49620 21143 49623
rect 22002 49620 22008 49632
rect 21131 49592 22008 49620
rect 21131 49589 21143 49592
rect 21085 49583 21143 49589
rect 22002 49580 22008 49592
rect 22060 49580 22066 49632
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 21634 49376 21640 49428
rect 21692 49416 21698 49428
rect 21729 49419 21787 49425
rect 21729 49416 21741 49419
rect 21692 49388 21741 49416
rect 21692 49376 21698 49388
rect 21729 49385 21741 49388
rect 21775 49385 21787 49419
rect 21729 49379 21787 49385
rect 17862 49172 17868 49224
rect 17920 49212 17926 49224
rect 21177 49215 21235 49221
rect 21177 49212 21189 49215
rect 17920 49184 21189 49212
rect 17920 49172 17926 49184
rect 21177 49181 21189 49184
rect 21223 49181 21235 49215
rect 21542 49212 21548 49224
rect 21503 49184 21548 49212
rect 21177 49175 21235 49181
rect 21542 49172 21548 49184
rect 21600 49172 21606 49224
rect 20438 49104 20444 49156
rect 20496 49144 20502 49156
rect 21361 49147 21419 49153
rect 21361 49144 21373 49147
rect 20496 49116 21373 49144
rect 20496 49104 20502 49116
rect 21361 49113 21373 49116
rect 21407 49113 21419 49147
rect 21361 49107 21419 49113
rect 21450 49104 21456 49156
rect 21508 49144 21514 49156
rect 57974 49144 57980 49156
rect 21508 49116 21553 49144
rect 57935 49116 57980 49144
rect 21508 49104 21514 49116
rect 57974 49104 57980 49116
rect 58032 49104 58038 49156
rect 58345 49147 58403 49153
rect 58345 49113 58357 49147
rect 58391 49144 58403 49147
rect 58894 49144 58900 49156
rect 58391 49116 58900 49144
rect 58391 49113 58403 49116
rect 58345 49107 58403 49113
rect 58894 49104 58900 49116
rect 58952 49104 58958 49156
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 6886 48844 22140 48872
rect 3326 48764 3332 48816
rect 3384 48804 3390 48816
rect 6886 48804 6914 48844
rect 3384 48776 6914 48804
rect 19981 48807 20039 48813
rect 3384 48764 3390 48776
rect 19981 48773 19993 48807
rect 20027 48804 20039 48807
rect 20346 48804 20352 48816
rect 20027 48776 20352 48804
rect 20027 48773 20039 48776
rect 19981 48767 20039 48773
rect 20346 48764 20352 48776
rect 20404 48764 20410 48816
rect 1670 48736 1676 48748
rect 1631 48708 1676 48736
rect 1670 48696 1676 48708
rect 1728 48696 1734 48748
rect 19705 48739 19763 48745
rect 19705 48736 19717 48739
rect 6886 48708 19717 48736
rect 1765 48535 1823 48541
rect 1765 48501 1777 48535
rect 1811 48532 1823 48535
rect 6886 48532 6914 48708
rect 19705 48705 19717 48708
rect 19751 48705 19763 48739
rect 19705 48699 19763 48705
rect 19889 48739 19947 48745
rect 19889 48705 19901 48739
rect 19935 48705 19947 48739
rect 19889 48699 19947 48705
rect 19904 48668 19932 48699
rect 20070 48696 20076 48748
rect 20128 48736 20134 48748
rect 20622 48736 20628 48748
rect 20128 48708 20628 48736
rect 20128 48696 20134 48708
rect 20622 48696 20628 48708
rect 20680 48696 20686 48748
rect 22002 48736 22008 48748
rect 21963 48708 22008 48736
rect 22002 48696 22008 48708
rect 22060 48696 22066 48748
rect 22112 48745 22140 48844
rect 22204 48776 22508 48804
rect 22098 48739 22156 48745
rect 22098 48705 22110 48739
rect 22144 48705 22156 48739
rect 22098 48699 22156 48705
rect 20438 48668 20444 48680
rect 19904 48640 20444 48668
rect 20438 48628 20444 48640
rect 20496 48628 20502 48680
rect 20714 48628 20720 48680
rect 20772 48668 20778 48680
rect 21542 48668 21548 48680
rect 20772 48640 21548 48668
rect 20772 48628 20778 48640
rect 21542 48628 21548 48640
rect 21600 48668 21606 48680
rect 22204 48668 22232 48776
rect 22480 48745 22508 48776
rect 22281 48739 22339 48745
rect 22281 48705 22293 48739
rect 22327 48705 22339 48739
rect 22281 48699 22339 48705
rect 22373 48739 22431 48745
rect 22373 48705 22385 48739
rect 22419 48705 22431 48739
rect 22373 48699 22431 48705
rect 22470 48739 22528 48745
rect 22470 48705 22482 48739
rect 22516 48705 22528 48739
rect 22470 48699 22528 48705
rect 21600 48640 22232 48668
rect 21600 48628 21606 48640
rect 19978 48560 19984 48612
rect 20036 48600 20042 48612
rect 22296 48600 22324 48699
rect 22388 48668 22416 48699
rect 23017 48671 23075 48677
rect 23017 48668 23029 48671
rect 22388 48640 23029 48668
rect 23017 48637 23029 48640
rect 23063 48668 23075 48671
rect 39298 48668 39304 48680
rect 23063 48640 39304 48668
rect 23063 48637 23075 48640
rect 23017 48631 23075 48637
rect 39298 48628 39304 48640
rect 39356 48628 39362 48680
rect 24762 48600 24768 48612
rect 20036 48572 24768 48600
rect 20036 48560 20042 48572
rect 24762 48560 24768 48572
rect 24820 48560 24826 48612
rect 20254 48532 20260 48544
rect 1811 48504 6914 48532
rect 20215 48504 20260 48532
rect 1811 48501 1823 48504
rect 1765 48495 1823 48501
rect 20254 48492 20260 48504
rect 20312 48492 20318 48544
rect 22370 48492 22376 48544
rect 22428 48532 22434 48544
rect 22649 48535 22707 48541
rect 22649 48532 22661 48535
rect 22428 48504 22661 48532
rect 22428 48492 22434 48504
rect 22649 48501 22661 48504
rect 22695 48501 22707 48535
rect 22649 48495 22707 48501
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 21726 48220 21732 48272
rect 21784 48260 21790 48272
rect 22278 48260 22284 48272
rect 21784 48232 22284 48260
rect 21784 48220 21790 48232
rect 22278 48220 22284 48232
rect 22336 48220 22342 48272
rect 56870 48084 56876 48136
rect 56928 48124 56934 48136
rect 56965 48127 57023 48133
rect 56965 48124 56977 48127
rect 56928 48096 56977 48124
rect 56928 48084 56934 48096
rect 56965 48093 56977 48096
rect 57011 48093 57023 48127
rect 56965 48087 57023 48093
rect 1670 48056 1676 48068
rect 1631 48028 1676 48056
rect 1670 48016 1676 48028
rect 1728 48016 1734 48068
rect 57241 48059 57299 48065
rect 57241 48025 57253 48059
rect 57287 48056 57299 48059
rect 57330 48056 57336 48068
rect 57287 48028 57336 48056
rect 57287 48025 57299 48028
rect 57241 48019 57299 48025
rect 57330 48016 57336 48028
rect 57388 48016 57394 48068
rect 57974 48056 57980 48068
rect 57935 48028 57980 48056
rect 57974 48016 57980 48028
rect 58032 48016 58038 48068
rect 58342 48056 58348 48068
rect 58303 48028 58348 48056
rect 58342 48016 58348 48028
rect 58400 48016 58406 48068
rect 1765 47991 1823 47997
rect 1765 47957 1777 47991
rect 1811 47988 1823 47991
rect 16574 47988 16580 48000
rect 1811 47960 16580 47988
rect 1811 47957 1823 47960
rect 1765 47951 1823 47957
rect 16574 47948 16580 47960
rect 16632 47948 16638 48000
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1670 47648 1676 47660
rect 1631 47620 1676 47648
rect 1670 47608 1676 47620
rect 1728 47608 1734 47660
rect 21450 47608 21456 47660
rect 21508 47648 21514 47660
rect 41598 47648 41604 47660
rect 21508 47620 41604 47648
rect 21508 47608 21514 47620
rect 41598 47608 41604 47620
rect 41656 47608 41662 47660
rect 20346 47540 20352 47592
rect 20404 47580 20410 47592
rect 57054 47580 57060 47592
rect 20404 47552 57060 47580
rect 20404 47540 20410 47552
rect 57054 47540 57060 47552
rect 57112 47540 57118 47592
rect 1486 47404 1492 47456
rect 1544 47444 1550 47456
rect 1765 47447 1823 47453
rect 1765 47444 1777 47447
rect 1544 47416 1777 47444
rect 1544 47404 1550 47416
rect 1765 47413 1777 47416
rect 1811 47413 1823 47447
rect 1765 47407 1823 47413
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 1857 47039 1915 47045
rect 1857 47005 1869 47039
rect 1903 47036 1915 47039
rect 17218 47036 17224 47048
rect 1903 47008 17224 47036
rect 1903 47005 1915 47008
rect 1857 46999 1915 47005
rect 17218 46996 17224 47008
rect 17276 46996 17282 47048
rect 57606 46996 57612 47048
rect 57664 47036 57670 47048
rect 57885 47039 57943 47045
rect 57885 47036 57897 47039
rect 57664 47008 57897 47036
rect 57664 46996 57670 47008
rect 57885 47005 57897 47008
rect 57931 47005 57943 47039
rect 57885 46999 57943 47005
rect 1670 46968 1676 46980
rect 1631 46940 1676 46968
rect 1670 46928 1676 46940
rect 1728 46928 1734 46980
rect 58161 46971 58219 46977
rect 58161 46968 58173 46971
rect 57900 46940 58173 46968
rect 57900 46912 57928 46940
rect 58161 46937 58173 46940
rect 58207 46937 58219 46971
rect 58161 46931 58219 46937
rect 57882 46860 57888 46912
rect 57940 46860 57946 46912
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 21634 45976 21640 46028
rect 21692 46016 21698 46028
rect 28350 46016 28356 46028
rect 21692 45988 28356 46016
rect 21692 45976 21698 45988
rect 23032 45957 23060 45988
rect 28350 45976 28356 45988
rect 28408 45976 28414 46028
rect 22833 45951 22891 45957
rect 22833 45948 22845 45951
rect 6886 45920 22845 45948
rect 1670 45880 1676 45892
rect 1631 45852 1676 45880
rect 1670 45840 1676 45852
rect 1728 45840 1734 45892
rect 1765 45815 1823 45821
rect 1765 45781 1777 45815
rect 1811 45812 1823 45815
rect 6886 45812 6914 45920
rect 22833 45917 22845 45920
rect 22879 45917 22891 45951
rect 22833 45911 22891 45917
rect 23017 45951 23075 45957
rect 23017 45917 23029 45951
rect 23063 45917 23075 45951
rect 23198 45948 23204 45960
rect 23159 45920 23204 45948
rect 23017 45911 23075 45917
rect 23198 45908 23204 45920
rect 23256 45908 23262 45960
rect 23109 45883 23167 45889
rect 23109 45849 23121 45883
rect 23155 45880 23167 45883
rect 56778 45880 56784 45892
rect 23155 45852 56784 45880
rect 23155 45849 23167 45852
rect 23109 45843 23167 45849
rect 1811 45784 6914 45812
rect 22557 45815 22615 45821
rect 1811 45781 1823 45784
rect 1765 45775 1823 45781
rect 22557 45781 22569 45815
rect 22603 45812 22615 45815
rect 23124 45812 23152 45843
rect 56778 45840 56784 45852
rect 56836 45840 56842 45892
rect 57974 45880 57980 45892
rect 57935 45852 57980 45880
rect 57974 45840 57980 45852
rect 58032 45840 58038 45892
rect 58345 45883 58403 45889
rect 58345 45849 58357 45883
rect 58391 45880 58403 45883
rect 58710 45880 58716 45892
rect 58391 45852 58716 45880
rect 58391 45849 58403 45852
rect 58345 45843 58403 45849
rect 58710 45840 58716 45852
rect 58768 45840 58774 45892
rect 22603 45784 23152 45812
rect 22603 45781 22615 45784
rect 22557 45775 22615 45781
rect 23290 45772 23296 45824
rect 23348 45812 23354 45824
rect 23385 45815 23443 45821
rect 23385 45812 23397 45815
rect 23348 45784 23397 45812
rect 23348 45772 23354 45784
rect 23385 45781 23397 45784
rect 23431 45781 23443 45815
rect 23385 45775 23443 45781
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 21542 45568 21548 45620
rect 21600 45608 21606 45620
rect 23198 45608 23204 45620
rect 21600 45580 23204 45608
rect 21600 45568 21606 45580
rect 23198 45568 23204 45580
rect 23256 45568 23262 45620
rect 1578 45472 1584 45484
rect 1539 45444 1584 45472
rect 1578 45432 1584 45444
rect 1636 45432 1642 45484
rect 1765 45271 1823 45277
rect 1765 45237 1777 45271
rect 1811 45268 1823 45271
rect 24118 45268 24124 45280
rect 1811 45240 24124 45268
rect 1811 45237 1823 45240
rect 1765 45231 1823 45237
rect 24118 45228 24124 45240
rect 24176 45228 24182 45280
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 1857 44999 1915 45005
rect 1857 44965 1869 44999
rect 1903 44996 1915 44999
rect 9030 44996 9036 45008
rect 1903 44968 9036 44996
rect 1903 44965 1915 44968
rect 1857 44959 1915 44965
rect 9030 44956 9036 44968
rect 9088 44956 9094 45008
rect 31478 44888 31484 44940
rect 31536 44928 31542 44940
rect 45922 44928 45928 44940
rect 31536 44900 45928 44928
rect 31536 44888 31542 44900
rect 45922 44888 45928 44900
rect 45980 44888 45986 44940
rect 9122 44820 9128 44872
rect 9180 44860 9186 44872
rect 19426 44860 19432 44872
rect 9180 44832 19432 44860
rect 9180 44820 9186 44832
rect 19426 44820 19432 44832
rect 19484 44820 19490 44872
rect 21266 44820 21272 44872
rect 21324 44860 21330 44872
rect 54478 44860 54484 44872
rect 21324 44832 54484 44860
rect 21324 44820 21330 44832
rect 54478 44820 54484 44832
rect 54536 44820 54542 44872
rect 55950 44820 55956 44872
rect 56008 44860 56014 44872
rect 56965 44863 57023 44869
rect 56965 44860 56977 44863
rect 56008 44832 56977 44860
rect 56008 44820 56014 44832
rect 56965 44829 56977 44832
rect 57011 44829 57023 44863
rect 56965 44823 57023 44829
rect 1670 44792 1676 44804
rect 1631 44764 1676 44792
rect 1670 44752 1676 44764
rect 1728 44752 1734 44804
rect 57238 44792 57244 44804
rect 57199 44764 57244 44792
rect 57238 44752 57244 44764
rect 57296 44752 57302 44804
rect 57882 44752 57888 44804
rect 57940 44792 57946 44804
rect 57977 44795 58035 44801
rect 57977 44792 57989 44795
rect 57940 44764 57989 44792
rect 57940 44752 57946 44764
rect 57977 44761 57989 44764
rect 58023 44761 58035 44795
rect 57977 44755 58035 44761
rect 58345 44795 58403 44801
rect 58345 44761 58357 44795
rect 58391 44792 58403 44795
rect 58434 44792 58440 44804
rect 58391 44764 58440 44792
rect 58391 44761 58403 44764
rect 58345 44755 58403 44761
rect 58434 44752 58440 44764
rect 58492 44752 58498 44804
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 1670 44384 1676 44396
rect 1631 44356 1676 44384
rect 1670 44344 1676 44356
rect 1728 44344 1734 44396
rect 1765 44183 1823 44189
rect 1765 44149 1777 44183
rect 1811 44180 1823 44183
rect 15470 44180 15476 44192
rect 1811 44152 15476 44180
rect 1811 44149 1823 44152
rect 1765 44143 1823 44149
rect 15470 44140 15476 44152
rect 15528 44140 15534 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 15470 43840 15476 43852
rect 15431 43812 15476 43840
rect 15470 43800 15476 43812
rect 15528 43800 15534 43852
rect 15657 43775 15715 43781
rect 15657 43741 15669 43775
rect 15703 43741 15715 43775
rect 16022 43772 16028 43784
rect 15983 43744 16028 43772
rect 15657 43735 15715 43741
rect 15672 43704 15700 43735
rect 16022 43732 16028 43744
rect 16080 43732 16086 43784
rect 16209 43775 16267 43781
rect 16209 43741 16221 43775
rect 16255 43772 16267 43775
rect 20070 43772 20076 43784
rect 16255 43744 20076 43772
rect 16255 43741 16267 43744
rect 16209 43735 16267 43741
rect 20070 43732 20076 43744
rect 20128 43732 20134 43784
rect 47578 43732 47584 43784
rect 47636 43772 47642 43784
rect 57885 43775 57943 43781
rect 57885 43772 57897 43775
rect 47636 43744 57897 43772
rect 47636 43732 47642 43744
rect 57885 43741 57897 43744
rect 57931 43741 57943 43775
rect 57885 43735 57943 43741
rect 20438 43704 20444 43716
rect 15672 43676 20444 43704
rect 20438 43664 20444 43676
rect 20496 43704 20502 43716
rect 20622 43704 20628 43716
rect 20496 43676 20628 43704
rect 20496 43664 20502 43676
rect 20622 43664 20628 43676
rect 20680 43664 20686 43716
rect 58158 43704 58164 43716
rect 58119 43676 58164 43704
rect 58158 43664 58164 43676
rect 58216 43664 58222 43716
rect 15102 43636 15108 43648
rect 15063 43608 15108 43636
rect 15102 43596 15108 43608
rect 15160 43596 15166 43648
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 1578 43296 1584 43308
rect 1539 43268 1584 43296
rect 1578 43256 1584 43268
rect 1636 43256 1642 43308
rect 1765 43095 1823 43101
rect 1765 43061 1777 43095
rect 1811 43092 1823 43095
rect 4062 43092 4068 43104
rect 1811 43064 4068 43092
rect 1811 43061 1823 43064
rect 1765 43055 1823 43061
rect 4062 43052 4068 43064
rect 4120 43052 4126 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 30558 42780 30564 42832
rect 30616 42820 30622 42832
rect 32214 42820 32220 42832
rect 30616 42792 32220 42820
rect 30616 42780 30622 42792
rect 32214 42780 32220 42792
rect 32272 42780 32278 42832
rect 20070 42712 20076 42764
rect 20128 42752 20134 42764
rect 22830 42752 22836 42764
rect 20128 42724 22836 42752
rect 20128 42712 20134 42724
rect 22830 42712 22836 42724
rect 22888 42752 22894 42764
rect 23293 42755 23351 42761
rect 23293 42752 23305 42755
rect 22888 42724 23305 42752
rect 22888 42712 22894 42724
rect 23293 42721 23305 42724
rect 23339 42721 23351 42755
rect 23293 42715 23351 42721
rect 22738 42644 22744 42696
rect 22796 42684 22802 42696
rect 23017 42687 23075 42693
rect 23017 42684 23029 42687
rect 22796 42656 23029 42684
rect 22796 42644 22802 42656
rect 23017 42653 23029 42656
rect 23063 42684 23075 42687
rect 31846 42684 31852 42696
rect 23063 42656 31852 42684
rect 23063 42653 23075 42656
rect 23017 42647 23075 42653
rect 31846 42644 31852 42656
rect 31904 42644 31910 42696
rect 56962 42684 56968 42696
rect 56923 42656 56968 42684
rect 56962 42644 56968 42656
rect 57020 42644 57026 42696
rect 57882 42684 57888 42696
rect 57843 42656 57888 42684
rect 57882 42644 57888 42656
rect 57940 42644 57946 42696
rect 1670 42616 1676 42628
rect 1631 42588 1676 42616
rect 1670 42576 1676 42588
rect 1728 42576 1734 42628
rect 2041 42619 2099 42625
rect 2041 42585 2053 42619
rect 2087 42616 2099 42619
rect 5534 42616 5540 42628
rect 2087 42588 5540 42616
rect 2087 42585 2099 42588
rect 2041 42579 2099 42585
rect 5534 42576 5540 42588
rect 5592 42576 5598 42628
rect 31754 42576 31760 42628
rect 31812 42616 31818 42628
rect 57241 42619 57299 42625
rect 57241 42616 57253 42619
rect 31812 42588 57253 42616
rect 31812 42576 31818 42588
rect 57241 42585 57253 42588
rect 57287 42585 57299 42619
rect 57241 42579 57299 42585
rect 58161 42619 58219 42625
rect 58161 42585 58173 42619
rect 58207 42616 58219 42619
rect 58618 42616 58624 42628
rect 58207 42588 58624 42616
rect 58207 42585 58219 42588
rect 58161 42579 58219 42585
rect 58618 42576 58624 42588
rect 58676 42576 58682 42628
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 3786 42304 3792 42356
rect 3844 42344 3850 42356
rect 3844 42316 4844 42344
rect 3844 42304 3850 42316
rect 1857 42279 1915 42285
rect 1857 42245 1869 42279
rect 1903 42276 1915 42279
rect 4709 42279 4767 42285
rect 4709 42276 4721 42279
rect 1903 42248 4721 42276
rect 1903 42245 1915 42248
rect 1857 42239 1915 42245
rect 4709 42245 4721 42248
rect 4755 42245 4767 42279
rect 4709 42239 4767 42245
rect 1670 42208 1676 42220
rect 1631 42180 1676 42208
rect 1670 42168 1676 42180
rect 1728 42168 1734 42220
rect 4433 42211 4491 42217
rect 4433 42177 4445 42211
rect 4479 42177 4491 42211
rect 4614 42208 4620 42220
rect 4575 42180 4620 42208
rect 4433 42171 4491 42177
rect 4448 42140 4476 42171
rect 4614 42168 4620 42180
rect 4672 42168 4678 42220
rect 4816 42217 4844 42316
rect 4801 42211 4859 42217
rect 4801 42177 4813 42211
rect 4847 42177 4859 42211
rect 4801 42171 4859 42177
rect 22646 42168 22652 42220
rect 22704 42208 22710 42220
rect 22925 42211 22983 42217
rect 22925 42208 22937 42211
rect 22704 42180 22937 42208
rect 22704 42168 22710 42180
rect 22925 42177 22937 42180
rect 22971 42177 22983 42211
rect 23106 42208 23112 42220
rect 23067 42180 23112 42208
rect 22925 42171 22983 42177
rect 23106 42168 23112 42180
rect 23164 42168 23170 42220
rect 4890 42140 4896 42152
rect 4448 42112 4896 42140
rect 4890 42100 4896 42112
rect 4948 42100 4954 42152
rect 23477 42143 23535 42149
rect 23477 42109 23489 42143
rect 23523 42140 23535 42143
rect 27522 42140 27528 42152
rect 23523 42112 27528 42140
rect 23523 42109 23535 42112
rect 23477 42103 23535 42109
rect 27522 42100 27528 42112
rect 27580 42100 27586 42152
rect 4062 42032 4068 42084
rect 4120 42072 4126 42084
rect 32766 42072 32772 42084
rect 4120 42044 32772 42072
rect 4120 42032 4126 42044
rect 32766 42032 32772 42044
rect 32824 42032 32830 42084
rect 4982 42004 4988 42016
rect 4943 41976 4988 42004
rect 4982 41964 4988 41976
rect 5040 41964 5046 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 22646 41800 22652 41812
rect 22607 41772 22652 41800
rect 22646 41760 22652 41772
rect 22704 41760 22710 41812
rect 4982 41692 4988 41744
rect 5040 41732 5046 41744
rect 5040 41704 23152 41732
rect 5040 41692 5046 41704
rect 22830 41596 22836 41608
rect 22791 41568 22836 41596
rect 22830 41556 22836 41568
rect 22888 41556 22894 41608
rect 22922 41556 22928 41608
rect 22980 41596 22986 41608
rect 23124 41605 23152 41704
rect 23109 41599 23167 41605
rect 22980 41568 23025 41596
rect 22980 41556 22986 41568
rect 23109 41565 23121 41599
rect 23155 41565 23167 41599
rect 23109 41559 23167 41565
rect 23201 41599 23259 41605
rect 23201 41565 23213 41599
rect 23247 41596 23259 41599
rect 24854 41596 24860 41608
rect 23247 41568 24860 41596
rect 23247 41565 23259 41568
rect 23201 41559 23259 41565
rect 24854 41556 24860 41568
rect 24912 41556 24918 41608
rect 49142 41556 49148 41608
rect 49200 41596 49206 41608
rect 56965 41599 57023 41605
rect 56965 41596 56977 41599
rect 49200 41568 56977 41596
rect 49200 41556 49206 41568
rect 56965 41565 56977 41568
rect 57011 41565 57023 41599
rect 56965 41559 57023 41565
rect 1670 41528 1676 41540
rect 1631 41500 1676 41528
rect 1670 41488 1676 41500
rect 1728 41488 1734 41540
rect 1857 41531 1915 41537
rect 1857 41497 1869 41531
rect 1903 41528 1915 41531
rect 3970 41528 3976 41540
rect 1903 41500 3976 41528
rect 1903 41497 1915 41500
rect 1857 41491 1915 41497
rect 3970 41488 3976 41500
rect 4028 41488 4034 41540
rect 57238 41528 57244 41540
rect 57199 41500 57244 41528
rect 57238 41488 57244 41500
rect 57296 41488 57302 41540
rect 57882 41488 57888 41540
rect 57940 41528 57946 41540
rect 57977 41531 58035 41537
rect 57977 41528 57989 41531
rect 57940 41500 57989 41528
rect 57940 41488 57946 41500
rect 57977 41497 57989 41500
rect 58023 41497 58035 41531
rect 57977 41491 58035 41497
rect 58345 41531 58403 41537
rect 58345 41497 58357 41531
rect 58391 41528 58403 41531
rect 58802 41528 58808 41540
rect 58391 41500 58808 41528
rect 58391 41497 58403 41500
rect 58345 41491 58403 41497
rect 58802 41488 58808 41500
rect 58860 41488 58866 41540
rect 3878 41420 3884 41472
rect 3936 41460 3942 41472
rect 4614 41460 4620 41472
rect 3936 41432 4620 41460
rect 3936 41420 3942 41432
rect 4614 41420 4620 41432
rect 4672 41420 4678 41472
rect 31846 41420 31852 41472
rect 31904 41460 31910 41472
rect 32398 41460 32404 41472
rect 31904 41432 32404 41460
rect 31904 41420 31910 41432
rect 32398 41420 32404 41432
rect 32456 41420 32462 41472
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 2958 41216 2964 41268
rect 3016 41256 3022 41268
rect 3786 41256 3792 41268
rect 3016 41228 3792 41256
rect 3016 41216 3022 41228
rect 3786 41216 3792 41228
rect 3844 41256 3850 41268
rect 3844 41228 4108 41256
rect 3844 41216 3850 41228
rect 3970 41188 3976 41200
rect 3931 41160 3976 41188
rect 3970 41148 3976 41160
rect 4028 41148 4034 41200
rect 1394 41080 1400 41132
rect 1452 41120 1458 41132
rect 1673 41123 1731 41129
rect 1673 41120 1685 41123
rect 1452 41092 1685 41120
rect 1452 41080 1458 41092
rect 1673 41089 1685 41092
rect 1719 41089 1731 41123
rect 1673 41083 1731 41089
rect 3697 41123 3755 41129
rect 3697 41089 3709 41123
rect 3743 41089 3755 41123
rect 3878 41120 3884 41132
rect 3839 41092 3884 41120
rect 3697 41083 3755 41089
rect 3712 41052 3740 41083
rect 3878 41080 3884 41092
rect 3936 41080 3942 41132
rect 4080 41129 4108 41228
rect 4070 41123 4128 41129
rect 4070 41089 4082 41123
rect 4116 41089 4128 41123
rect 4070 41083 4128 41089
rect 4798 41052 4804 41064
rect 3712 41024 4804 41052
rect 4798 41012 4804 41024
rect 4856 41012 4862 41064
rect 5534 41012 5540 41064
rect 5592 41052 5598 41064
rect 5592 41024 12434 41052
rect 5592 41012 5598 41024
rect 1857 40987 1915 40993
rect 1857 40953 1869 40987
rect 1903 40984 1915 40987
rect 12406 40984 12434 41024
rect 18598 41012 18604 41064
rect 18656 41052 18662 41064
rect 22554 41052 22560 41064
rect 18656 41024 22560 41052
rect 18656 41012 18662 41024
rect 22554 41012 22560 41024
rect 22612 41012 22618 41064
rect 34422 40984 34428 40996
rect 1903 40956 11836 40984
rect 12406 40956 34428 40984
rect 1903 40953 1915 40956
rect 1857 40947 1915 40953
rect 4249 40919 4307 40925
rect 4249 40885 4261 40919
rect 4295 40916 4307 40919
rect 11698 40916 11704 40928
rect 4295 40888 11704 40916
rect 4295 40885 4307 40888
rect 4249 40879 4307 40885
rect 11698 40876 11704 40888
rect 11756 40876 11762 40928
rect 11808 40916 11836 40956
rect 34422 40944 34428 40956
rect 34480 40944 34486 40996
rect 22646 40916 22652 40928
rect 11808 40888 22652 40916
rect 22646 40876 22652 40888
rect 22704 40876 22710 40928
rect 27614 40876 27620 40928
rect 27672 40916 27678 40928
rect 34330 40916 34336 40928
rect 27672 40888 34336 40916
rect 27672 40876 27678 40888
rect 34330 40876 34336 40888
rect 34388 40876 34394 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 11698 40672 11704 40724
rect 11756 40712 11762 40724
rect 18046 40712 18052 40724
rect 11756 40684 18052 40712
rect 11756 40672 11762 40684
rect 18046 40672 18052 40684
rect 18104 40672 18110 40724
rect 22646 40508 22652 40520
rect 22607 40480 22652 40508
rect 22646 40468 22652 40480
rect 22704 40468 22710 40520
rect 23014 40508 23020 40520
rect 22975 40480 23020 40508
rect 23014 40468 23020 40480
rect 23072 40468 23078 40520
rect 48222 40468 48228 40520
rect 48280 40508 48286 40520
rect 57885 40511 57943 40517
rect 57885 40508 57897 40511
rect 48280 40480 57897 40508
rect 48280 40468 48286 40480
rect 57885 40477 57897 40480
rect 57931 40477 57943 40511
rect 57885 40471 57943 40477
rect 1670 40440 1676 40452
rect 1631 40412 1676 40440
rect 1670 40400 1676 40412
rect 1728 40400 1734 40452
rect 22830 40440 22836 40452
rect 22791 40412 22836 40440
rect 22830 40400 22836 40412
rect 22888 40400 22894 40452
rect 22925 40443 22983 40449
rect 22925 40409 22937 40443
rect 22971 40440 22983 40443
rect 28258 40440 28264 40452
rect 22971 40412 28264 40440
rect 22971 40409 22983 40412
rect 22925 40403 22983 40409
rect 28258 40400 28264 40412
rect 28316 40400 28322 40452
rect 58161 40443 58219 40449
rect 58161 40440 58173 40443
rect 57900 40412 58173 40440
rect 57900 40384 57928 40412
rect 58161 40409 58173 40412
rect 58207 40409 58219 40443
rect 58161 40403 58219 40409
rect 1765 40375 1823 40381
rect 1765 40341 1777 40375
rect 1811 40372 1823 40375
rect 2774 40372 2780 40384
rect 1811 40344 2780 40372
rect 1811 40341 1823 40344
rect 1765 40335 1823 40341
rect 2774 40332 2780 40344
rect 2832 40332 2838 40384
rect 23201 40375 23259 40381
rect 23201 40341 23213 40375
rect 23247 40372 23259 40375
rect 23474 40372 23480 40384
rect 23247 40344 23480 40372
rect 23247 40341 23259 40344
rect 23201 40335 23259 40341
rect 23474 40332 23480 40344
rect 23532 40332 23538 40384
rect 57882 40332 57888 40384
rect 57940 40332 57946 40384
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 3878 40168 3884 40180
rect 2608 40140 3884 40168
rect 1578 40060 1584 40112
rect 1636 40100 1642 40112
rect 1673 40103 1731 40109
rect 1673 40100 1685 40103
rect 1636 40072 1685 40100
rect 1636 40060 1642 40072
rect 1673 40069 1685 40072
rect 1719 40069 1731 40103
rect 1673 40063 1731 40069
rect 2406 40060 2412 40112
rect 2464 40100 2470 40112
rect 2464 40072 2544 40100
rect 2464 40060 2470 40072
rect 2516 40041 2544 40072
rect 2501 40035 2559 40041
rect 2501 40001 2513 40035
rect 2547 40001 2559 40035
rect 2608 40032 2636 40140
rect 3878 40128 3884 40140
rect 3936 40128 3942 40180
rect 2774 40100 2780 40112
rect 2735 40072 2780 40100
rect 2774 40060 2780 40072
rect 2832 40060 2838 40112
rect 58158 40100 58164 40112
rect 58119 40072 58164 40100
rect 58158 40060 58164 40072
rect 58216 40060 58222 40112
rect 2682 40032 2688 40044
rect 2608 40004 2688 40032
rect 2501 39995 2559 40001
rect 2682 39992 2688 40004
rect 2740 40032 2746 40044
rect 2958 40041 2964 40044
rect 2921 40035 2964 40041
rect 2740 40004 2833 40032
rect 2740 39992 2746 40004
rect 2921 40001 2933 40035
rect 2921 39995 2964 40001
rect 2958 39992 2964 39995
rect 3016 39992 3022 40044
rect 1857 39899 1915 39905
rect 1857 39865 1869 39899
rect 1903 39896 1915 39899
rect 1903 39868 6914 39896
rect 1903 39865 1915 39868
rect 1857 39859 1915 39865
rect 3050 39828 3056 39840
rect 3011 39800 3056 39828
rect 3050 39788 3056 39800
rect 3108 39788 3114 39840
rect 6886 39828 6914 39868
rect 22646 39828 22652 39840
rect 6886 39800 22652 39828
rect 22646 39788 22652 39800
rect 22704 39788 22710 39840
rect 56042 39788 56048 39840
rect 56100 39828 56106 39840
rect 58253 39831 58311 39837
rect 58253 39828 58265 39831
rect 56100 39800 58265 39828
rect 56100 39788 56106 39800
rect 58253 39797 58265 39800
rect 58299 39797 58311 39831
rect 58253 39791 58311 39797
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 3050 39584 3056 39636
rect 3108 39624 3114 39636
rect 22278 39624 22284 39636
rect 3108 39596 22284 39624
rect 3108 39584 3114 39596
rect 22278 39584 22284 39596
rect 22336 39584 22342 39636
rect 16574 39516 16580 39568
rect 16632 39556 16638 39568
rect 21910 39556 21916 39568
rect 16632 39528 21916 39556
rect 16632 39516 16638 39528
rect 21910 39516 21916 39528
rect 21968 39516 21974 39568
rect 23014 39448 23020 39500
rect 23072 39488 23078 39500
rect 23385 39491 23443 39497
rect 23385 39488 23397 39491
rect 23072 39460 23397 39488
rect 23072 39448 23078 39460
rect 23385 39457 23397 39460
rect 23431 39457 23443 39491
rect 23385 39451 23443 39457
rect 23106 39420 23112 39432
rect 23067 39392 23112 39420
rect 23106 39380 23112 39392
rect 23164 39380 23170 39432
rect 1394 39312 1400 39364
rect 1452 39352 1458 39364
rect 1673 39355 1731 39361
rect 1673 39352 1685 39355
rect 1452 39324 1685 39352
rect 1452 39312 1458 39324
rect 1673 39321 1685 39324
rect 1719 39321 1731 39355
rect 1673 39315 1731 39321
rect 1857 39355 1915 39361
rect 1857 39321 1869 39355
rect 1903 39352 1915 39355
rect 2498 39352 2504 39364
rect 1903 39324 2504 39352
rect 1903 39321 1915 39324
rect 1857 39315 1915 39321
rect 2498 39312 2504 39324
rect 2556 39312 2562 39364
rect 24854 39312 24860 39364
rect 24912 39352 24918 39364
rect 42518 39352 42524 39364
rect 24912 39324 42524 39352
rect 24912 39312 24918 39324
rect 42518 39312 42524 39324
rect 42576 39312 42582 39364
rect 57054 39352 57060 39364
rect 57015 39324 57060 39352
rect 57054 39312 57060 39324
rect 57112 39312 57118 39364
rect 57974 39352 57980 39364
rect 57935 39324 57980 39352
rect 57974 39312 57980 39324
rect 58032 39312 58038 39364
rect 58345 39355 58403 39361
rect 58345 39321 58357 39355
rect 58391 39352 58403 39355
rect 58526 39352 58532 39364
rect 58391 39324 58532 39352
rect 58391 39321 58403 39324
rect 58345 39315 58403 39321
rect 58526 39312 58532 39324
rect 58584 39312 58590 39364
rect 29638 39244 29644 39296
rect 29696 39284 29702 39296
rect 31754 39284 31760 39296
rect 29696 39256 31760 39284
rect 29696 39244 29702 39256
rect 31754 39244 31760 39256
rect 31812 39244 31818 39296
rect 37918 39244 37924 39296
rect 37976 39284 37982 39296
rect 57149 39287 57207 39293
rect 57149 39284 57161 39287
rect 37976 39256 57161 39284
rect 37976 39244 37982 39256
rect 57149 39253 57161 39256
rect 57195 39253 57207 39287
rect 57149 39247 57207 39253
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 20530 39040 20536 39092
rect 20588 39080 20594 39092
rect 22738 39080 22744 39092
rect 20588 39052 22744 39080
rect 20588 39040 20594 39052
rect 22738 39040 22744 39052
rect 22796 39040 22802 39092
rect 10318 38972 10324 39024
rect 10376 39012 10382 39024
rect 20809 39015 20867 39021
rect 20809 39012 20821 39015
rect 10376 38984 20821 39012
rect 10376 38972 10382 38984
rect 20809 38981 20821 38984
rect 20855 38981 20867 39015
rect 20809 38975 20867 38981
rect 22925 39015 22983 39021
rect 22925 38981 22937 39015
rect 22971 39012 22983 39015
rect 26878 39012 26884 39024
rect 22971 38984 26884 39012
rect 22971 38981 22983 38984
rect 22925 38975 22983 38981
rect 26878 38972 26884 38984
rect 26936 38972 26942 39024
rect 1670 38944 1676 38956
rect 1631 38916 1676 38944
rect 1670 38904 1676 38916
rect 1728 38904 1734 38956
rect 20438 38944 20444 38956
rect 20399 38916 20444 38944
rect 20438 38904 20444 38916
rect 20496 38904 20502 38956
rect 20589 38947 20647 38953
rect 20589 38913 20601 38947
rect 20635 38944 20647 38947
rect 20635 38913 20668 38944
rect 20589 38907 20668 38913
rect 20640 38876 20668 38907
rect 20714 38904 20720 38956
rect 20772 38944 20778 38956
rect 20990 38953 20996 38956
rect 20947 38947 20996 38953
rect 20772 38916 20817 38944
rect 20772 38904 20778 38916
rect 20947 38913 20959 38947
rect 20993 38913 20996 38947
rect 20947 38907 20996 38913
rect 20990 38904 20996 38907
rect 21048 38904 21054 38956
rect 22646 38944 22652 38956
rect 22607 38916 22652 38944
rect 22646 38904 22652 38916
rect 22704 38904 22710 38956
rect 22830 38944 22836 38956
rect 22791 38916 22836 38944
rect 22830 38904 22836 38916
rect 22888 38904 22894 38956
rect 23014 38904 23020 38956
rect 23072 38953 23078 38956
rect 23072 38944 23080 38953
rect 23072 38916 23117 38944
rect 23072 38907 23080 38916
rect 23072 38904 23078 38907
rect 26142 38876 26148 38888
rect 20640 38848 26148 38876
rect 26142 38836 26148 38848
rect 26200 38836 26206 38888
rect 20714 38768 20720 38820
rect 20772 38808 20778 38820
rect 24946 38808 24952 38820
rect 20772 38780 24952 38808
rect 20772 38768 20778 38780
rect 24946 38768 24952 38780
rect 25004 38768 25010 38820
rect 1765 38743 1823 38749
rect 1765 38709 1777 38743
rect 1811 38740 1823 38743
rect 11698 38740 11704 38752
rect 1811 38712 11704 38740
rect 1811 38709 1823 38712
rect 1765 38703 1823 38709
rect 11698 38700 11704 38712
rect 11756 38700 11762 38752
rect 21082 38740 21088 38752
rect 21043 38712 21088 38740
rect 21082 38700 21088 38712
rect 21140 38700 21146 38752
rect 23201 38743 23259 38749
rect 23201 38709 23213 38743
rect 23247 38740 23259 38743
rect 23842 38740 23848 38752
rect 23247 38712 23848 38740
rect 23247 38709 23259 38712
rect 23201 38703 23259 38709
rect 23842 38700 23848 38712
rect 23900 38700 23906 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 2958 38468 2964 38480
rect 2424 38440 2964 38468
rect 2424 38341 2452 38440
rect 2958 38428 2964 38440
rect 3016 38468 3022 38480
rect 3694 38468 3700 38480
rect 3016 38440 3700 38468
rect 3016 38428 3022 38440
rect 3694 38428 3700 38440
rect 3752 38428 3758 38480
rect 21082 38428 21088 38480
rect 21140 38468 21146 38480
rect 21453 38471 21511 38477
rect 21453 38468 21465 38471
rect 21140 38440 21465 38468
rect 21140 38428 21146 38440
rect 21453 38437 21465 38440
rect 21499 38437 21511 38471
rect 21453 38431 21511 38437
rect 21634 38428 21640 38480
rect 21692 38428 21698 38480
rect 2590 38360 2596 38412
rect 2648 38400 2654 38412
rect 2648 38372 3280 38400
rect 2648 38360 2654 38372
rect 2409 38335 2467 38341
rect 2409 38301 2421 38335
rect 2455 38301 2467 38335
rect 2409 38295 2467 38301
rect 2498 38292 2504 38344
rect 2556 38332 2562 38344
rect 2556 38304 2601 38332
rect 2556 38292 2562 38304
rect 2682 38292 2688 38344
rect 2740 38332 2746 38344
rect 2777 38335 2835 38341
rect 2777 38332 2789 38335
rect 2740 38304 2789 38332
rect 2740 38292 2746 38304
rect 2777 38301 2789 38304
rect 2823 38301 2835 38335
rect 2777 38295 2835 38301
rect 2866 38292 2872 38344
rect 2924 38332 2930 38344
rect 3252 38341 3280 38372
rect 18874 38360 18880 38412
rect 18932 38400 18938 38412
rect 20257 38403 20315 38409
rect 20257 38400 20269 38403
rect 18932 38372 20269 38400
rect 18932 38360 18938 38372
rect 20257 38369 20269 38372
rect 20303 38400 20315 38403
rect 20622 38400 20628 38412
rect 20303 38372 20628 38400
rect 20303 38369 20315 38372
rect 20257 38363 20315 38369
rect 20622 38360 20628 38372
rect 20680 38360 20686 38412
rect 21652 38400 21680 38428
rect 21197 38372 21680 38400
rect 3053 38335 3111 38341
rect 3053 38332 3065 38335
rect 2924 38304 3065 38332
rect 2924 38292 2930 38304
rect 3053 38301 3065 38304
rect 3099 38301 3111 38335
rect 3053 38295 3111 38301
rect 3237 38335 3295 38341
rect 3237 38301 3249 38335
rect 3283 38301 3295 38335
rect 3237 38295 3295 38301
rect 20073 38335 20131 38341
rect 20073 38301 20085 38335
rect 20119 38332 20131 38335
rect 21197 38332 21225 38372
rect 21468 38344 21496 38372
rect 21358 38332 21364 38344
rect 20119 38304 21225 38332
rect 21319 38304 21364 38332
rect 20119 38301 20131 38304
rect 20073 38295 20131 38301
rect 21358 38292 21364 38304
rect 21416 38292 21422 38344
rect 21450 38292 21456 38344
rect 21508 38292 21514 38344
rect 21634 38332 21640 38344
rect 21595 38304 21640 38332
rect 21634 38292 21640 38304
rect 21692 38292 21698 38344
rect 56965 38335 57023 38341
rect 56965 38301 56977 38335
rect 57011 38301 57023 38335
rect 57882 38332 57888 38344
rect 57843 38304 57888 38332
rect 56965 38295 57023 38301
rect 13906 38224 13912 38276
rect 13964 38264 13970 38276
rect 20990 38264 20996 38276
rect 13964 38236 20996 38264
rect 13964 38224 13970 38236
rect 20990 38224 20996 38236
rect 21048 38224 21054 38276
rect 2041 38199 2099 38205
rect 2041 38165 2053 38199
rect 2087 38196 2099 38199
rect 13998 38196 14004 38208
rect 2087 38168 14004 38196
rect 2087 38165 2099 38168
rect 2041 38159 2099 38165
rect 13998 38156 14004 38168
rect 14056 38156 14062 38208
rect 21818 38196 21824 38208
rect 21779 38168 21824 38196
rect 21818 38156 21824 38168
rect 21876 38156 21882 38208
rect 56980 38196 57008 38295
rect 57882 38292 57888 38304
rect 57940 38292 57946 38344
rect 57238 38264 57244 38276
rect 57199 38236 57244 38264
rect 57238 38224 57244 38236
rect 57296 38224 57302 38276
rect 58161 38267 58219 38273
rect 58161 38233 58173 38267
rect 58207 38264 58219 38267
rect 59078 38264 59084 38276
rect 58207 38236 59084 38264
rect 58207 38233 58219 38236
rect 58161 38227 58219 38233
rect 59078 38224 59084 38236
rect 59136 38224 59142 38276
rect 58250 38196 58256 38208
rect 56980 38168 58256 38196
rect 58250 38156 58256 38168
rect 58308 38156 58314 38208
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 2682 37992 2688 38004
rect 2643 37964 2688 37992
rect 2682 37952 2688 37964
rect 2740 37952 2746 38004
rect 56318 37992 56324 38004
rect 6886 37964 56324 37992
rect 1946 37884 1952 37936
rect 2004 37924 2010 37936
rect 2409 37927 2467 37933
rect 2409 37924 2421 37927
rect 2004 37896 2421 37924
rect 2004 37884 2010 37896
rect 2409 37893 2421 37896
rect 2455 37893 2467 37927
rect 6886 37924 6914 37964
rect 56318 37952 56324 37964
rect 56376 37952 56382 38004
rect 11974 37924 11980 37936
rect 2409 37887 2467 37893
rect 3620 37896 6914 37924
rect 11935 37896 11980 37924
rect 2133 37859 2191 37865
rect 2133 37825 2145 37859
rect 2179 37825 2191 37859
rect 2314 37856 2320 37868
rect 2275 37828 2320 37856
rect 2133 37819 2191 37825
rect 1857 37791 1915 37797
rect 1857 37757 1869 37791
rect 1903 37788 1915 37791
rect 2148 37788 2176 37819
rect 2314 37816 2320 37828
rect 2372 37816 2378 37868
rect 2498 37816 2504 37868
rect 2556 37856 2562 37868
rect 2556 37828 2601 37856
rect 2556 37816 2562 37828
rect 3620 37788 3648 37896
rect 11974 37884 11980 37896
rect 12032 37884 12038 37936
rect 13906 37924 13912 37936
rect 12084 37896 13912 37924
rect 3694 37816 3700 37868
rect 3752 37856 3758 37868
rect 11698 37856 11704 37868
rect 3752 37828 6914 37856
rect 11659 37828 11704 37856
rect 3752 37816 3758 37828
rect 1903 37760 3648 37788
rect 6886 37788 6914 37828
rect 11698 37816 11704 37828
rect 11756 37816 11762 37868
rect 12084 37865 12112 37896
rect 13906 37884 13912 37896
rect 13964 37884 13970 37936
rect 13998 37884 14004 37936
rect 14056 37924 14062 37936
rect 14056 37896 22876 37924
rect 14056 37884 14062 37896
rect 11885 37859 11943 37865
rect 11885 37825 11897 37859
rect 11931 37825 11943 37859
rect 11885 37819 11943 37825
rect 12069 37859 12127 37865
rect 12069 37825 12081 37859
rect 12115 37825 12127 37859
rect 12069 37819 12127 37825
rect 11330 37788 11336 37800
rect 6886 37760 11336 37788
rect 1903 37757 1915 37760
rect 1857 37751 1915 37757
rect 11330 37748 11336 37760
rect 11388 37788 11394 37800
rect 11900 37788 11928 37819
rect 17218 37816 17224 37868
rect 17276 37856 17282 37868
rect 18693 37859 18751 37865
rect 18693 37856 18705 37859
rect 17276 37828 18705 37856
rect 17276 37816 17282 37828
rect 18693 37825 18705 37828
rect 18739 37825 18751 37859
rect 18874 37856 18880 37868
rect 18835 37828 18880 37856
rect 18693 37819 18751 37825
rect 18874 37816 18880 37828
rect 18932 37816 18938 37868
rect 18966 37816 18972 37868
rect 19024 37856 19030 37868
rect 19107 37859 19165 37865
rect 19024 37828 19069 37856
rect 19024 37816 19030 37828
rect 19107 37825 19119 37859
rect 19153 37856 19165 37859
rect 19153 37828 19334 37856
rect 19153 37825 19165 37828
rect 19107 37819 19165 37825
rect 11388 37760 11928 37788
rect 18417 37791 18475 37797
rect 11388 37748 11394 37760
rect 18417 37757 18429 37791
rect 18463 37788 18475 37791
rect 18984 37788 19012 37816
rect 18463 37760 19012 37788
rect 19306 37788 19334 37828
rect 19702 37816 19708 37868
rect 19760 37856 19766 37868
rect 21450 37856 21456 37868
rect 19760 37828 19805 37856
rect 21411 37828 21456 37856
rect 19760 37816 19766 37828
rect 21450 37816 21456 37828
rect 21508 37816 21514 37868
rect 22186 37816 22192 37868
rect 22244 37856 22250 37868
rect 22281 37859 22339 37865
rect 22281 37856 22293 37859
rect 22244 37828 22293 37856
rect 22244 37816 22250 37828
rect 22281 37825 22293 37828
rect 22327 37856 22339 37859
rect 22646 37856 22652 37868
rect 22327 37828 22652 37856
rect 22327 37825 22339 37828
rect 22281 37819 22339 37825
rect 22646 37816 22652 37828
rect 22704 37816 22710 37868
rect 22848 37865 22876 37896
rect 26142 37884 26148 37936
rect 26200 37924 26206 37936
rect 41506 37924 41512 37936
rect 26200 37896 41512 37924
rect 26200 37884 26206 37896
rect 41506 37884 41512 37896
rect 41564 37884 41570 37936
rect 22741 37859 22799 37865
rect 22741 37825 22753 37859
rect 22787 37825 22799 37859
rect 22741 37819 22799 37825
rect 22833 37859 22891 37865
rect 22833 37825 22845 37859
rect 22879 37825 22891 37859
rect 23198 37856 23204 37868
rect 23159 37828 23204 37856
rect 22833 37819 22891 37825
rect 20806 37788 20812 37800
rect 19306 37760 20812 37788
rect 18463 37757 18475 37760
rect 18417 37751 18475 37757
rect 20806 37748 20812 37760
rect 20864 37748 20870 37800
rect 20898 37748 20904 37800
rect 20956 37788 20962 37800
rect 22756 37788 22784 37819
rect 23198 37816 23204 37828
rect 23256 37816 23262 37868
rect 23477 37791 23535 37797
rect 20956 37760 22094 37788
rect 22756 37760 22876 37788
rect 20956 37748 20962 37760
rect 12253 37723 12311 37729
rect 12253 37689 12265 37723
rect 12299 37720 12311 37723
rect 18782 37720 18788 37732
rect 12299 37692 18788 37720
rect 12299 37689 12311 37692
rect 12253 37683 12311 37689
rect 18782 37680 18788 37692
rect 18840 37680 18846 37732
rect 19245 37723 19303 37729
rect 19245 37689 19257 37723
rect 19291 37720 19303 37723
rect 20438 37720 20444 37732
rect 19291 37692 20444 37720
rect 19291 37689 19303 37692
rect 19245 37683 19303 37689
rect 20438 37680 20444 37692
rect 20496 37680 20502 37732
rect 17954 37612 17960 37664
rect 18012 37652 18018 37664
rect 18874 37652 18880 37664
rect 18012 37624 18880 37652
rect 18012 37612 18018 37624
rect 18874 37612 18880 37624
rect 18932 37612 18938 37664
rect 19702 37612 19708 37664
rect 19760 37652 19766 37664
rect 20346 37652 20352 37664
rect 19760 37624 20352 37652
rect 19760 37612 19766 37624
rect 20346 37612 20352 37624
rect 20404 37612 20410 37664
rect 22066 37652 22094 37760
rect 22848 37652 22876 37760
rect 23477 37757 23489 37791
rect 23523 37788 23535 37791
rect 26510 37788 26516 37800
rect 23523 37760 26516 37788
rect 23523 37757 23535 37760
rect 23477 37751 23535 37757
rect 26510 37748 26516 37760
rect 26568 37748 26574 37800
rect 22066 37624 22876 37652
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 20622 37408 20628 37460
rect 20680 37448 20686 37460
rect 21358 37448 21364 37460
rect 20680 37420 21364 37448
rect 20680 37408 20686 37420
rect 21358 37408 21364 37420
rect 21416 37408 21422 37460
rect 22465 37451 22523 37457
rect 22465 37417 22477 37451
rect 22511 37448 22523 37451
rect 23198 37448 23204 37460
rect 22511 37420 23204 37448
rect 22511 37417 22523 37420
rect 22465 37411 22523 37417
rect 23198 37408 23204 37420
rect 23256 37408 23262 37460
rect 41690 37408 41696 37460
rect 41748 37448 41754 37460
rect 48222 37448 48228 37460
rect 41748 37420 48228 37448
rect 41748 37408 41754 37420
rect 48222 37408 48228 37420
rect 48280 37408 48286 37460
rect 18966 37340 18972 37392
rect 19024 37380 19030 37392
rect 46934 37380 46940 37392
rect 19024 37352 46940 37380
rect 19024 37340 19030 37352
rect 46934 37340 46940 37352
rect 46992 37340 46998 37392
rect 2593 37315 2651 37321
rect 2593 37281 2605 37315
rect 2639 37312 2651 37315
rect 2639 37284 19472 37312
rect 2639 37281 2651 37284
rect 2593 37275 2651 37281
rect 1578 37244 1584 37256
rect 1539 37216 1584 37244
rect 1578 37204 1584 37216
rect 1636 37204 1642 37256
rect 19444 37253 19472 37284
rect 19996 37284 20668 37312
rect 19429 37247 19487 37253
rect 19429 37213 19441 37247
rect 19475 37213 19487 37247
rect 19702 37244 19708 37256
rect 19663 37216 19708 37244
rect 19429 37207 19487 37213
rect 19702 37204 19708 37216
rect 19760 37204 19766 37256
rect 19797 37247 19855 37253
rect 19797 37213 19809 37247
rect 19843 37244 19855 37247
rect 19996 37244 20024 37284
rect 20530 37244 20536 37256
rect 19843 37216 20024 37244
rect 20491 37216 20536 37244
rect 19843 37213 19855 37216
rect 19797 37207 19855 37213
rect 20530 37204 20536 37216
rect 20588 37204 20594 37256
rect 20640 37244 20668 37284
rect 20806 37272 20812 37324
rect 20864 37312 20870 37324
rect 20864 37284 22324 37312
rect 20864 37272 20870 37284
rect 21542 37244 21548 37256
rect 20640 37216 21548 37244
rect 21542 37204 21548 37216
rect 21600 37204 21606 37256
rect 21910 37244 21916 37256
rect 21871 37216 21916 37244
rect 21910 37204 21916 37216
rect 21968 37204 21974 37256
rect 22296 37253 22324 37284
rect 45020 37284 45324 37312
rect 22281 37247 22339 37253
rect 22281 37213 22293 37247
rect 22327 37244 22339 37247
rect 23014 37244 23020 37256
rect 22327 37216 23020 37244
rect 22327 37213 22339 37216
rect 22281 37207 22339 37213
rect 23014 37204 23020 37216
rect 23072 37204 23078 37256
rect 24118 37204 24124 37256
rect 24176 37244 24182 37256
rect 25590 37244 25596 37256
rect 24176 37216 25596 37244
rect 24176 37204 24182 37216
rect 25590 37204 25596 37216
rect 25648 37204 25654 37256
rect 36446 37204 36452 37256
rect 36504 37244 36510 37256
rect 45020 37244 45048 37284
rect 45186 37244 45192 37256
rect 36504 37216 45048 37244
rect 45147 37216 45192 37244
rect 36504 37204 36510 37216
rect 45186 37204 45192 37216
rect 45244 37204 45250 37256
rect 45296 37244 45324 37284
rect 45370 37272 45376 37324
rect 45428 37312 45434 37324
rect 45428 37284 46612 37312
rect 45428 37272 45434 37284
rect 45465 37247 45523 37253
rect 45465 37244 45477 37247
rect 45296 37216 45477 37244
rect 45465 37213 45477 37216
rect 45511 37213 45523 37247
rect 45465 37207 45523 37213
rect 45557 37247 45615 37253
rect 45557 37213 45569 37247
rect 45603 37213 45615 37247
rect 46477 37247 46535 37253
rect 46477 37244 46489 37247
rect 45557 37207 45615 37213
rect 45756 37216 46489 37244
rect 2406 37176 2412 37188
rect 2367 37148 2412 37176
rect 2406 37136 2412 37148
rect 2464 37136 2470 37188
rect 11330 37136 11336 37188
rect 11388 37176 11394 37188
rect 19613 37179 19671 37185
rect 19613 37176 19625 37179
rect 11388 37148 19625 37176
rect 11388 37136 11394 37148
rect 19613 37145 19625 37148
rect 19659 37145 19671 37179
rect 21269 37179 21327 37185
rect 21269 37176 21281 37179
rect 19613 37139 19671 37145
rect 19812 37148 21281 37176
rect 1765 37111 1823 37117
rect 1765 37077 1777 37111
rect 1811 37108 1823 37111
rect 2130 37108 2136 37120
rect 1811 37080 2136 37108
rect 1811 37077 1823 37080
rect 1765 37071 1823 37077
rect 2130 37068 2136 37080
rect 2188 37068 2194 37120
rect 19628 37108 19656 37139
rect 19812 37108 19840 37148
rect 21269 37145 21281 37148
rect 21315 37145 21327 37179
rect 21269 37139 21327 37145
rect 19628 37080 19840 37108
rect 19981 37111 20039 37117
rect 19981 37077 19993 37111
rect 20027 37108 20039 37111
rect 20714 37108 20720 37120
rect 20027 37080 20720 37108
rect 20027 37077 20039 37080
rect 19981 37071 20039 37077
rect 20714 37068 20720 37080
rect 20772 37068 20778 37120
rect 21284 37108 21312 37139
rect 21358 37136 21364 37188
rect 21416 37176 21422 37188
rect 22097 37179 22155 37185
rect 22097 37176 22109 37179
rect 21416 37148 22109 37176
rect 21416 37136 21422 37148
rect 22097 37145 22109 37148
rect 22143 37145 22155 37179
rect 22097 37139 22155 37145
rect 22186 37136 22192 37188
rect 22244 37176 22250 37188
rect 22244 37148 22289 37176
rect 22244 37136 22250 37148
rect 44082 37136 44088 37188
rect 44140 37176 44146 37188
rect 45373 37179 45431 37185
rect 45373 37176 45385 37179
rect 44140 37148 45385 37176
rect 44140 37136 44146 37148
rect 45373 37145 45385 37148
rect 45419 37145 45431 37179
rect 45373 37139 45431 37145
rect 22830 37108 22836 37120
rect 21284 37080 22836 37108
rect 22830 37068 22836 37080
rect 22888 37068 22894 37120
rect 43898 37068 43904 37120
rect 43956 37108 43962 37120
rect 45572 37108 45600 37207
rect 45646 37108 45652 37120
rect 43956 37080 45652 37108
rect 43956 37068 43962 37080
rect 45646 37068 45652 37080
rect 45704 37068 45710 37120
rect 45756 37117 45784 37216
rect 46477 37213 46489 37216
rect 46523 37213 46535 37247
rect 46584 37244 46612 37284
rect 46753 37247 46811 37253
rect 46753 37244 46765 37247
rect 46584 37216 46765 37244
rect 46477 37207 46535 37213
rect 46753 37213 46765 37216
rect 46799 37213 46811 37247
rect 46753 37207 46811 37213
rect 57698 37204 57704 37256
rect 57756 37244 57762 37256
rect 57885 37247 57943 37253
rect 57885 37244 57897 37247
rect 57756 37216 57897 37244
rect 57756 37204 57762 37216
rect 57885 37213 57897 37216
rect 57931 37213 57943 37247
rect 57885 37207 57943 37213
rect 46290 37176 46296 37188
rect 46251 37148 46296 37176
rect 46290 37136 46296 37148
rect 46348 37136 46354 37188
rect 58158 37176 58164 37188
rect 58119 37148 58164 37176
rect 58158 37136 58164 37148
rect 58216 37136 58222 37188
rect 45741 37111 45799 37117
rect 45741 37077 45753 37111
rect 45787 37077 45799 37111
rect 45741 37071 45799 37077
rect 46661 37111 46719 37117
rect 46661 37077 46673 37111
rect 46707 37108 46719 37111
rect 59170 37108 59176 37120
rect 46707 37080 59176 37108
rect 46707 37077 46719 37080
rect 46661 37071 46719 37077
rect 59170 37068 59176 37080
rect 59228 37068 59234 37120
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 18414 36864 18420 36916
rect 18472 36904 18478 36916
rect 20530 36904 20536 36916
rect 18472 36876 20536 36904
rect 18472 36864 18478 36876
rect 20530 36864 20536 36876
rect 20588 36864 20594 36916
rect 21361 36907 21419 36913
rect 20916 36876 21220 36904
rect 1762 36796 1768 36848
rect 1820 36836 1826 36848
rect 20441 36839 20499 36845
rect 1820 36808 6914 36836
rect 1820 36796 1826 36808
rect 1394 36728 1400 36780
rect 1452 36768 1458 36780
rect 1673 36771 1731 36777
rect 1673 36768 1685 36771
rect 1452 36740 1685 36768
rect 1452 36728 1458 36740
rect 1673 36737 1685 36740
rect 1719 36737 1731 36771
rect 1673 36731 1731 36737
rect 6886 36700 6914 36808
rect 20441 36805 20453 36839
rect 20487 36836 20499 36839
rect 20916 36836 20944 36876
rect 21082 36836 21088 36848
rect 20487 36808 20944 36836
rect 21043 36808 21088 36836
rect 20487 36805 20499 36808
rect 20441 36799 20499 36805
rect 20714 36768 20720 36780
rect 20675 36740 20720 36768
rect 20714 36728 20720 36740
rect 20772 36728 20778 36780
rect 20916 36777 20944 36808
rect 21082 36796 21088 36808
rect 21140 36796 21146 36848
rect 21192 36836 21220 36876
rect 21361 36873 21373 36907
rect 21407 36904 21419 36907
rect 21634 36904 21640 36916
rect 21407 36876 21640 36904
rect 21407 36873 21419 36876
rect 21361 36867 21419 36873
rect 21634 36864 21640 36876
rect 21692 36864 21698 36916
rect 26878 36904 26884 36916
rect 22066 36876 26884 36904
rect 22066 36836 22094 36876
rect 26878 36864 26884 36876
rect 26936 36864 26942 36916
rect 38930 36864 38936 36916
rect 38988 36904 38994 36916
rect 45370 36904 45376 36916
rect 38988 36876 45376 36904
rect 38988 36864 38994 36876
rect 45370 36864 45376 36876
rect 45428 36864 45434 36916
rect 21192 36808 22094 36836
rect 22186 36796 22192 36848
rect 22244 36836 22250 36848
rect 22244 36808 45554 36836
rect 22244 36796 22250 36808
rect 20865 36771 20944 36777
rect 20865 36737 20877 36771
rect 20911 36740 20944 36771
rect 20911 36737 20923 36740
rect 20865 36731 20923 36737
rect 20990 36728 20996 36780
rect 21048 36768 21054 36780
rect 21048 36740 21093 36768
rect 21048 36728 21054 36740
rect 21174 36728 21180 36780
rect 21232 36777 21238 36780
rect 21232 36768 21240 36777
rect 21232 36740 21277 36768
rect 21232 36731 21240 36740
rect 21232 36728 21238 36731
rect 23014 36728 23020 36780
rect 23072 36768 23078 36780
rect 23109 36771 23167 36777
rect 23109 36768 23121 36771
rect 23072 36740 23121 36768
rect 23072 36728 23078 36740
rect 23109 36737 23121 36740
rect 23155 36737 23167 36771
rect 23109 36731 23167 36737
rect 23201 36771 23259 36777
rect 23201 36737 23213 36771
rect 23247 36737 23259 36771
rect 23382 36768 23388 36780
rect 23343 36740 23388 36768
rect 23201 36731 23259 36737
rect 23216 36700 23244 36731
rect 23382 36728 23388 36740
rect 23440 36728 23446 36780
rect 23474 36728 23480 36780
rect 23532 36768 23538 36780
rect 23532 36740 23577 36768
rect 23532 36728 23538 36740
rect 43162 36728 43168 36780
rect 43220 36768 43226 36780
rect 45373 36771 45431 36777
rect 45373 36768 45385 36771
rect 43220 36740 45385 36768
rect 43220 36728 43226 36740
rect 45373 36737 45385 36740
rect 45419 36737 45431 36771
rect 45526 36768 45554 36808
rect 45646 36796 45652 36848
rect 45704 36836 45710 36848
rect 45704 36808 45749 36836
rect 45704 36796 45710 36808
rect 48682 36768 48688 36780
rect 45526 36740 48688 36768
rect 45373 36731 45431 36737
rect 48682 36728 48688 36740
rect 48740 36728 48746 36780
rect 36538 36700 36544 36712
rect 6886 36672 16712 36700
rect 23216 36672 36544 36700
rect 1765 36567 1823 36573
rect 1765 36533 1777 36567
rect 1811 36564 1823 36567
rect 12342 36564 12348 36576
rect 1811 36536 12348 36564
rect 1811 36533 1823 36536
rect 1765 36527 1823 36533
rect 12342 36524 12348 36536
rect 12400 36524 12406 36576
rect 16684 36564 16712 36672
rect 36538 36660 36544 36672
rect 36596 36660 36602 36712
rect 16758 36592 16764 36644
rect 16816 36632 16822 36644
rect 21082 36632 21088 36644
rect 16816 36604 21088 36632
rect 16816 36592 16822 36604
rect 21082 36592 21088 36604
rect 21140 36592 21146 36644
rect 26878 36592 26884 36644
rect 26936 36632 26942 36644
rect 58986 36632 58992 36644
rect 26936 36604 58992 36632
rect 26936 36592 26942 36604
rect 58986 36592 58992 36604
rect 59044 36592 59050 36644
rect 21634 36564 21640 36576
rect 16684 36536 21640 36564
rect 21634 36524 21640 36536
rect 21692 36524 21698 36576
rect 22646 36524 22652 36576
rect 22704 36564 22710 36576
rect 22925 36567 22983 36573
rect 22925 36564 22937 36567
rect 22704 36536 22937 36564
rect 22704 36524 22710 36536
rect 22925 36533 22937 36536
rect 22971 36533 22983 36567
rect 22925 36527 22983 36533
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1762 36360 1768 36372
rect 1723 36332 1768 36360
rect 1762 36320 1768 36332
rect 1820 36320 1826 36372
rect 12406 36332 18552 36360
rect 1854 36252 1860 36304
rect 1912 36292 1918 36304
rect 12406 36292 12434 36332
rect 1912 36264 12434 36292
rect 1912 36252 1918 36264
rect 2314 36184 2320 36236
rect 2372 36224 2378 36236
rect 2590 36224 2596 36236
rect 2372 36196 2596 36224
rect 2372 36184 2378 36196
rect 2590 36184 2596 36196
rect 2648 36224 2654 36236
rect 18524 36224 18552 36332
rect 27338 36320 27344 36372
rect 27396 36360 27402 36372
rect 46290 36360 46296 36372
rect 27396 36332 46296 36360
rect 27396 36320 27402 36332
rect 46290 36320 46296 36332
rect 46348 36320 46354 36372
rect 21913 36295 21971 36301
rect 21913 36261 21925 36295
rect 21959 36292 21971 36295
rect 22465 36295 22523 36301
rect 22465 36292 22477 36295
rect 21959 36264 22477 36292
rect 21959 36261 21971 36264
rect 21913 36255 21971 36261
rect 22465 36261 22477 36264
rect 22511 36261 22523 36295
rect 25130 36292 25136 36304
rect 25091 36264 25136 36292
rect 22465 36255 22523 36261
rect 25130 36252 25136 36264
rect 25188 36252 25194 36304
rect 32950 36292 32956 36304
rect 31726 36264 32956 36292
rect 31726 36224 31754 36264
rect 32950 36252 32956 36264
rect 33008 36252 33014 36304
rect 2648 36196 18368 36224
rect 18524 36196 24624 36224
rect 2648 36184 2654 36196
rect 18233 36159 18291 36165
rect 18233 36125 18245 36159
rect 18279 36125 18291 36159
rect 18233 36119 18291 36125
rect 1670 36088 1676 36100
rect 1631 36060 1676 36088
rect 1670 36048 1676 36060
rect 1728 36048 1734 36100
rect 18248 36020 18276 36119
rect 18340 36088 18368 36196
rect 18598 36156 18604 36168
rect 18559 36128 18604 36156
rect 18598 36116 18604 36128
rect 18656 36116 18662 36168
rect 21266 36116 21272 36168
rect 21324 36156 21330 36168
rect 21361 36159 21419 36165
rect 21361 36156 21373 36159
rect 21324 36128 21373 36156
rect 21324 36116 21330 36128
rect 21361 36125 21373 36128
rect 21407 36125 21419 36159
rect 21634 36156 21640 36168
rect 21595 36128 21640 36156
rect 21361 36119 21419 36125
rect 21634 36116 21640 36128
rect 21692 36116 21698 36168
rect 21729 36159 21787 36165
rect 21729 36125 21741 36159
rect 21775 36125 21787 36159
rect 22370 36156 22376 36168
rect 22331 36128 22376 36156
rect 21729 36119 21787 36125
rect 20990 36088 20996 36100
rect 18340 36060 20996 36088
rect 20990 36048 20996 36060
rect 21048 36048 21054 36100
rect 21450 36048 21456 36100
rect 21508 36088 21514 36100
rect 21545 36091 21603 36097
rect 21545 36088 21557 36091
rect 21508 36060 21557 36088
rect 21508 36048 21514 36060
rect 21545 36057 21557 36060
rect 21591 36057 21603 36091
rect 21744 36088 21772 36119
rect 22370 36116 22376 36128
rect 22428 36116 22434 36168
rect 22646 36156 22652 36168
rect 22607 36128 22652 36156
rect 22646 36116 22652 36128
rect 22704 36116 22710 36168
rect 24596 36165 24624 36196
rect 24780 36196 31754 36224
rect 24581 36159 24639 36165
rect 24581 36125 24593 36159
rect 24627 36125 24639 36159
rect 24581 36119 24639 36125
rect 24780 36100 24808 36196
rect 24946 36156 24952 36168
rect 24907 36128 24952 36156
rect 24946 36116 24952 36128
rect 25004 36116 25010 36168
rect 21545 36051 21603 36057
rect 21652 36060 21772 36088
rect 23109 36091 23167 36097
rect 20438 36020 20444 36032
rect 18248 35992 20444 36020
rect 20438 35980 20444 35992
rect 20496 35980 20502 36032
rect 21266 35980 21272 36032
rect 21324 36020 21330 36032
rect 21652 36020 21680 36060
rect 23109 36057 23121 36091
rect 23155 36057 23167 36091
rect 24762 36088 24768 36100
rect 24723 36060 24768 36088
rect 23109 36051 23167 36057
rect 21324 35992 21680 36020
rect 23124 36020 23152 36051
rect 24762 36048 24768 36060
rect 24820 36048 24826 36100
rect 24857 36091 24915 36097
rect 24857 36057 24869 36091
rect 24903 36088 24915 36091
rect 40862 36088 40868 36100
rect 24903 36060 40868 36088
rect 24903 36057 24915 36060
rect 24857 36051 24915 36057
rect 40862 36048 40868 36060
rect 40920 36048 40926 36100
rect 57974 36088 57980 36100
rect 57935 36060 57980 36088
rect 57974 36048 57980 36060
rect 58032 36048 58038 36100
rect 58345 36091 58403 36097
rect 58345 36057 58357 36091
rect 58391 36088 58403 36091
rect 59170 36088 59176 36100
rect 58391 36060 59176 36088
rect 58391 36057 58403 36060
rect 58345 36051 58403 36057
rect 59170 36048 59176 36060
rect 59228 36048 59234 36100
rect 26418 36020 26424 36032
rect 23124 35992 26424 36020
rect 21324 35980 21330 35992
rect 26418 35980 26424 35992
rect 26476 35980 26482 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 2222 35776 2228 35828
rect 2280 35816 2286 35828
rect 17954 35816 17960 35828
rect 2280 35788 17960 35816
rect 2280 35776 2286 35788
rect 17954 35776 17960 35788
rect 18012 35776 18018 35828
rect 20622 35816 20628 35828
rect 18156 35788 20628 35816
rect 1854 35708 1860 35760
rect 1912 35748 1918 35760
rect 2317 35751 2375 35757
rect 2317 35748 2329 35751
rect 1912 35720 2329 35748
rect 1912 35708 1918 35720
rect 2317 35717 2329 35720
rect 2363 35717 2375 35751
rect 18156 35748 18184 35788
rect 20622 35776 20628 35788
rect 20680 35776 20686 35828
rect 21453 35819 21511 35825
rect 21453 35785 21465 35819
rect 21499 35816 21511 35819
rect 22186 35816 22192 35828
rect 21499 35788 22192 35816
rect 21499 35785 21511 35788
rect 21453 35779 21511 35785
rect 22186 35776 22192 35788
rect 22244 35776 22250 35828
rect 35434 35776 35440 35828
rect 35492 35816 35498 35828
rect 38930 35816 38936 35828
rect 35492 35788 38936 35816
rect 35492 35776 35498 35788
rect 38930 35776 38936 35788
rect 38988 35776 38994 35828
rect 2317 35711 2375 35717
rect 6886 35720 18184 35748
rect 18233 35751 18291 35757
rect 2038 35680 2044 35692
rect 1999 35652 2044 35680
rect 2038 35640 2044 35652
rect 2096 35640 2102 35692
rect 2225 35683 2283 35689
rect 2225 35649 2237 35683
rect 2271 35649 2283 35683
rect 2225 35643 2283 35649
rect 2240 35612 2268 35643
rect 2406 35640 2412 35692
rect 2464 35689 2470 35692
rect 2464 35680 2472 35689
rect 2464 35652 2509 35680
rect 2464 35643 2472 35652
rect 2464 35640 2470 35643
rect 2682 35612 2688 35624
rect 2240 35584 2688 35612
rect 2682 35572 2688 35584
rect 2740 35612 2746 35624
rect 6886 35612 6914 35720
rect 18233 35717 18245 35751
rect 18279 35748 18291 35751
rect 20070 35748 20076 35760
rect 18279 35720 20076 35748
rect 18279 35717 18291 35720
rect 18233 35711 18291 35717
rect 20070 35708 20076 35720
rect 20128 35708 20134 35760
rect 20990 35708 20996 35760
rect 21048 35748 21054 35760
rect 21085 35751 21143 35757
rect 21085 35748 21097 35751
rect 21048 35720 21097 35748
rect 21048 35708 21054 35720
rect 21085 35717 21097 35720
rect 21131 35748 21143 35751
rect 36354 35748 36360 35760
rect 21131 35720 21496 35748
rect 21131 35717 21143 35720
rect 21085 35711 21143 35717
rect 18417 35683 18475 35689
rect 18417 35649 18429 35683
rect 18463 35649 18475 35683
rect 18417 35643 18475 35649
rect 2740 35584 6914 35612
rect 18432 35612 18460 35643
rect 18506 35640 18512 35692
rect 18564 35680 18570 35692
rect 18693 35683 18751 35689
rect 18564 35652 18609 35680
rect 18564 35640 18570 35652
rect 18693 35649 18705 35683
rect 18739 35649 18751 35683
rect 18693 35643 18751 35649
rect 18598 35612 18604 35624
rect 18432 35584 18604 35612
rect 2740 35572 2746 35584
rect 18598 35572 18604 35584
rect 18656 35572 18662 35624
rect 2593 35479 2651 35485
rect 2593 35445 2605 35479
rect 2639 35476 2651 35479
rect 4706 35476 4712 35488
rect 2639 35448 4712 35476
rect 2639 35445 2651 35448
rect 2593 35439 2651 35445
rect 4706 35436 4712 35448
rect 4764 35436 4770 35488
rect 18708 35476 18736 35643
rect 18782 35640 18788 35692
rect 18840 35680 18846 35692
rect 20806 35680 20812 35692
rect 18840 35652 18885 35680
rect 20767 35652 20812 35680
rect 18840 35640 18846 35652
rect 20806 35640 20812 35652
rect 20864 35640 20870 35692
rect 20902 35683 20960 35689
rect 20902 35649 20914 35683
rect 20948 35649 20960 35683
rect 20902 35643 20960 35649
rect 21177 35683 21235 35689
rect 21177 35649 21189 35683
rect 21223 35649 21235 35683
rect 21177 35643 21235 35649
rect 20533 35547 20591 35553
rect 20533 35513 20545 35547
rect 20579 35544 20591 35547
rect 20916 35544 20944 35643
rect 20990 35572 20996 35624
rect 21048 35612 21054 35624
rect 21192 35612 21220 35643
rect 21266 35640 21272 35692
rect 21324 35689 21330 35692
rect 21324 35680 21332 35689
rect 21324 35652 21369 35680
rect 21324 35643 21332 35652
rect 21324 35640 21330 35643
rect 21468 35624 21496 35720
rect 22020 35720 36360 35748
rect 22020 35692 22048 35720
rect 36354 35708 36360 35720
rect 36412 35708 36418 35760
rect 22002 35680 22008 35692
rect 21963 35652 22008 35680
rect 22002 35640 22008 35652
rect 22060 35640 22066 35692
rect 24854 35640 24860 35692
rect 24912 35680 24918 35692
rect 24949 35683 25007 35689
rect 24949 35680 24961 35683
rect 24912 35652 24961 35680
rect 24912 35640 24918 35652
rect 24949 35649 24961 35652
rect 24995 35649 25007 35683
rect 24949 35643 25007 35649
rect 25041 35683 25099 35689
rect 25041 35649 25053 35683
rect 25087 35680 25099 35683
rect 25130 35680 25136 35692
rect 25087 35652 25136 35680
rect 25087 35649 25099 35652
rect 25041 35643 25099 35649
rect 25130 35640 25136 35652
rect 25188 35640 25194 35692
rect 25314 35680 25320 35692
rect 25275 35652 25320 35680
rect 25314 35640 25320 35652
rect 25372 35640 25378 35692
rect 21048 35584 21220 35612
rect 21048 35572 21054 35584
rect 21450 35572 21456 35624
rect 21508 35612 21514 35624
rect 23201 35615 23259 35621
rect 23201 35612 23213 35615
rect 21508 35584 23213 35612
rect 21508 35572 21514 35584
rect 23201 35581 23213 35584
rect 23247 35612 23259 35615
rect 24026 35612 24032 35624
rect 23247 35584 24032 35612
rect 23247 35581 23259 35584
rect 23201 35575 23259 35581
rect 24026 35572 24032 35584
rect 24084 35572 24090 35624
rect 25406 35612 25412 35624
rect 25367 35584 25412 35612
rect 25406 35572 25412 35584
rect 25464 35572 25470 35624
rect 26878 35544 26884 35556
rect 20579 35516 26884 35544
rect 20579 35513 20591 35516
rect 20533 35507 20591 35513
rect 26878 35504 26884 35516
rect 26936 35504 26942 35556
rect 23566 35476 23572 35488
rect 18708 35448 23572 35476
rect 23566 35436 23572 35448
rect 23624 35436 23630 35488
rect 24302 35436 24308 35488
rect 24360 35476 24366 35488
rect 24397 35479 24455 35485
rect 24397 35476 24409 35479
rect 24360 35448 24409 35476
rect 24360 35436 24366 35448
rect 24397 35445 24409 35448
rect 24443 35445 24455 35479
rect 24397 35439 24455 35445
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 4706 35232 4712 35284
rect 4764 35272 4770 35284
rect 4764 35244 22094 35272
rect 4764 35232 4770 35244
rect 2593 35207 2651 35213
rect 2593 35173 2605 35207
rect 2639 35204 2651 35207
rect 2639 35176 21404 35204
rect 2639 35173 2651 35176
rect 2593 35167 2651 35173
rect 16390 35096 16396 35148
rect 16448 35136 16454 35148
rect 16448 35108 17080 35136
rect 16448 35096 16454 35108
rect 1486 35028 1492 35080
rect 1544 35068 1550 35080
rect 2041 35071 2099 35077
rect 2041 35068 2053 35071
rect 1544 35040 2053 35068
rect 1544 35028 1550 35040
rect 2041 35037 2053 35040
rect 2087 35037 2099 35071
rect 2222 35068 2228 35080
rect 2183 35040 2228 35068
rect 2041 35031 2099 35037
rect 2222 35028 2228 35040
rect 2280 35028 2286 35080
rect 2406 35028 2412 35080
rect 2464 35077 2470 35080
rect 2464 35068 2472 35077
rect 16206 35068 16212 35080
rect 2464 35040 16212 35068
rect 2464 35031 2472 35040
rect 2464 35028 2470 35031
rect 16206 35028 16212 35040
rect 16264 35028 16270 35080
rect 16298 35028 16304 35080
rect 16356 35068 16362 35080
rect 17052 35077 17080 35108
rect 21376 35077 21404 35176
rect 21542 35096 21548 35148
rect 21600 35136 21606 35148
rect 22066 35136 22094 35244
rect 22186 35232 22192 35284
rect 22244 35281 22250 35284
rect 22244 35275 22293 35281
rect 22244 35241 22247 35275
rect 22281 35241 22293 35275
rect 22244 35235 22293 35241
rect 22244 35232 22250 35235
rect 22370 35232 22376 35284
rect 22428 35272 22434 35284
rect 24854 35272 24860 35284
rect 22428 35244 22473 35272
rect 24815 35244 24860 35272
rect 22428 35232 22434 35244
rect 24854 35232 24860 35244
rect 24912 35232 24918 35284
rect 25222 35272 25228 35284
rect 25056 35244 25228 35272
rect 23753 35207 23811 35213
rect 23753 35173 23765 35207
rect 23799 35204 23811 35207
rect 24946 35204 24952 35216
rect 23799 35176 24952 35204
rect 23799 35173 23811 35176
rect 23753 35167 23811 35173
rect 24946 35164 24952 35176
rect 25004 35164 25010 35216
rect 22462 35136 22468 35148
rect 21600 35108 21680 35136
rect 22066 35108 22324 35136
rect 22423 35108 22468 35136
rect 21600 35096 21606 35108
rect 21652 35077 21680 35108
rect 16577 35071 16635 35077
rect 16356 35040 16401 35068
rect 16356 35028 16362 35040
rect 16577 35037 16589 35071
rect 16623 35037 16635 35071
rect 16577 35031 16635 35037
rect 16853 35071 16911 35077
rect 16853 35037 16865 35071
rect 16899 35037 16911 35071
rect 16853 35031 16911 35037
rect 17037 35071 17095 35077
rect 17037 35037 17049 35071
rect 17083 35037 17095 35071
rect 17037 35031 17095 35037
rect 21361 35071 21419 35077
rect 21361 35037 21373 35071
rect 21407 35037 21419 35071
rect 21361 35031 21419 35037
rect 21637 35071 21695 35077
rect 21637 35037 21649 35071
rect 21683 35037 21695 35071
rect 21637 35031 21695 35037
rect 2314 34960 2320 35012
rect 2372 35000 2378 35012
rect 2372 34972 2417 35000
rect 2372 34960 2378 34972
rect 15378 34960 15384 35012
rect 15436 35000 15442 35012
rect 15436 34972 15976 35000
rect 15436 34960 15442 34972
rect 15838 34932 15844 34944
rect 15799 34904 15844 34932
rect 15838 34892 15844 34904
rect 15896 34892 15902 34944
rect 15948 34932 15976 34972
rect 16592 34932 16620 35031
rect 16868 35000 16896 35031
rect 22094 35028 22100 35080
rect 22152 35068 22158 35080
rect 22296 35068 22324 35108
rect 22462 35096 22468 35108
rect 22520 35096 22526 35148
rect 24762 35136 24768 35148
rect 23860 35108 24768 35136
rect 23753 35071 23811 35077
rect 23753 35068 23765 35071
rect 22152 35040 22197 35068
rect 22296 35040 23765 35068
rect 22152 35028 22158 35040
rect 23753 35037 23765 35040
rect 23799 35037 23811 35071
rect 23753 35031 23811 35037
rect 18690 35000 18696 35012
rect 16868 34972 18696 35000
rect 18690 34960 18696 34972
rect 18748 34960 18754 35012
rect 20901 35003 20959 35009
rect 20901 34969 20913 35003
rect 20947 35000 20959 35003
rect 21545 35003 21603 35009
rect 21545 35000 21557 35003
rect 20947 34972 21557 35000
rect 20947 34969 20959 34972
rect 20901 34963 20959 34969
rect 21545 34969 21557 34972
rect 21591 35000 21603 35003
rect 23860 35000 23888 35108
rect 24762 35096 24768 35108
rect 24820 35096 24826 35148
rect 24026 35028 24032 35080
rect 24084 35068 24090 35080
rect 24854 35068 24860 35080
rect 24084 35040 24860 35068
rect 24084 35028 24090 35040
rect 24854 35028 24860 35040
rect 24912 35028 24918 35080
rect 25056 35077 25084 35244
rect 25222 35232 25228 35244
rect 25280 35232 25286 35284
rect 25332 35176 31754 35204
rect 25332 35136 25360 35176
rect 25204 35108 25360 35136
rect 25204 35078 25232 35108
rect 25498 35096 25504 35148
rect 25556 35096 25562 35148
rect 25148 35077 25232 35078
rect 25041 35071 25099 35077
rect 25041 35037 25053 35071
rect 25087 35037 25099 35071
rect 25041 35031 25099 35037
rect 25133 35071 25232 35077
rect 25133 35037 25145 35071
rect 25179 35050 25232 35071
rect 25317 35071 25375 35077
rect 25179 35037 25191 35050
rect 25133 35031 25191 35037
rect 25317 35037 25329 35071
rect 25363 35037 25375 35071
rect 25317 35031 25375 35037
rect 25409 35071 25467 35077
rect 25409 35037 25421 35071
rect 25455 35068 25467 35071
rect 25516 35068 25544 35096
rect 25455 35040 25544 35068
rect 31726 35068 31754 35176
rect 36538 35164 36544 35216
rect 36596 35204 36602 35216
rect 49878 35204 49884 35216
rect 36596 35176 49884 35204
rect 36596 35164 36602 35176
rect 49878 35164 49884 35176
rect 49936 35164 49942 35216
rect 47670 35068 47676 35080
rect 31726 35040 47676 35068
rect 25455 35037 25467 35040
rect 25409 35031 25467 35037
rect 21591 34972 23888 35000
rect 23937 35003 23995 35009
rect 21591 34969 21603 34972
rect 21545 34963 21603 34969
rect 23937 34969 23949 35003
rect 23983 35000 23995 35003
rect 24118 35000 24124 35012
rect 23983 34972 24124 35000
rect 23983 34969 23995 34972
rect 23937 34963 23995 34969
rect 21174 34932 21180 34944
rect 15948 34904 16620 34932
rect 21135 34904 21180 34932
rect 21174 34892 21180 34904
rect 21232 34892 21238 34944
rect 22738 34932 22744 34944
rect 22699 34904 22744 34932
rect 22738 34892 22744 34904
rect 22796 34892 22802 34944
rect 23477 34935 23535 34941
rect 23477 34901 23489 34935
rect 23523 34932 23535 34935
rect 23952 34932 23980 34963
rect 24118 34960 24124 34972
rect 24176 34960 24182 35012
rect 24210 34960 24216 35012
rect 24268 35000 24274 35012
rect 25332 35000 25360 35031
rect 47670 35028 47676 35040
rect 47728 35028 47734 35080
rect 51718 35028 51724 35080
rect 51776 35068 51782 35080
rect 57885 35071 57943 35077
rect 57885 35068 57897 35071
rect 51776 35040 57897 35068
rect 51776 35028 51782 35040
rect 57885 35037 57897 35040
rect 57931 35037 57943 35071
rect 58066 35068 58072 35080
rect 57885 35031 57943 35037
rect 57992 35040 58072 35068
rect 24268 34972 25360 35000
rect 24268 34960 24274 34972
rect 25498 34960 25504 35012
rect 25556 35000 25562 35012
rect 57992 35000 58020 35040
rect 58066 35028 58072 35040
rect 58124 35028 58130 35080
rect 58158 35000 58164 35012
rect 25556 34972 58020 35000
rect 58119 34972 58164 35000
rect 25556 34960 25562 34972
rect 58158 34960 58164 34972
rect 58216 34960 58222 35012
rect 23523 34904 23980 34932
rect 23523 34901 23535 34904
rect 23477 34895 23535 34901
rect 24762 34892 24768 34944
rect 24820 34932 24826 34944
rect 57146 34932 57152 34944
rect 24820 34904 57152 34932
rect 24820 34892 24826 34904
rect 57146 34892 57152 34904
rect 57204 34892 57210 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 15838 34688 15844 34740
rect 15896 34728 15902 34740
rect 27614 34728 27620 34740
rect 15896 34700 27620 34728
rect 15896 34688 15902 34700
rect 27614 34688 27620 34700
rect 27672 34688 27678 34740
rect 1857 34663 1915 34669
rect 1857 34629 1869 34663
rect 1903 34660 1915 34663
rect 20990 34660 20996 34672
rect 1903 34632 20996 34660
rect 1903 34629 1915 34632
rect 1857 34623 1915 34629
rect 20990 34620 20996 34632
rect 21048 34620 21054 34672
rect 21266 34660 21272 34672
rect 21100 34632 21272 34660
rect 1670 34592 1676 34604
rect 1631 34564 1676 34592
rect 1670 34552 1676 34564
rect 1728 34552 1734 34604
rect 16206 34552 16212 34604
rect 16264 34592 16270 34604
rect 17954 34592 17960 34604
rect 16264 34564 17960 34592
rect 16264 34552 16270 34564
rect 17954 34552 17960 34564
rect 18012 34592 18018 34604
rect 21100 34592 21128 34632
rect 21266 34620 21272 34632
rect 21324 34620 21330 34672
rect 24762 34660 24768 34672
rect 22296 34632 24768 34660
rect 18012 34564 21128 34592
rect 18012 34552 18018 34564
rect 21174 34552 21180 34604
rect 21232 34592 21238 34604
rect 22296 34601 22324 34632
rect 24762 34620 24768 34632
rect 24820 34620 24826 34672
rect 24854 34620 24860 34672
rect 24912 34660 24918 34672
rect 35434 34660 35440 34672
rect 24912 34632 35440 34660
rect 24912 34620 24918 34632
rect 35434 34620 35440 34632
rect 35492 34620 35498 34672
rect 22005 34595 22063 34601
rect 22005 34592 22017 34595
rect 21232 34564 22017 34592
rect 21232 34552 21238 34564
rect 22005 34561 22017 34564
rect 22051 34561 22063 34595
rect 22005 34555 22063 34561
rect 22281 34595 22339 34601
rect 22281 34561 22293 34595
rect 22327 34561 22339 34595
rect 22281 34555 22339 34561
rect 22664 34564 23244 34592
rect 18690 34484 18696 34536
rect 18748 34524 18754 34536
rect 21910 34524 21916 34536
rect 18748 34496 21916 34524
rect 18748 34484 18754 34496
rect 21910 34484 21916 34496
rect 21968 34524 21974 34536
rect 22664 34524 22692 34564
rect 21968 34496 22692 34524
rect 22741 34527 22799 34533
rect 21968 34484 21974 34496
rect 22741 34493 22753 34527
rect 22787 34524 22799 34527
rect 23106 34524 23112 34536
rect 22787 34496 23112 34524
rect 22787 34493 22799 34496
rect 22741 34487 22799 34493
rect 23106 34484 23112 34496
rect 23164 34484 23170 34536
rect 23216 34524 23244 34564
rect 23382 34552 23388 34604
rect 23440 34592 23446 34604
rect 23658 34592 23664 34604
rect 23440 34564 23664 34592
rect 23440 34552 23446 34564
rect 23658 34552 23664 34564
rect 23716 34552 23722 34604
rect 23842 34592 23848 34604
rect 23803 34564 23848 34592
rect 23842 34552 23848 34564
rect 23900 34552 23906 34604
rect 24397 34595 24455 34601
rect 24397 34561 24409 34595
rect 24443 34592 24455 34595
rect 24946 34592 24952 34604
rect 24443 34564 24808 34592
rect 24907 34564 24952 34592
rect 24443 34561 24455 34564
rect 24397 34555 24455 34561
rect 23216 34496 24440 34524
rect 20070 34416 20076 34468
rect 20128 34456 20134 34468
rect 22097 34459 22155 34465
rect 22097 34456 22109 34459
rect 20128 34428 22109 34456
rect 20128 34416 20134 34428
rect 22097 34425 22109 34428
rect 22143 34425 22155 34459
rect 22097 34419 22155 34425
rect 23658 34416 23664 34468
rect 23716 34456 23722 34468
rect 24210 34456 24216 34468
rect 23716 34428 24216 34456
rect 23716 34416 23722 34428
rect 24210 34416 24216 34428
rect 24268 34416 24274 34468
rect 24412 34456 24440 34496
rect 24486 34484 24492 34536
rect 24544 34524 24550 34536
rect 24581 34527 24639 34533
rect 24581 34524 24593 34527
rect 24544 34496 24593 34524
rect 24544 34484 24550 34496
rect 24581 34493 24593 34496
rect 24627 34493 24639 34527
rect 24780 34524 24808 34564
rect 24946 34552 24952 34564
rect 25004 34552 25010 34604
rect 25682 34524 25688 34536
rect 24780 34496 25688 34524
rect 24581 34487 24639 34493
rect 25682 34484 25688 34496
rect 25740 34484 25746 34536
rect 26878 34484 26884 34536
rect 26936 34524 26942 34536
rect 56410 34524 56416 34536
rect 26936 34496 56416 34524
rect 26936 34484 26942 34496
rect 56410 34484 56416 34496
rect 56468 34484 56474 34536
rect 25406 34456 25412 34468
rect 24412 34428 25412 34456
rect 25406 34416 25412 34428
rect 25464 34416 25470 34468
rect 32950 34348 32956 34400
rect 33008 34388 33014 34400
rect 34606 34388 34612 34400
rect 33008 34360 34612 34388
rect 33008 34348 33014 34360
rect 34606 34348 34612 34360
rect 34664 34388 34670 34400
rect 43254 34388 43260 34400
rect 34664 34360 43260 34388
rect 34664 34348 34670 34360
rect 43254 34348 43260 34360
rect 43312 34348 43318 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 20254 34144 20260 34196
rect 20312 34184 20318 34196
rect 21174 34184 21180 34196
rect 20312 34156 21180 34184
rect 20312 34144 20318 34156
rect 21174 34144 21180 34156
rect 21232 34144 21238 34196
rect 21634 34144 21640 34196
rect 21692 34184 21698 34196
rect 21692 34156 22232 34184
rect 21692 34144 21698 34156
rect 1854 34116 1860 34128
rect 1815 34088 1860 34116
rect 1854 34076 1860 34088
rect 1912 34076 1918 34128
rect 5718 34076 5724 34128
rect 5776 34116 5782 34128
rect 22204 34116 22232 34156
rect 22462 34144 22468 34196
rect 22520 34184 22526 34196
rect 22557 34187 22615 34193
rect 22557 34184 22569 34187
rect 22520 34156 22569 34184
rect 22520 34144 22526 34156
rect 22557 34153 22569 34156
rect 22603 34153 22615 34187
rect 22557 34147 22615 34153
rect 23124 34156 41368 34184
rect 23124 34116 23152 34156
rect 5776 34088 21956 34116
rect 22204 34088 23152 34116
rect 5776 34076 5782 34088
rect 12342 34008 12348 34060
rect 12400 34048 12406 34060
rect 17681 34051 17739 34057
rect 17681 34048 17693 34051
rect 12400 34020 17693 34048
rect 12400 34008 12406 34020
rect 17681 34017 17693 34020
rect 17727 34017 17739 34051
rect 17681 34011 17739 34017
rect 17770 34008 17776 34060
rect 17828 34048 17834 34060
rect 21634 34048 21640 34060
rect 17828 34020 21640 34048
rect 17828 34008 17834 34020
rect 21634 34008 21640 34020
rect 21692 34008 21698 34060
rect 17218 33980 17224 33992
rect 17179 33952 17224 33980
rect 17218 33940 17224 33952
rect 17276 33940 17282 33992
rect 17405 33983 17463 33989
rect 17405 33949 17417 33983
rect 17451 33980 17463 33983
rect 17862 33980 17868 33992
rect 17451 33952 17868 33980
rect 17451 33949 17463 33952
rect 17405 33943 17463 33949
rect 17862 33940 17868 33952
rect 17920 33940 17926 33992
rect 19334 33940 19340 33992
rect 19392 33980 19398 33992
rect 20165 33983 20223 33989
rect 20165 33980 20177 33983
rect 19392 33952 20177 33980
rect 19392 33940 19398 33952
rect 20165 33949 20177 33952
rect 20211 33949 20223 33983
rect 20165 33943 20223 33949
rect 20254 33940 20260 33992
rect 20312 33980 20318 33992
rect 20533 33983 20591 33989
rect 20533 33980 20545 33983
rect 20312 33952 20545 33980
rect 20312 33940 20318 33952
rect 20533 33949 20545 33952
rect 20579 33949 20591 33983
rect 20533 33943 20591 33949
rect 1670 33912 1676 33924
rect 1631 33884 1676 33912
rect 1670 33872 1676 33884
rect 1728 33872 1734 33924
rect 17310 33912 17316 33924
rect 17271 33884 17316 33912
rect 17310 33872 17316 33884
rect 17368 33872 17374 33924
rect 17543 33915 17601 33921
rect 17543 33881 17555 33915
rect 17589 33912 17601 33915
rect 17954 33912 17960 33924
rect 17589 33884 17960 33912
rect 17589 33881 17601 33884
rect 17543 33875 17601 33881
rect 17954 33872 17960 33884
rect 18012 33872 18018 33924
rect 19352 33884 20300 33912
rect 19352 33856 19380 33884
rect 17037 33847 17095 33853
rect 17037 33813 17049 33847
rect 17083 33844 17095 33847
rect 18966 33844 18972 33856
rect 17083 33816 18972 33844
rect 17083 33813 17095 33816
rect 17037 33807 17095 33813
rect 18966 33804 18972 33816
rect 19024 33804 19030 33856
rect 19334 33804 19340 33856
rect 19392 33804 19398 33856
rect 20070 33844 20076 33856
rect 20031 33816 20076 33844
rect 20070 33804 20076 33816
rect 20128 33804 20134 33856
rect 20272 33853 20300 33884
rect 20257 33847 20315 33853
rect 20257 33813 20269 33847
rect 20303 33813 20315 33847
rect 20257 33807 20315 33813
rect 20346 33804 20352 33856
rect 20404 33844 20410 33856
rect 21928 33844 21956 34088
rect 22281 33983 22339 33989
rect 22281 33949 22293 33983
rect 22327 33949 22339 33983
rect 22281 33943 22339 33949
rect 22373 33983 22431 33989
rect 22373 33949 22385 33983
rect 22419 33980 22431 33983
rect 22922 33980 22928 33992
rect 22419 33952 22928 33980
rect 22419 33949 22431 33952
rect 22373 33943 22431 33949
rect 22296 33912 22324 33943
rect 22922 33940 22928 33952
rect 22980 33940 22986 33992
rect 23124 33989 23152 34088
rect 25038 34076 25044 34128
rect 25096 34116 25102 34128
rect 25774 34116 25780 34128
rect 25096 34088 25780 34116
rect 25096 34076 25102 34088
rect 25774 34076 25780 34088
rect 25832 34076 25838 34128
rect 40328 34088 41000 34116
rect 24762 34008 24768 34060
rect 24820 34048 24826 34060
rect 24820 34020 31754 34048
rect 24820 34008 24826 34020
rect 23109 33983 23167 33989
rect 23109 33949 23121 33983
rect 23155 33949 23167 33983
rect 23109 33943 23167 33949
rect 24581 33983 24639 33989
rect 24581 33949 24593 33983
rect 24627 33949 24639 33983
rect 24581 33943 24639 33949
rect 22830 33912 22836 33924
rect 22296 33884 22836 33912
rect 22830 33872 22836 33884
rect 22888 33872 22894 33924
rect 22940 33912 22968 33940
rect 23477 33915 23535 33921
rect 23477 33912 23489 33915
rect 22940 33884 23489 33912
rect 23477 33881 23489 33884
rect 23523 33881 23535 33915
rect 24596 33912 24624 33943
rect 24670 33940 24676 33992
rect 24728 33980 24734 33992
rect 24728 33952 24773 33980
rect 24728 33940 24734 33952
rect 24854 33940 24860 33992
rect 24912 33980 24918 33992
rect 25087 33983 25145 33989
rect 24912 33952 24957 33980
rect 24912 33940 24918 33952
rect 25087 33949 25099 33983
rect 25133 33980 25145 33983
rect 25406 33980 25412 33992
rect 25133 33952 25412 33980
rect 25133 33949 25145 33952
rect 25087 33943 25145 33949
rect 25406 33940 25412 33952
rect 25464 33980 25470 33992
rect 26050 33980 26056 33992
rect 25464 33952 26056 33980
rect 25464 33940 25470 33952
rect 26050 33940 26056 33952
rect 26108 33940 26114 33992
rect 23477 33875 23535 33881
rect 23768 33884 24624 33912
rect 24949 33915 25007 33921
rect 23768 33844 23796 33884
rect 24949 33881 24961 33915
rect 24995 33881 25007 33915
rect 24949 33875 25007 33881
rect 20404 33816 20449 33844
rect 21928 33816 23796 33844
rect 20404 33804 20410 33816
rect 23934 33804 23940 33856
rect 23992 33844 23998 33856
rect 24964 33844 24992 33875
rect 25222 33844 25228 33856
rect 23992 33816 24992 33844
rect 25183 33816 25228 33844
rect 23992 33804 23998 33816
rect 25222 33804 25228 33816
rect 25280 33804 25286 33856
rect 31726 33844 31754 34020
rect 40034 33940 40040 33992
rect 40092 33980 40098 33992
rect 40328 33989 40356 34088
rect 40420 34020 40908 34048
rect 40420 33989 40448 34020
rect 40129 33983 40187 33989
rect 40129 33980 40141 33983
rect 40092 33952 40141 33980
rect 40092 33940 40098 33952
rect 40129 33949 40141 33952
rect 40175 33949 40187 33983
rect 40129 33943 40187 33949
rect 40277 33983 40356 33989
rect 40277 33949 40289 33983
rect 40323 33952 40356 33983
rect 40405 33983 40463 33989
rect 40323 33949 40335 33952
rect 40277 33943 40335 33949
rect 40405 33949 40417 33983
rect 40451 33949 40463 33983
rect 40405 33943 40463 33949
rect 40586 33940 40592 33992
rect 40644 33989 40650 33992
rect 40644 33980 40652 33989
rect 40644 33952 40689 33980
rect 40644 33943 40652 33952
rect 40644 33940 40650 33943
rect 40494 33872 40500 33924
rect 40552 33912 40558 33924
rect 40552 33884 40597 33912
rect 40552 33872 40558 33884
rect 40773 33847 40831 33853
rect 40773 33844 40785 33847
rect 31726 33816 40785 33844
rect 40773 33813 40785 33816
rect 40819 33813 40831 33847
rect 40880 33844 40908 34020
rect 40972 33912 41000 34088
rect 41340 33989 41368 34156
rect 41325 33983 41383 33989
rect 41325 33949 41337 33983
rect 41371 33949 41383 33983
rect 57974 33980 57980 33992
rect 57935 33952 57980 33980
rect 41325 33943 41383 33949
rect 57974 33940 57980 33952
rect 58032 33940 58038 33992
rect 50982 33912 50988 33924
rect 40972 33884 50988 33912
rect 50982 33872 50988 33884
rect 51040 33872 51046 33924
rect 58345 33915 58403 33921
rect 58345 33881 58357 33915
rect 58391 33912 58403 33915
rect 58986 33912 58992 33924
rect 58391 33884 58992 33912
rect 58391 33881 58403 33884
rect 58345 33875 58403 33881
rect 58986 33872 58992 33884
rect 59044 33872 59050 33924
rect 41509 33847 41567 33853
rect 41509 33844 41521 33847
rect 40880 33816 41521 33844
rect 40773 33807 40831 33813
rect 41509 33813 41521 33816
rect 41555 33844 41567 33847
rect 44082 33844 44088 33856
rect 41555 33816 44088 33844
rect 41555 33813 41567 33816
rect 41509 33807 41567 33813
rect 44082 33804 44088 33816
rect 44140 33804 44146 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 19058 33600 19064 33652
rect 19116 33640 19122 33652
rect 20257 33643 20315 33649
rect 20257 33640 20269 33643
rect 19116 33612 20269 33640
rect 19116 33600 19122 33612
rect 20257 33609 20269 33612
rect 20303 33609 20315 33643
rect 20257 33603 20315 33609
rect 20349 33643 20407 33649
rect 20349 33609 20361 33643
rect 20395 33640 20407 33643
rect 20530 33640 20536 33652
rect 20395 33612 20536 33640
rect 20395 33609 20407 33612
rect 20349 33603 20407 33609
rect 20530 33600 20536 33612
rect 20588 33600 20594 33652
rect 32858 33640 32864 33652
rect 21100 33612 32864 33640
rect 1857 33575 1915 33581
rect 1857 33541 1869 33575
rect 1903 33572 1915 33575
rect 1946 33572 1952 33584
rect 1903 33544 1952 33572
rect 1903 33541 1915 33544
rect 1857 33535 1915 33541
rect 1946 33532 1952 33544
rect 2004 33532 2010 33584
rect 20070 33532 20076 33584
rect 20128 33572 20134 33584
rect 21100 33572 21128 33612
rect 32858 33600 32864 33612
rect 32916 33600 32922 33652
rect 35342 33640 35348 33652
rect 32968 33612 35348 33640
rect 20128 33544 21128 33572
rect 20128 33532 20134 33544
rect 21174 33532 21180 33584
rect 21232 33572 21238 33584
rect 25314 33572 25320 33584
rect 21232 33544 25084 33572
rect 25275 33544 25320 33572
rect 21232 33532 21238 33544
rect 1670 33504 1676 33516
rect 1631 33476 1676 33504
rect 1670 33464 1676 33476
rect 1728 33464 1734 33516
rect 17773 33507 17831 33513
rect 17773 33473 17785 33507
rect 17819 33504 17831 33507
rect 18874 33504 18880 33516
rect 17819 33476 18880 33504
rect 17819 33473 17831 33476
rect 17773 33467 17831 33473
rect 18874 33464 18880 33476
rect 18932 33464 18938 33516
rect 19426 33464 19432 33516
rect 19484 33504 19490 33516
rect 20165 33507 20223 33513
rect 20165 33504 20177 33507
rect 19484 33476 20177 33504
rect 19484 33464 19490 33476
rect 20165 33473 20177 33476
rect 20211 33473 20223 33507
rect 20165 33467 20223 33473
rect 20254 33464 20260 33516
rect 20312 33504 20318 33516
rect 20533 33507 20591 33513
rect 20533 33504 20545 33507
rect 20312 33476 20545 33504
rect 20312 33464 20318 33476
rect 20533 33473 20545 33476
rect 20579 33473 20591 33507
rect 23566 33504 23572 33516
rect 23527 33476 23572 33504
rect 20533 33467 20591 33473
rect 23566 33464 23572 33476
rect 23624 33464 23630 33516
rect 25056 33513 25084 33544
rect 25314 33532 25320 33544
rect 25372 33572 25378 33584
rect 32968 33572 32996 33612
rect 35342 33600 35348 33612
rect 35400 33600 35406 33652
rect 25372 33544 32996 33572
rect 25372 33532 25378 33544
rect 25041 33507 25099 33513
rect 25041 33473 25053 33507
rect 25087 33473 25099 33507
rect 25041 33467 25099 33473
rect 25189 33507 25247 33513
rect 25189 33473 25201 33507
rect 25235 33504 25247 33507
rect 25235 33476 25360 33504
rect 25235 33473 25247 33476
rect 25189 33467 25247 33473
rect 17954 33436 17960 33448
rect 17915 33408 17960 33436
rect 17954 33396 17960 33408
rect 18012 33396 18018 33448
rect 23658 33396 23664 33448
rect 23716 33436 23722 33448
rect 23934 33436 23940 33448
rect 23716 33408 23940 33436
rect 23716 33396 23722 33408
rect 23934 33396 23940 33408
rect 23992 33396 23998 33448
rect 25332 33436 25360 33476
rect 25406 33464 25412 33516
rect 25464 33504 25470 33516
rect 25547 33507 25605 33513
rect 25464 33476 25509 33504
rect 25464 33464 25470 33476
rect 25547 33473 25559 33507
rect 25593 33504 25605 33507
rect 25774 33504 25780 33516
rect 25593 33476 25780 33504
rect 25593 33473 25605 33476
rect 25547 33467 25605 33473
rect 25774 33464 25780 33476
rect 25832 33464 25838 33516
rect 27338 33504 27344 33516
rect 27299 33476 27344 33504
rect 27338 33464 27344 33476
rect 27396 33464 27402 33516
rect 27522 33504 27528 33516
rect 27483 33476 27528 33504
rect 27522 33464 27528 33476
rect 27580 33464 27586 33516
rect 27614 33464 27620 33516
rect 27672 33504 27678 33516
rect 27893 33507 27951 33513
rect 27893 33504 27905 33507
rect 27672 33476 27905 33504
rect 27672 33464 27678 33476
rect 27893 33473 27905 33476
rect 27939 33473 27951 33507
rect 28442 33504 28448 33516
rect 28403 33476 28448 33504
rect 27893 33467 27951 33473
rect 28442 33464 28448 33476
rect 28500 33464 28506 33516
rect 29181 33507 29239 33513
rect 29181 33473 29193 33507
rect 29227 33504 29239 33507
rect 32122 33504 32128 33516
rect 29227 33476 32128 33504
rect 29227 33473 29239 33476
rect 29181 33467 29239 33473
rect 32122 33464 32128 33476
rect 32180 33464 32186 33516
rect 32766 33504 32772 33516
rect 32727 33476 32772 33504
rect 32766 33464 32772 33476
rect 32824 33464 32830 33516
rect 32950 33504 32956 33516
rect 32911 33476 32956 33504
rect 32950 33464 32956 33476
rect 33008 33464 33014 33516
rect 33042 33464 33048 33516
rect 33100 33513 33106 33516
rect 33100 33504 33111 33513
rect 33183 33507 33241 33513
rect 33100 33476 33145 33504
rect 33100 33467 33111 33476
rect 33183 33473 33195 33507
rect 33229 33504 33241 33507
rect 34054 33504 34060 33516
rect 33229 33476 34060 33504
rect 33229 33473 33241 33476
rect 33183 33467 33241 33473
rect 33100 33464 33106 33467
rect 34054 33464 34060 33476
rect 34112 33504 34118 33516
rect 36078 33504 36084 33516
rect 34112 33476 36084 33504
rect 34112 33464 34118 33476
rect 36078 33464 36084 33476
rect 36136 33504 36142 33516
rect 40586 33504 40592 33516
rect 36136 33476 40592 33504
rect 36136 33464 36142 33476
rect 40586 33464 40592 33476
rect 40644 33464 40650 33516
rect 26602 33436 26608 33448
rect 25332 33408 26608 33436
rect 26602 33396 26608 33408
rect 26660 33396 26666 33448
rect 28460 33436 28488 33464
rect 29457 33439 29515 33445
rect 29457 33436 29469 33439
rect 28460 33408 29469 33436
rect 29457 33405 29469 33408
rect 29503 33405 29515 33439
rect 29457 33399 29515 33405
rect 19981 33371 20039 33377
rect 19981 33337 19993 33371
rect 20027 33368 20039 33371
rect 32766 33368 32772 33380
rect 20027 33340 32772 33368
rect 20027 33337 20039 33340
rect 19981 33331 20039 33337
rect 32766 33328 32772 33340
rect 32824 33328 32830 33380
rect 32858 33328 32864 33380
rect 32916 33368 32922 33380
rect 34698 33368 34704 33380
rect 32916 33340 34704 33368
rect 32916 33328 32922 33340
rect 34698 33328 34704 33340
rect 34756 33328 34762 33380
rect 17310 33260 17316 33312
rect 17368 33300 17374 33312
rect 17954 33300 17960 33312
rect 17368 33272 17960 33300
rect 17368 33260 17374 33272
rect 17954 33260 17960 33272
rect 18012 33260 18018 33312
rect 19426 33260 19432 33312
rect 19484 33300 19490 33312
rect 20346 33300 20352 33312
rect 19484 33272 20352 33300
rect 19484 33260 19490 33272
rect 20346 33260 20352 33272
rect 20404 33260 20410 33312
rect 25682 33300 25688 33312
rect 25643 33272 25688 33300
rect 25682 33260 25688 33272
rect 25740 33260 25746 33312
rect 28629 33303 28687 33309
rect 28629 33269 28641 33303
rect 28675 33300 28687 33303
rect 29546 33300 29552 33312
rect 28675 33272 29552 33300
rect 28675 33269 28687 33272
rect 28629 33263 28687 33269
rect 29546 33260 29552 33272
rect 29604 33260 29610 33312
rect 33321 33303 33379 33309
rect 33321 33269 33333 33303
rect 33367 33300 33379 33303
rect 33410 33300 33416 33312
rect 33367 33272 33416 33300
rect 33367 33269 33379 33272
rect 33321 33263 33379 33269
rect 33410 33260 33416 33272
rect 33468 33260 33474 33312
rect 46934 33260 46940 33312
rect 46992 33300 46998 33312
rect 48958 33300 48964 33312
rect 46992 33272 48964 33300
rect 46992 33260 46998 33272
rect 48958 33260 48964 33272
rect 49016 33260 49022 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 16761 33099 16819 33105
rect 16761 33065 16773 33099
rect 16807 33065 16819 33099
rect 16761 33059 16819 33065
rect 16945 33099 17003 33105
rect 16945 33065 16957 33099
rect 16991 33096 17003 33099
rect 17218 33096 17224 33108
rect 16991 33068 17224 33096
rect 16991 33065 17003 33068
rect 16945 33059 17003 33065
rect 16776 33028 16804 33059
rect 17218 33056 17224 33068
rect 17276 33056 17282 33108
rect 17310 33056 17316 33108
rect 17368 33096 17374 33108
rect 22373 33099 22431 33105
rect 17368 33068 22324 33096
rect 17368 33056 17374 33068
rect 19610 33028 19616 33040
rect 16776 33000 19616 33028
rect 19610 32988 19616 33000
rect 19668 32988 19674 33040
rect 19720 33000 20025 33028
rect 14458 32920 14464 32972
rect 14516 32960 14522 32972
rect 17218 32960 17224 32972
rect 14516 32932 17224 32960
rect 14516 32920 14522 32932
rect 17218 32920 17224 32932
rect 17276 32920 17282 32972
rect 18966 32920 18972 32972
rect 19024 32960 19030 32972
rect 19720 32960 19748 33000
rect 19024 32932 19748 32960
rect 19997 32960 20025 33000
rect 19997 32932 20760 32960
rect 19024 32920 19030 32932
rect 8938 32852 8944 32904
rect 8996 32892 9002 32904
rect 16577 32895 16635 32901
rect 16577 32892 16589 32895
rect 8996 32864 16589 32892
rect 8996 32852 9002 32864
rect 16577 32861 16589 32864
rect 16623 32861 16635 32895
rect 16577 32855 16635 32861
rect 16761 32895 16819 32901
rect 16761 32861 16773 32895
rect 16807 32892 16819 32895
rect 17589 32895 17647 32901
rect 17589 32892 17601 32895
rect 16807 32864 17601 32892
rect 16807 32861 16819 32864
rect 16761 32855 16819 32861
rect 17589 32861 17601 32864
rect 17635 32861 17647 32895
rect 17862 32892 17868 32904
rect 17823 32864 17868 32892
rect 17589 32855 17647 32861
rect 17604 32824 17632 32855
rect 17862 32852 17868 32864
rect 17920 32852 17926 32904
rect 17954 32852 17960 32904
rect 18012 32892 18018 32904
rect 18012 32864 18057 32892
rect 18012 32852 18018 32864
rect 18322 32852 18328 32904
rect 18380 32892 18386 32904
rect 18417 32895 18475 32901
rect 18417 32892 18429 32895
rect 18380 32864 18429 32892
rect 18380 32852 18386 32864
rect 18417 32861 18429 32864
rect 18463 32861 18475 32895
rect 18417 32855 18475 32861
rect 18782 32852 18788 32904
rect 18840 32892 18846 32904
rect 19334 32892 19340 32904
rect 18840 32864 19340 32892
rect 18840 32852 18846 32864
rect 19334 32852 19340 32864
rect 19392 32892 19398 32904
rect 19613 32895 19671 32901
rect 19613 32892 19625 32895
rect 19392 32864 19625 32892
rect 19392 32852 19398 32864
rect 19613 32861 19625 32864
rect 19659 32861 19671 32895
rect 19779 32895 19837 32901
rect 19779 32892 19791 32895
rect 19613 32855 19671 32861
rect 19720 32864 19791 32892
rect 19518 32824 19524 32836
rect 17604 32796 19524 32824
rect 19518 32784 19524 32796
rect 19576 32784 19582 32836
rect 17218 32716 17224 32768
rect 17276 32756 17282 32768
rect 17497 32759 17555 32765
rect 17497 32756 17509 32759
rect 17276 32728 17509 32756
rect 17276 32716 17282 32728
rect 17497 32725 17509 32728
rect 17543 32725 17555 32759
rect 17497 32719 17555 32725
rect 18046 32716 18052 32768
rect 18104 32756 18110 32768
rect 19334 32756 19340 32768
rect 18104 32728 19340 32756
rect 18104 32716 18110 32728
rect 19334 32716 19340 32728
rect 19392 32716 19398 32768
rect 19426 32716 19432 32768
rect 19484 32756 19490 32768
rect 19720 32756 19748 32864
rect 19779 32861 19791 32864
rect 19825 32861 19837 32895
rect 19982 32895 20040 32901
rect 19779 32855 19837 32861
rect 19890 32873 19948 32879
rect 19890 32839 19902 32873
rect 19936 32839 19948 32873
rect 19982 32861 19994 32895
rect 20028 32894 20040 32895
rect 20070 32894 20076 32904
rect 20028 32866 20076 32894
rect 20028 32861 20040 32866
rect 19982 32855 20040 32861
rect 20070 32852 20076 32866
rect 20128 32852 20134 32904
rect 20254 32852 20260 32904
rect 20312 32892 20318 32904
rect 20732 32892 20760 32932
rect 20806 32920 20812 32972
rect 20864 32960 20870 32972
rect 22296 32960 22324 33068
rect 22373 33065 22385 33099
rect 22419 33096 22431 33099
rect 33502 33096 33508 33108
rect 22419 33068 33508 33096
rect 22419 33065 22431 33068
rect 22373 33059 22431 33065
rect 33502 33056 33508 33068
rect 33560 33056 33566 33108
rect 34054 33096 34060 33108
rect 34015 33068 34060 33096
rect 34054 33056 34060 33068
rect 34112 33056 34118 33108
rect 26145 33031 26203 33037
rect 26145 32997 26157 33031
rect 26191 33028 26203 33031
rect 26789 33031 26847 33037
rect 26789 33028 26801 33031
rect 26191 33000 26801 33028
rect 26191 32997 26203 33000
rect 26145 32991 26203 32997
rect 26789 32997 26801 33000
rect 26835 33028 26847 33031
rect 27522 33028 27528 33040
rect 26835 33000 27528 33028
rect 26835 32997 26847 33000
rect 26789 32991 26847 32997
rect 27522 32988 27528 33000
rect 27580 32988 27586 33040
rect 32766 32988 32772 33040
rect 32824 33028 32830 33040
rect 43990 33028 43996 33040
rect 32824 33000 43996 33028
rect 32824 32988 32830 33000
rect 43990 32988 43996 33000
rect 44048 32988 44054 33040
rect 58158 32960 58164 32972
rect 20864 32932 21588 32960
rect 22296 32932 33180 32960
rect 58119 32932 58164 32960
rect 20864 32920 20870 32932
rect 21560 32904 21588 32932
rect 20993 32895 21051 32901
rect 20993 32892 21005 32895
rect 20312 32864 20668 32892
rect 20732 32864 21005 32892
rect 20312 32852 20318 32864
rect 19890 32836 19948 32839
rect 19886 32784 19892 32836
rect 19944 32784 19950 32836
rect 20640 32824 20668 32864
rect 20993 32861 21005 32864
rect 21039 32861 21051 32895
rect 21174 32892 21180 32904
rect 21135 32864 21180 32892
rect 20993 32855 21051 32861
rect 21174 32852 21180 32864
rect 21232 32852 21238 32904
rect 21542 32892 21548 32904
rect 21503 32864 21548 32892
rect 21542 32852 21548 32864
rect 21600 32852 21606 32904
rect 21726 32892 21732 32904
rect 21687 32864 21732 32892
rect 21726 32852 21732 32864
rect 21784 32852 21790 32904
rect 21910 32892 21916 32904
rect 21871 32864 21916 32892
rect 21910 32852 21916 32864
rect 21968 32852 21974 32904
rect 23566 32852 23572 32904
rect 23624 32892 23630 32904
rect 25498 32892 25504 32904
rect 23624 32864 25504 32892
rect 23624 32852 23630 32864
rect 25498 32852 25504 32864
rect 25556 32852 25562 32904
rect 25590 32852 25596 32904
rect 25648 32892 25654 32904
rect 25648 32864 25693 32892
rect 25648 32852 25654 32864
rect 25958 32852 25964 32904
rect 26016 32901 26022 32904
rect 26016 32892 26024 32901
rect 26016 32864 26061 32892
rect 26016 32855 26024 32864
rect 26016 32852 26022 32855
rect 26142 32852 26148 32904
rect 26200 32852 26206 32904
rect 26697 32895 26755 32901
rect 26697 32861 26709 32895
rect 26743 32861 26755 32895
rect 26697 32855 26755 32861
rect 26973 32895 27031 32901
rect 26973 32861 26985 32895
rect 27019 32892 27031 32895
rect 27338 32892 27344 32904
rect 27019 32864 27344 32892
rect 27019 32861 27031 32864
rect 26973 32855 27031 32861
rect 20806 32824 20812 32836
rect 20640 32796 20812 32824
rect 20806 32784 20812 32796
rect 20864 32784 20870 32836
rect 21358 32784 21364 32836
rect 21416 32824 21422 32836
rect 25777 32827 25835 32833
rect 25777 32824 25789 32827
rect 21416 32796 25789 32824
rect 21416 32784 21422 32796
rect 25777 32793 25789 32796
rect 25823 32793 25835 32827
rect 25777 32787 25835 32793
rect 25869 32827 25927 32833
rect 25869 32793 25881 32827
rect 25915 32824 25927 32827
rect 26160 32824 26188 32852
rect 25915 32796 26188 32824
rect 26712 32824 26740 32855
rect 27338 32852 27344 32864
rect 27396 32852 27402 32904
rect 27433 32895 27491 32901
rect 27433 32861 27445 32895
rect 27479 32892 27491 32895
rect 27522 32892 27528 32904
rect 27479 32864 27528 32892
rect 27479 32861 27491 32864
rect 27433 32855 27491 32861
rect 27522 32852 27528 32864
rect 27580 32852 27586 32904
rect 33042 32892 33048 32904
rect 33003 32864 33048 32892
rect 33042 32852 33048 32864
rect 33100 32852 33106 32904
rect 33152 32901 33180 32932
rect 58158 32920 58164 32932
rect 58216 32920 58222 32972
rect 33137 32895 33195 32901
rect 33137 32861 33149 32895
rect 33183 32861 33195 32895
rect 33137 32855 33195 32861
rect 33321 32895 33379 32901
rect 33321 32861 33333 32895
rect 33367 32861 33379 32895
rect 33321 32855 33379 32861
rect 27614 32824 27620 32836
rect 26712 32796 27620 32824
rect 25915 32793 25927 32796
rect 25869 32787 25927 32793
rect 27614 32784 27620 32796
rect 27672 32784 27678 32836
rect 33336 32824 33364 32855
rect 33410 32852 33416 32904
rect 33468 32892 33474 32904
rect 42886 32892 42892 32904
rect 33468 32864 33513 32892
rect 42847 32864 42892 32892
rect 33468 32852 33474 32864
rect 42886 32852 42892 32864
rect 42944 32852 42950 32904
rect 43070 32901 43076 32904
rect 43037 32895 43076 32901
rect 43037 32861 43049 32895
rect 43037 32855 43076 32861
rect 43070 32852 43076 32855
rect 43128 32852 43134 32904
rect 43346 32852 43352 32904
rect 43404 32901 43410 32904
rect 43404 32892 43412 32901
rect 43404 32864 43449 32892
rect 43404 32855 43412 32864
rect 43404 32852 43410 32855
rect 57514 32852 57520 32904
rect 57572 32892 57578 32904
rect 57885 32895 57943 32901
rect 57885 32892 57897 32895
rect 57572 32864 57897 32892
rect 57572 32852 57578 32864
rect 57885 32861 57897 32864
rect 57931 32861 57943 32895
rect 57885 32855 57943 32861
rect 33962 32824 33968 32836
rect 31726 32796 33364 32824
rect 33923 32796 33968 32824
rect 19484 32728 19748 32756
rect 19484 32716 19490 32728
rect 25498 32716 25504 32768
rect 25556 32756 25562 32768
rect 31726 32756 31754 32796
rect 33962 32784 33968 32796
rect 34020 32784 34026 32836
rect 35342 32784 35348 32836
rect 35400 32824 35406 32836
rect 43165 32827 43223 32833
rect 43165 32824 43177 32827
rect 35400 32796 43177 32824
rect 35400 32784 35406 32796
rect 43165 32793 43177 32796
rect 43211 32793 43223 32827
rect 43165 32787 43223 32793
rect 43257 32827 43315 32833
rect 43257 32793 43269 32827
rect 43303 32824 43315 32827
rect 44266 32824 44272 32836
rect 43303 32796 44272 32824
rect 43303 32793 43315 32796
rect 43257 32787 43315 32793
rect 44266 32784 44272 32796
rect 44324 32784 44330 32836
rect 57054 32824 57060 32836
rect 57015 32796 57060 32824
rect 57054 32784 57060 32796
rect 57112 32784 57118 32836
rect 25556 32728 31754 32756
rect 32861 32759 32919 32765
rect 25556 32716 25562 32728
rect 32861 32725 32873 32759
rect 32907 32756 32919 32759
rect 33778 32756 33784 32768
rect 32907 32728 33784 32756
rect 32907 32725 32919 32728
rect 32861 32719 32919 32725
rect 33778 32716 33784 32728
rect 33836 32716 33842 32768
rect 36538 32716 36544 32768
rect 36596 32756 36602 32768
rect 43533 32759 43591 32765
rect 43533 32756 43545 32759
rect 36596 32728 43545 32756
rect 36596 32716 36602 32728
rect 43533 32725 43545 32728
rect 43579 32725 43591 32759
rect 43533 32719 43591 32725
rect 48038 32716 48044 32768
rect 48096 32756 48102 32768
rect 57149 32759 57207 32765
rect 57149 32756 57161 32759
rect 48096 32728 57161 32756
rect 48096 32716 48102 32728
rect 57149 32725 57161 32728
rect 57195 32725 57207 32759
rect 57149 32719 57207 32725
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 17954 32512 17960 32564
rect 18012 32552 18018 32564
rect 18782 32552 18788 32564
rect 18012 32524 18788 32552
rect 18012 32512 18018 32524
rect 18782 32512 18788 32524
rect 18840 32512 18846 32564
rect 19334 32512 19340 32564
rect 19392 32552 19398 32564
rect 19978 32552 19984 32564
rect 19392 32524 19984 32552
rect 19392 32512 19398 32524
rect 19978 32512 19984 32524
rect 20036 32512 20042 32564
rect 36538 32552 36544 32564
rect 31726 32524 36544 32552
rect 1857 32487 1915 32493
rect 1857 32453 1869 32487
rect 1903 32484 1915 32487
rect 2314 32484 2320 32496
rect 1903 32456 2320 32484
rect 1903 32453 1915 32456
rect 1857 32447 1915 32453
rect 2314 32444 2320 32456
rect 2372 32444 2378 32496
rect 17862 32444 17868 32496
rect 17920 32484 17926 32496
rect 18233 32487 18291 32493
rect 18233 32484 18245 32487
rect 17920 32456 18245 32484
rect 17920 32444 17926 32456
rect 18233 32453 18245 32456
rect 18279 32484 18291 32487
rect 19426 32484 19432 32496
rect 18279 32456 19432 32484
rect 18279 32453 18291 32456
rect 18233 32447 18291 32453
rect 19426 32444 19432 32456
rect 19484 32484 19490 32496
rect 19797 32487 19855 32493
rect 19797 32484 19809 32487
rect 19484 32456 19809 32484
rect 19484 32444 19490 32456
rect 19797 32453 19809 32456
rect 19843 32453 19855 32487
rect 20441 32487 20499 32493
rect 20441 32484 20453 32487
rect 19797 32447 19855 32453
rect 19904 32456 20453 32484
rect 1670 32416 1676 32428
rect 1631 32388 1676 32416
rect 1670 32376 1676 32388
rect 1728 32376 1734 32428
rect 17402 32376 17408 32428
rect 17460 32416 17466 32428
rect 18693 32419 18751 32425
rect 18693 32416 18705 32419
rect 17460 32388 18705 32416
rect 17460 32376 17466 32388
rect 18693 32385 18705 32388
rect 18739 32385 18751 32419
rect 18693 32379 18751 32385
rect 18230 32308 18236 32360
rect 18288 32348 18294 32360
rect 18325 32351 18383 32357
rect 18325 32348 18337 32351
rect 18288 32320 18337 32348
rect 18288 32308 18294 32320
rect 18325 32317 18337 32320
rect 18371 32348 18383 32351
rect 18414 32348 18420 32360
rect 18371 32320 18420 32348
rect 18371 32317 18383 32320
rect 18325 32311 18383 32317
rect 18414 32308 18420 32320
rect 18472 32308 18478 32360
rect 18708 32280 18736 32379
rect 18782 32376 18788 32428
rect 18840 32416 18846 32428
rect 19904 32416 19932 32456
rect 20441 32453 20453 32456
rect 20487 32484 20499 32487
rect 20622 32484 20628 32496
rect 20487 32456 20628 32484
rect 20487 32453 20499 32456
rect 20441 32447 20499 32453
rect 20622 32444 20628 32456
rect 20680 32444 20686 32496
rect 25222 32444 25228 32496
rect 25280 32484 25286 32496
rect 25409 32487 25467 32493
rect 25409 32484 25421 32487
rect 25280 32456 25421 32484
rect 25280 32444 25286 32456
rect 25409 32453 25421 32456
rect 25455 32453 25467 32487
rect 25409 32447 25467 32453
rect 25961 32487 26019 32493
rect 25961 32453 25973 32487
rect 26007 32484 26019 32487
rect 27338 32484 27344 32496
rect 26007 32456 27344 32484
rect 26007 32453 26019 32456
rect 25961 32447 26019 32453
rect 27338 32444 27344 32456
rect 27396 32444 27402 32496
rect 18840 32388 19932 32416
rect 18840 32376 18846 32388
rect 19978 32376 19984 32428
rect 20036 32416 20042 32428
rect 20254 32416 20260 32428
rect 20036 32388 20260 32416
rect 20036 32376 20042 32388
rect 20254 32376 20260 32388
rect 20312 32376 20318 32428
rect 20349 32419 20407 32425
rect 20349 32385 20361 32419
rect 20395 32385 20407 32419
rect 22186 32416 22192 32428
rect 22147 32388 22192 32416
rect 20349 32379 20407 32385
rect 19242 32348 19248 32360
rect 19203 32320 19248 32348
rect 19242 32308 19248 32320
rect 19300 32308 19306 32360
rect 19886 32348 19892 32360
rect 19847 32320 19892 32348
rect 19886 32308 19892 32320
rect 19944 32308 19950 32360
rect 19426 32280 19432 32292
rect 18708 32252 19432 32280
rect 19426 32240 19432 32252
rect 19484 32280 19490 32292
rect 20364 32280 20392 32379
rect 22186 32376 22192 32388
rect 22244 32376 22250 32428
rect 22281 32419 22339 32425
rect 22281 32385 22293 32419
rect 22327 32385 22339 32419
rect 22281 32379 22339 32385
rect 22373 32419 22431 32425
rect 22373 32385 22385 32419
rect 22419 32385 22431 32419
rect 22554 32416 22560 32428
rect 22515 32388 22560 32416
rect 22373 32379 22431 32385
rect 22296 32348 22324 32379
rect 19484 32252 20392 32280
rect 20456 32320 22324 32348
rect 19484 32240 19490 32252
rect 19058 32172 19064 32224
rect 19116 32212 19122 32224
rect 20456 32212 20484 32320
rect 20530 32240 20536 32292
rect 20588 32280 20594 32292
rect 22388 32280 22416 32379
rect 22554 32376 22560 32388
rect 22612 32376 22618 32428
rect 22649 32419 22707 32425
rect 22649 32385 22661 32419
rect 22695 32385 22707 32419
rect 22649 32379 22707 32385
rect 25593 32419 25651 32425
rect 25593 32385 25605 32419
rect 25639 32416 25651 32419
rect 31726 32416 31754 32524
rect 36538 32512 36544 32524
rect 36596 32512 36602 32564
rect 42794 32552 42800 32564
rect 41386 32524 42800 32552
rect 41386 32484 41414 32524
rect 42794 32512 42800 32524
rect 42852 32512 42858 32564
rect 33060 32456 41414 32484
rect 33060 32425 33088 32456
rect 44082 32444 44088 32496
rect 44140 32484 44146 32496
rect 44913 32487 44971 32493
rect 44913 32484 44925 32487
rect 44140 32456 44925 32484
rect 44140 32444 44146 32456
rect 44913 32453 44925 32456
rect 44959 32453 44971 32487
rect 44913 32447 44971 32453
rect 45005 32487 45063 32493
rect 45005 32453 45017 32487
rect 45051 32484 45063 32487
rect 46106 32484 46112 32496
rect 45051 32456 46112 32484
rect 45051 32453 45063 32456
rect 45005 32447 45063 32453
rect 46106 32444 46112 32456
rect 46164 32444 46170 32496
rect 25639 32388 31754 32416
rect 33045 32419 33103 32425
rect 25639 32385 25651 32388
rect 25593 32379 25651 32385
rect 33045 32385 33057 32419
rect 33091 32385 33103 32419
rect 33502 32416 33508 32428
rect 33463 32388 33508 32416
rect 33045 32379 33103 32385
rect 22664 32348 22692 32379
rect 33502 32376 33508 32388
rect 33560 32376 33566 32428
rect 33870 32376 33876 32428
rect 33928 32416 33934 32428
rect 44726 32416 44732 32428
rect 33928 32388 41414 32416
rect 44687 32388 44732 32416
rect 33928 32376 33934 32388
rect 33137 32351 33195 32357
rect 22664 32320 31754 32348
rect 20588 32252 22416 32280
rect 20588 32240 20594 32252
rect 23014 32240 23020 32292
rect 23072 32280 23078 32292
rect 25958 32280 25964 32292
rect 23072 32252 25964 32280
rect 23072 32240 23078 32252
rect 25958 32240 25964 32252
rect 26016 32240 26022 32292
rect 27154 32240 27160 32292
rect 27212 32280 27218 32292
rect 27522 32280 27528 32292
rect 27212 32252 27528 32280
rect 27212 32240 27218 32252
rect 27522 32240 27528 32252
rect 27580 32240 27586 32292
rect 19116 32184 20484 32212
rect 22005 32215 22063 32221
rect 19116 32172 19122 32184
rect 22005 32181 22017 32215
rect 22051 32212 22063 32215
rect 24762 32212 24768 32224
rect 22051 32184 24768 32212
rect 22051 32181 22063 32184
rect 22005 32175 22063 32181
rect 24762 32172 24768 32184
rect 24820 32172 24826 32224
rect 31726 32212 31754 32320
rect 33137 32317 33149 32351
rect 33183 32317 33195 32351
rect 34146 32348 34152 32360
rect 33810 32320 34152 32348
rect 33137 32311 33195 32317
rect 33152 32280 33180 32311
rect 34146 32308 34152 32320
rect 34204 32308 34210 32360
rect 41386 32348 41414 32388
rect 44726 32376 44732 32388
rect 44784 32376 44790 32428
rect 45102 32419 45160 32425
rect 45102 32416 45114 32419
rect 45020 32388 45114 32416
rect 43346 32348 43352 32360
rect 41386 32320 43352 32348
rect 43346 32308 43352 32320
rect 43404 32308 43410 32360
rect 44450 32308 44456 32360
rect 44508 32348 44514 32360
rect 45020 32348 45048 32388
rect 45102 32385 45114 32388
rect 45148 32385 45160 32419
rect 45102 32379 45160 32385
rect 45738 32348 45744 32360
rect 44508 32320 45744 32348
rect 44508 32308 44514 32320
rect 45738 32308 45744 32320
rect 45796 32308 45802 32360
rect 33502 32280 33508 32292
rect 33152 32252 33508 32280
rect 33502 32240 33508 32252
rect 33560 32240 33566 32292
rect 33873 32283 33931 32289
rect 33873 32249 33885 32283
rect 33919 32280 33931 32283
rect 36998 32280 37004 32292
rect 33919 32252 37004 32280
rect 33919 32249 33931 32252
rect 33873 32243 33931 32249
rect 36998 32240 37004 32252
rect 37056 32240 37062 32292
rect 42610 32240 42616 32292
rect 42668 32280 42674 32292
rect 49694 32280 49700 32292
rect 42668 32252 49700 32280
rect 42668 32240 42674 32252
rect 49694 32240 49700 32252
rect 49752 32240 49758 32292
rect 45281 32215 45339 32221
rect 45281 32212 45293 32215
rect 31726 32184 45293 32212
rect 45281 32181 45293 32184
rect 45327 32181 45339 32215
rect 45281 32175 45339 32181
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 17494 31968 17500 32020
rect 17552 32008 17558 32020
rect 19794 32008 19800 32020
rect 17552 31980 19800 32008
rect 17552 31968 17558 31980
rect 19794 31968 19800 31980
rect 19852 31968 19858 32020
rect 19886 31968 19892 32020
rect 19944 32008 19950 32020
rect 20438 32008 20444 32020
rect 19944 31980 20444 32008
rect 19944 31968 19950 31980
rect 20438 31968 20444 31980
rect 20496 31968 20502 32020
rect 20898 31968 20904 32020
rect 20956 32008 20962 32020
rect 23109 32011 23167 32017
rect 23109 32008 23121 32011
rect 20956 31980 23121 32008
rect 20956 31968 20962 31980
rect 23109 31977 23121 31980
rect 23155 31977 23167 32011
rect 23109 31971 23167 31977
rect 38654 31968 38660 32020
rect 38712 32008 38718 32020
rect 44637 32011 44695 32017
rect 44637 32008 44649 32011
rect 38712 31980 44649 32008
rect 38712 31968 38718 31980
rect 44637 31977 44649 31980
rect 44683 31977 44695 32011
rect 44637 31971 44695 31977
rect 16482 31900 16488 31952
rect 16540 31940 16546 31952
rect 21361 31943 21419 31949
rect 16540 31912 20116 31940
rect 16540 31900 16546 31912
rect 1857 31875 1915 31881
rect 1857 31841 1869 31875
rect 1903 31872 1915 31875
rect 16758 31872 16764 31884
rect 1903 31844 16764 31872
rect 1903 31841 1915 31844
rect 1857 31835 1915 31841
rect 16758 31832 16764 31844
rect 16816 31832 16822 31884
rect 17954 31872 17960 31884
rect 17788 31844 17960 31872
rect 1670 31804 1676 31816
rect 1631 31776 1676 31804
rect 1670 31764 1676 31776
rect 1728 31764 1734 31816
rect 17402 31804 17408 31816
rect 17363 31776 17408 31804
rect 17402 31764 17408 31776
rect 17460 31764 17466 31816
rect 17494 31696 17500 31748
rect 17552 31736 17558 31748
rect 17788 31736 17816 31844
rect 17954 31832 17960 31844
rect 18012 31872 18018 31884
rect 18012 31844 18092 31872
rect 18012 31832 18018 31844
rect 18064 31813 18092 31844
rect 19334 31832 19340 31884
rect 19392 31872 19398 31884
rect 20088 31872 20116 31912
rect 21361 31909 21373 31943
rect 21407 31940 21419 31943
rect 22646 31940 22652 31952
rect 21407 31912 22652 31940
rect 21407 31909 21419 31912
rect 21361 31903 21419 31909
rect 22646 31900 22652 31912
rect 22704 31900 22710 31952
rect 23569 31943 23627 31949
rect 23569 31909 23581 31943
rect 23615 31940 23627 31943
rect 25866 31940 25872 31952
rect 23615 31912 25872 31940
rect 23615 31909 23627 31912
rect 23569 31903 23627 31909
rect 25866 31900 25872 31912
rect 25924 31900 25930 31952
rect 33502 31900 33508 31952
rect 33560 31940 33566 31952
rect 36170 31940 36176 31952
rect 33560 31912 36176 31940
rect 33560 31900 33566 31912
rect 36170 31900 36176 31912
rect 36228 31940 36234 31952
rect 36228 31912 38654 31940
rect 36228 31900 36234 31912
rect 23014 31872 23020 31884
rect 19392 31844 19932 31872
rect 20088 31844 23020 31872
rect 19392 31832 19398 31844
rect 19904 31813 19932 31844
rect 23014 31832 23020 31844
rect 23072 31832 23078 31884
rect 23201 31875 23259 31881
rect 23201 31841 23213 31875
rect 23247 31872 23259 31875
rect 24394 31872 24400 31884
rect 23247 31844 24400 31872
rect 23247 31841 23259 31844
rect 23201 31835 23259 31841
rect 24394 31832 24400 31844
rect 24452 31832 24458 31884
rect 25240 31844 25820 31872
rect 17865 31807 17923 31813
rect 17865 31773 17877 31807
rect 17911 31804 17923 31807
rect 18049 31807 18107 31813
rect 17911 31776 18000 31804
rect 17911 31773 17923 31776
rect 17865 31767 17923 31773
rect 17552 31708 17816 31736
rect 17972 31736 18000 31776
rect 18049 31773 18061 31807
rect 18095 31773 18107 31807
rect 18049 31767 18107 31773
rect 18877 31807 18935 31813
rect 18877 31773 18889 31807
rect 18923 31804 18935 31807
rect 19889 31807 19947 31813
rect 18923 31776 19840 31804
rect 18923 31773 18935 31776
rect 18877 31767 18935 31773
rect 18138 31736 18144 31748
rect 17972 31708 18144 31736
rect 17552 31696 17558 31708
rect 18138 31696 18144 31708
rect 18196 31736 18202 31748
rect 18322 31736 18328 31748
rect 18196 31708 18328 31736
rect 18196 31696 18202 31708
rect 18322 31696 18328 31708
rect 18380 31736 18386 31748
rect 19242 31736 19248 31748
rect 18380 31708 19248 31736
rect 18380 31696 18386 31708
rect 19242 31696 19248 31708
rect 19300 31696 19306 31748
rect 19812 31736 19840 31776
rect 19889 31773 19901 31807
rect 19935 31773 19947 31807
rect 19889 31767 19947 31773
rect 20441 31807 20499 31813
rect 20441 31773 20453 31807
rect 20487 31804 20499 31807
rect 20714 31804 20720 31816
rect 20487 31776 20720 31804
rect 20487 31773 20499 31776
rect 20441 31767 20499 31773
rect 20714 31764 20720 31776
rect 20772 31764 20778 31816
rect 20806 31764 20812 31816
rect 20864 31804 20870 31816
rect 21545 31807 21603 31813
rect 21545 31804 21557 31807
rect 20864 31776 21557 31804
rect 20864 31764 20870 31776
rect 21545 31773 21557 31776
rect 21591 31773 21603 31807
rect 21910 31804 21916 31816
rect 21871 31776 21916 31804
rect 21545 31767 21603 31773
rect 20530 31736 20536 31748
rect 19812 31708 20536 31736
rect 20530 31696 20536 31708
rect 20588 31696 20594 31748
rect 21560 31736 21588 31767
rect 21910 31764 21916 31776
rect 21968 31764 21974 31816
rect 22005 31807 22063 31813
rect 22005 31773 22017 31807
rect 22051 31804 22063 31807
rect 22186 31804 22192 31816
rect 22051 31776 22192 31804
rect 22051 31773 22063 31776
rect 22005 31767 22063 31773
rect 22186 31764 22192 31776
rect 22244 31764 22250 31816
rect 23109 31807 23167 31813
rect 23109 31773 23121 31807
rect 23155 31804 23167 31807
rect 23155 31776 23244 31804
rect 23155 31773 23167 31776
rect 23109 31767 23167 31773
rect 22554 31736 22560 31748
rect 21560 31708 22560 31736
rect 22554 31696 22560 31708
rect 22612 31696 22618 31748
rect 23216 31736 23244 31776
rect 23290 31764 23296 31816
rect 23348 31804 23354 31816
rect 23385 31807 23443 31813
rect 23385 31804 23397 31807
rect 23348 31776 23397 31804
rect 23348 31764 23354 31776
rect 23385 31773 23397 31776
rect 23431 31773 23443 31807
rect 25133 31807 25191 31813
rect 25133 31804 25145 31807
rect 25043 31776 25145 31804
rect 23385 31767 23443 31773
rect 25133 31773 25145 31776
rect 25179 31804 25191 31807
rect 25240 31804 25268 31844
rect 25179 31776 25268 31804
rect 25792 31804 25820 31844
rect 25958 31832 25964 31884
rect 26016 31872 26022 31884
rect 33870 31872 33876 31884
rect 26016 31844 33876 31872
rect 26016 31832 26022 31844
rect 32876 31813 32904 31844
rect 33870 31832 33876 31844
rect 33928 31832 33934 31884
rect 38626 31872 38654 31912
rect 42334 31900 42340 31952
rect 42392 31940 42398 31952
rect 42889 31943 42947 31949
rect 42889 31940 42901 31943
rect 42392 31912 42901 31940
rect 42392 31900 42398 31912
rect 42889 31909 42901 31912
rect 42935 31909 42947 31943
rect 44450 31940 44456 31952
rect 42889 31903 42947 31909
rect 44284 31912 44456 31940
rect 44284 31872 44312 31912
rect 44450 31900 44456 31912
rect 44508 31900 44514 31952
rect 44726 31900 44732 31952
rect 44784 31940 44790 31952
rect 49234 31940 49240 31952
rect 44784 31912 49240 31940
rect 44784 31900 44790 31912
rect 49234 31900 49240 31912
rect 49292 31900 49298 31952
rect 38626 31844 44312 31872
rect 32861 31807 32919 31813
rect 25792 31776 32812 31804
rect 25179 31773 25191 31776
rect 25133 31767 25191 31773
rect 23566 31736 23572 31748
rect 23216 31708 23572 31736
rect 23566 31696 23572 31708
rect 23624 31696 23630 31748
rect 14366 31628 14372 31680
rect 14424 31668 14430 31680
rect 17313 31671 17371 31677
rect 17313 31668 17325 31671
rect 14424 31640 17325 31668
rect 14424 31628 14430 31640
rect 17313 31637 17325 31640
rect 17359 31668 17371 31671
rect 25148 31668 25176 31767
rect 25685 31739 25743 31745
rect 25685 31705 25697 31739
rect 25731 31736 25743 31739
rect 25774 31736 25780 31748
rect 25731 31708 25780 31736
rect 25731 31705 25743 31708
rect 25685 31699 25743 31705
rect 25774 31696 25780 31708
rect 25832 31696 25838 31748
rect 25958 31696 25964 31748
rect 26016 31736 26022 31748
rect 31754 31736 31760 31748
rect 26016 31708 31760 31736
rect 26016 31696 26022 31708
rect 31754 31696 31760 31708
rect 31812 31736 31818 31748
rect 32784 31736 32812 31776
rect 32861 31773 32873 31807
rect 32907 31773 32919 31807
rect 33962 31804 33968 31816
rect 32861 31767 32919 31773
rect 32968 31776 33968 31804
rect 32968 31736 32996 31776
rect 33962 31764 33968 31776
rect 34020 31764 34026 31816
rect 34698 31764 34704 31816
rect 34756 31804 34762 31816
rect 42426 31813 42432 31816
rect 42245 31807 42303 31813
rect 42245 31804 42257 31807
rect 34756 31776 42257 31804
rect 34756 31764 34762 31776
rect 42245 31773 42257 31776
rect 42291 31773 42303 31807
rect 42245 31767 42303 31773
rect 42393 31807 42432 31813
rect 42393 31773 42405 31807
rect 42393 31767 42432 31773
rect 42426 31764 42432 31767
rect 42484 31764 42490 31816
rect 42610 31804 42616 31816
rect 42571 31776 42616 31804
rect 42610 31764 42616 31776
rect 42668 31764 42674 31816
rect 42720 31813 42748 31844
rect 42710 31807 42768 31813
rect 42710 31773 42722 31807
rect 42756 31773 42768 31807
rect 43438 31804 43444 31816
rect 42710 31767 42768 31773
rect 42812 31776 43444 31804
rect 31812 31708 32168 31736
rect 32784 31708 32996 31736
rect 31812 31696 31818 31708
rect 17359 31640 25176 31668
rect 17359 31637 17371 31640
rect 17313 31631 17371 31637
rect 26050 31628 26056 31680
rect 26108 31668 26114 31680
rect 32030 31668 32036 31680
rect 26108 31640 32036 31668
rect 26108 31628 26114 31640
rect 32030 31628 32036 31640
rect 32088 31628 32094 31680
rect 32140 31668 32168 31708
rect 33502 31696 33508 31748
rect 33560 31736 33566 31748
rect 33689 31739 33747 31745
rect 33689 31736 33701 31739
rect 33560 31708 33701 31736
rect 33560 31696 33566 31708
rect 33689 31705 33701 31708
rect 33735 31705 33747 31739
rect 38470 31736 38476 31748
rect 33689 31699 33747 31705
rect 33980 31708 38476 31736
rect 33042 31668 33048 31680
rect 32140 31640 33048 31668
rect 33042 31628 33048 31640
rect 33100 31628 33106 31680
rect 33594 31628 33600 31680
rect 33652 31668 33658 31680
rect 33980 31668 34008 31708
rect 38470 31696 38476 31708
rect 38528 31696 38534 31748
rect 42521 31739 42579 31745
rect 42521 31705 42533 31739
rect 42567 31736 42579 31739
rect 42812 31736 42840 31776
rect 43438 31764 43444 31776
rect 43496 31804 43502 31816
rect 43990 31804 43996 31816
rect 43496 31776 43852 31804
rect 43951 31776 43996 31804
rect 43496 31764 43502 31776
rect 42567 31708 42840 31736
rect 43824 31736 43852 31776
rect 43990 31764 43996 31776
rect 44048 31764 44054 31816
rect 44082 31764 44088 31816
rect 44140 31804 44146 31816
rect 44468 31813 44496 31900
rect 46750 31872 46756 31884
rect 44560 31844 46756 31872
rect 44269 31807 44327 31813
rect 44140 31776 44185 31804
rect 44140 31764 44146 31776
rect 44269 31773 44281 31807
rect 44315 31773 44327 31807
rect 44269 31767 44327 31773
rect 44458 31807 44516 31813
rect 44458 31773 44470 31807
rect 44504 31773 44516 31807
rect 44458 31767 44516 31773
rect 44174 31736 44180 31748
rect 43824 31708 44180 31736
rect 42567 31705 42579 31708
rect 42521 31699 42579 31705
rect 44174 31696 44180 31708
rect 44232 31736 44238 31748
rect 44284 31736 44312 31767
rect 44232 31708 44312 31736
rect 44361 31739 44419 31745
rect 44232 31696 44238 31708
rect 44361 31705 44373 31739
rect 44407 31736 44419 31739
rect 44560 31736 44588 31844
rect 46750 31832 46756 31844
rect 46808 31832 46814 31884
rect 45830 31764 45836 31816
rect 45888 31804 45894 31816
rect 47578 31804 47584 31816
rect 45888 31776 47584 31804
rect 45888 31764 45894 31776
rect 47578 31764 47584 31776
rect 47636 31764 47642 31816
rect 57422 31764 57428 31816
rect 57480 31804 57486 31816
rect 57885 31807 57943 31813
rect 57885 31804 57897 31807
rect 57480 31776 57897 31804
rect 57480 31764 57486 31776
rect 57885 31773 57897 31776
rect 57931 31773 57943 31807
rect 58158 31804 58164 31816
rect 58119 31776 58164 31804
rect 57885 31767 57943 31773
rect 58158 31764 58164 31776
rect 58216 31764 58222 31816
rect 44407 31708 44588 31736
rect 44407 31705 44419 31708
rect 44361 31699 44419 31705
rect 33652 31640 34008 31668
rect 33652 31628 33658 31640
rect 34054 31628 34060 31680
rect 34112 31668 34118 31680
rect 53926 31668 53932 31680
rect 34112 31640 53932 31668
rect 34112 31628 34118 31640
rect 53926 31628 53932 31640
rect 53984 31628 53990 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 24578 31424 24584 31476
rect 24636 31464 24642 31476
rect 24636 31436 31754 31464
rect 24636 31424 24642 31436
rect 17954 31356 17960 31408
rect 18012 31396 18018 31408
rect 19245 31399 19303 31405
rect 18012 31368 18552 31396
rect 18012 31356 18018 31368
rect 1670 31328 1676 31340
rect 1631 31300 1676 31328
rect 1670 31288 1676 31300
rect 1728 31288 1734 31340
rect 18138 31328 18144 31340
rect 18099 31300 18144 31328
rect 18138 31288 18144 31300
rect 18196 31288 18202 31340
rect 18524 31337 18552 31368
rect 19245 31365 19257 31399
rect 19291 31396 19303 31399
rect 19291 31368 22324 31396
rect 19291 31365 19303 31368
rect 19245 31359 19303 31365
rect 18509 31331 18567 31337
rect 18509 31297 18521 31331
rect 18555 31297 18567 31331
rect 19058 31328 19064 31340
rect 19019 31300 19064 31328
rect 18509 31291 18567 31297
rect 19058 31288 19064 31300
rect 19116 31288 19122 31340
rect 19426 31288 19432 31340
rect 19484 31328 19490 31340
rect 19613 31331 19671 31337
rect 19613 31328 19625 31331
rect 19484 31300 19625 31328
rect 19484 31288 19490 31300
rect 19613 31297 19625 31300
rect 19659 31297 19671 31331
rect 19613 31291 19671 31297
rect 20257 31331 20315 31337
rect 20257 31297 20269 31331
rect 20303 31328 20315 31331
rect 20438 31328 20444 31340
rect 20303 31300 20444 31328
rect 20303 31297 20315 31300
rect 20257 31291 20315 31297
rect 20438 31288 20444 31300
rect 20496 31288 20502 31340
rect 22296 31337 22324 31368
rect 25130 31356 25136 31408
rect 25188 31396 25194 31408
rect 25866 31396 25872 31408
rect 25188 31368 25233 31396
rect 25827 31368 25872 31396
rect 25188 31356 25194 31368
rect 25866 31356 25872 31368
rect 25924 31356 25930 31408
rect 31726 31396 31754 31436
rect 32398 31424 32404 31476
rect 32456 31464 32462 31476
rect 32456 31436 36400 31464
rect 32456 31424 32462 31436
rect 31726 31368 34192 31396
rect 24946 31337 24952 31340
rect 22281 31331 22339 31337
rect 22281 31297 22293 31331
rect 22327 31328 22339 31331
rect 24765 31331 24823 31337
rect 22327 31300 23520 31328
rect 22327 31297 22339 31300
rect 22281 31291 22339 31297
rect 20530 31260 20536 31272
rect 20491 31232 20536 31260
rect 20530 31220 20536 31232
rect 20588 31220 20594 31272
rect 22094 31220 22100 31272
rect 22152 31260 22158 31272
rect 22557 31263 22615 31269
rect 22557 31260 22569 31263
rect 22152 31232 22569 31260
rect 22152 31220 22158 31232
rect 22557 31229 22569 31232
rect 22603 31229 22615 31263
rect 23492 31260 23520 31300
rect 24765 31297 24777 31331
rect 24811 31297 24823 31331
rect 24765 31291 24823 31297
rect 24913 31331 24952 31337
rect 24913 31297 24925 31331
rect 24913 31291 24952 31297
rect 24578 31260 24584 31272
rect 23492 31232 24584 31260
rect 22557 31223 22615 31229
rect 24578 31220 24584 31232
rect 24636 31220 24642 31272
rect 21542 31152 21548 31204
rect 21600 31192 21606 31204
rect 24780 31192 24808 31291
rect 24946 31288 24952 31291
rect 25004 31288 25010 31340
rect 25041 31331 25099 31337
rect 25041 31297 25053 31331
rect 25087 31297 25099 31331
rect 25041 31291 25099 31297
rect 25271 31331 25329 31337
rect 25271 31297 25283 31331
rect 25317 31328 25329 31331
rect 26050 31328 26056 31340
rect 25317 31300 25912 31328
rect 26011 31300 26056 31328
rect 25317 31297 25329 31300
rect 25271 31291 25329 31297
rect 25056 31260 25084 31291
rect 25774 31260 25780 31272
rect 25056 31232 25780 31260
rect 25774 31220 25780 31232
rect 25832 31220 25838 31272
rect 25884 31260 25912 31300
rect 26050 31288 26056 31300
rect 26108 31288 26114 31340
rect 32030 31288 32036 31340
rect 32088 31328 32094 31340
rect 33594 31328 33600 31340
rect 32088 31300 33600 31328
rect 32088 31288 32094 31300
rect 33594 31288 33600 31300
rect 33652 31288 33658 31340
rect 33778 31328 33784 31340
rect 33739 31300 33784 31328
rect 33778 31288 33784 31300
rect 33836 31288 33842 31340
rect 34054 31328 34060 31340
rect 34015 31300 34060 31328
rect 34054 31288 34060 31300
rect 34112 31288 34118 31340
rect 34164 31328 34192 31368
rect 34790 31356 34796 31408
rect 34848 31396 34854 31408
rect 35250 31396 35256 31408
rect 34848 31368 35020 31396
rect 35211 31368 35256 31396
rect 34848 31356 34854 31368
rect 34992 31337 35020 31368
rect 35250 31356 35256 31368
rect 35308 31356 35314 31408
rect 35158 31337 35164 31340
rect 34977 31331 35035 31337
rect 34164 31300 34928 31328
rect 25958 31260 25964 31272
rect 25884 31232 25964 31260
rect 25958 31220 25964 31232
rect 26016 31220 26022 31272
rect 26326 31260 26332 31272
rect 26287 31232 26332 31260
rect 26326 31220 26332 31232
rect 26384 31220 26390 31272
rect 33134 31220 33140 31272
rect 33192 31260 33198 31272
rect 34241 31263 34299 31269
rect 34241 31260 34253 31263
rect 33192 31232 34253 31260
rect 33192 31220 33198 31232
rect 34241 31229 34253 31232
rect 34287 31229 34299 31263
rect 34900 31260 34928 31300
rect 34977 31297 34989 31331
rect 35023 31297 35035 31331
rect 34977 31291 35035 31297
rect 35125 31331 35164 31337
rect 35125 31297 35137 31331
rect 35125 31291 35164 31297
rect 35158 31288 35164 31291
rect 35216 31288 35222 31340
rect 35342 31328 35348 31340
rect 35303 31300 35348 31328
rect 35342 31288 35348 31300
rect 35400 31288 35406 31340
rect 36372 31337 36400 31436
rect 35442 31331 35500 31337
rect 35442 31297 35454 31331
rect 35488 31297 35500 31331
rect 35442 31291 35500 31297
rect 36357 31331 36415 31337
rect 36357 31297 36369 31331
rect 36403 31297 36415 31331
rect 36357 31291 36415 31297
rect 35452 31260 35480 31291
rect 34900 31232 35480 31260
rect 34241 31223 34299 31229
rect 36262 31220 36268 31272
rect 36320 31260 36326 31272
rect 36541 31263 36599 31269
rect 36541 31260 36553 31263
rect 36320 31232 36553 31260
rect 36320 31220 36326 31232
rect 36541 31229 36553 31232
rect 36587 31260 36599 31263
rect 37458 31260 37464 31272
rect 36587 31232 37464 31260
rect 36587 31229 36599 31232
rect 36541 31223 36599 31229
rect 37458 31220 37464 31232
rect 37516 31220 37522 31272
rect 43070 31220 43076 31272
rect 43128 31260 43134 31272
rect 52270 31260 52276 31272
rect 43128 31232 52276 31260
rect 43128 31220 43134 31232
rect 52270 31220 52276 31232
rect 52328 31220 52334 31272
rect 31110 31192 31116 31204
rect 21600 31164 31116 31192
rect 21600 31152 21606 31164
rect 31110 31152 31116 31164
rect 31168 31152 31174 31204
rect 33873 31195 33931 31201
rect 33873 31161 33885 31195
rect 33919 31192 33931 31195
rect 35621 31195 35679 31201
rect 35621 31192 35633 31195
rect 33919 31164 35633 31192
rect 33919 31161 33931 31164
rect 33873 31155 33931 31161
rect 35621 31161 35633 31164
rect 35667 31161 35679 31195
rect 35621 31155 35679 31161
rect 44082 31152 44088 31204
rect 44140 31192 44146 31204
rect 53006 31192 53012 31204
rect 44140 31164 53012 31192
rect 44140 31152 44146 31164
rect 53006 31152 53012 31164
rect 53064 31152 53070 31204
rect 1765 31127 1823 31133
rect 1765 31093 1777 31127
rect 1811 31124 1823 31127
rect 23290 31124 23296 31136
rect 1811 31096 23296 31124
rect 1811 31093 1823 31096
rect 1765 31087 1823 31093
rect 23290 31084 23296 31096
rect 23348 31084 23354 31136
rect 24578 31084 24584 31136
rect 24636 31124 24642 31136
rect 25409 31127 25467 31133
rect 25409 31124 25421 31127
rect 24636 31096 25421 31124
rect 24636 31084 24642 31096
rect 25409 31093 25421 31096
rect 25455 31093 25467 31127
rect 25409 31087 25467 31093
rect 29822 31084 29828 31136
rect 29880 31124 29886 31136
rect 37274 31124 37280 31136
rect 29880 31096 37280 31124
rect 29880 31084 29886 31096
rect 37274 31084 37280 31096
rect 37332 31084 37338 31136
rect 42426 31084 42432 31136
rect 42484 31124 42490 31136
rect 52914 31124 52920 31136
rect 42484 31096 52920 31124
rect 42484 31084 42490 31096
rect 52914 31084 52920 31096
rect 52972 31084 52978 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 6914 30880 6920 30932
rect 6972 30920 6978 30932
rect 35342 30920 35348 30932
rect 6972 30892 35348 30920
rect 6972 30880 6978 30892
rect 35342 30880 35348 30892
rect 35400 30880 35406 30932
rect 35802 30880 35808 30932
rect 35860 30920 35866 30932
rect 38289 30923 38347 30929
rect 38289 30920 38301 30923
rect 35860 30892 38301 30920
rect 35860 30880 35866 30892
rect 38289 30889 38301 30892
rect 38335 30889 38347 30923
rect 38289 30883 38347 30889
rect 17954 30812 17960 30864
rect 18012 30812 18018 30864
rect 18874 30812 18880 30864
rect 18932 30852 18938 30864
rect 23566 30852 23572 30864
rect 18932 30824 23428 30852
rect 23527 30824 23572 30852
rect 18932 30812 18938 30824
rect 17494 30784 17500 30796
rect 17455 30756 17500 30784
rect 17494 30744 17500 30756
rect 17552 30744 17558 30796
rect 17972 30784 18000 30812
rect 20070 30784 20076 30796
rect 17972 30756 18092 30784
rect 18064 30725 18092 30756
rect 19720 30756 20076 30784
rect 17957 30719 18015 30725
rect 17957 30685 17969 30719
rect 18003 30685 18015 30719
rect 17957 30679 18015 30685
rect 18049 30719 18107 30725
rect 18049 30685 18061 30719
rect 18095 30716 18107 30719
rect 18322 30716 18328 30728
rect 18095 30688 18328 30716
rect 18095 30685 18107 30688
rect 18049 30679 18107 30685
rect 1670 30648 1676 30660
rect 1631 30620 1676 30648
rect 1670 30608 1676 30620
rect 1728 30608 1734 30660
rect 17402 30608 17408 30660
rect 17460 30648 17466 30660
rect 17589 30651 17647 30657
rect 17589 30648 17601 30651
rect 17460 30620 17601 30648
rect 17460 30608 17466 30620
rect 17589 30617 17601 30620
rect 17635 30648 17647 30651
rect 17770 30648 17776 30660
rect 17635 30620 17776 30648
rect 17635 30617 17647 30620
rect 17589 30611 17647 30617
rect 17770 30608 17776 30620
rect 17828 30608 17834 30660
rect 17972 30648 18000 30679
rect 18322 30676 18328 30688
rect 18380 30676 18386 30728
rect 18509 30719 18567 30725
rect 18509 30685 18521 30719
rect 18555 30716 18567 30719
rect 19426 30716 19432 30728
rect 18555 30688 19432 30716
rect 18555 30685 18567 30688
rect 18509 30679 18567 30685
rect 19426 30676 19432 30688
rect 19484 30676 19490 30728
rect 19720 30725 19748 30756
rect 20070 30744 20076 30756
rect 20128 30744 20134 30796
rect 21542 30784 21548 30796
rect 21503 30756 21548 30784
rect 21542 30744 21548 30756
rect 21600 30744 21606 30796
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30685 19763 30719
rect 19978 30716 19984 30728
rect 19939 30688 19984 30716
rect 19705 30679 19763 30685
rect 19978 30676 19984 30688
rect 20036 30676 20042 30728
rect 20441 30719 20499 30725
rect 20441 30685 20453 30719
rect 20487 30716 20499 30719
rect 20530 30716 20536 30728
rect 20487 30688 20536 30716
rect 20487 30685 20499 30688
rect 20441 30679 20499 30685
rect 18340 30648 18368 30676
rect 20456 30648 20484 30679
rect 20530 30676 20536 30688
rect 20588 30676 20594 30728
rect 20622 30676 20628 30728
rect 20680 30716 20686 30728
rect 20717 30719 20775 30725
rect 20717 30716 20729 30719
rect 20680 30688 20729 30716
rect 20680 30676 20686 30688
rect 20717 30685 20729 30688
rect 20763 30685 20775 30719
rect 20717 30679 20775 30685
rect 22005 30719 22063 30725
rect 22005 30685 22017 30719
rect 22051 30685 22063 30719
rect 22186 30716 22192 30728
rect 22147 30688 22192 30716
rect 22005 30679 22063 30685
rect 17972 30620 18092 30648
rect 18340 30620 20484 30648
rect 1765 30583 1823 30589
rect 1765 30549 1777 30583
rect 1811 30580 1823 30583
rect 16298 30580 16304 30592
rect 1811 30552 16304 30580
rect 1811 30549 1823 30552
rect 1765 30543 1823 30549
rect 16298 30540 16304 30552
rect 16356 30540 16362 30592
rect 18064 30580 18092 30620
rect 18138 30580 18144 30592
rect 18051 30552 18144 30580
rect 18138 30540 18144 30552
rect 18196 30580 18202 30592
rect 18782 30580 18788 30592
rect 18196 30552 18788 30580
rect 18196 30540 18202 30552
rect 18782 30540 18788 30552
rect 18840 30540 18846 30592
rect 19334 30540 19340 30592
rect 19392 30580 19398 30592
rect 20530 30580 20536 30592
rect 19392 30552 20536 30580
rect 19392 30540 19398 30552
rect 20530 30540 20536 30552
rect 20588 30580 20594 30592
rect 20625 30583 20683 30589
rect 20625 30580 20637 30583
rect 20588 30552 20637 30580
rect 20588 30540 20594 30552
rect 20625 30549 20637 30552
rect 20671 30549 20683 30583
rect 20625 30543 20683 30549
rect 20990 30540 20996 30592
rect 21048 30580 21054 30592
rect 22020 30580 22048 30679
rect 22186 30676 22192 30688
rect 22244 30676 22250 30728
rect 22373 30719 22431 30725
rect 22373 30685 22385 30719
rect 22419 30716 22431 30719
rect 23014 30716 23020 30728
rect 22419 30688 23020 30716
rect 22419 30685 22431 30688
rect 22373 30679 22431 30685
rect 23014 30676 23020 30688
rect 23072 30676 23078 30728
rect 23290 30716 23296 30728
rect 23251 30688 23296 30716
rect 23290 30676 23296 30688
rect 23348 30676 23354 30728
rect 23400 30725 23428 30824
rect 23566 30812 23572 30824
rect 23624 30812 23630 30864
rect 43806 30852 43812 30864
rect 30668 30824 43812 30852
rect 30466 30784 30472 30796
rect 30427 30756 30472 30784
rect 30466 30744 30472 30756
rect 30524 30744 30530 30796
rect 23385 30719 23443 30725
rect 23385 30685 23397 30719
rect 23431 30685 23443 30719
rect 24578 30716 24584 30728
rect 24539 30688 24584 30716
rect 23385 30679 23443 30685
rect 24578 30676 24584 30688
rect 24636 30676 24642 30728
rect 24762 30716 24768 30728
rect 24723 30688 24768 30716
rect 24762 30676 24768 30688
rect 24820 30676 24826 30728
rect 28534 30676 28540 30728
rect 28592 30716 28598 30728
rect 30377 30719 30435 30725
rect 28592 30688 29868 30716
rect 28592 30676 28598 30688
rect 22204 30648 22232 30676
rect 23201 30651 23259 30657
rect 23201 30648 23213 30651
rect 22204 30620 23213 30648
rect 23201 30617 23213 30620
rect 23247 30617 23259 30651
rect 29730 30648 29736 30660
rect 29691 30620 29736 30648
rect 23201 30611 23259 30617
rect 29730 30608 29736 30620
rect 29788 30608 29794 30660
rect 29840 30648 29868 30688
rect 30377 30685 30389 30719
rect 30423 30716 30435 30719
rect 30668 30716 30696 30824
rect 43806 30812 43812 30824
rect 43864 30812 43870 30864
rect 31110 30744 31116 30796
rect 31168 30784 31174 30796
rect 31168 30756 35664 30784
rect 31168 30744 31174 30756
rect 35636 30728 35664 30756
rect 36096 30756 37228 30784
rect 36096 30728 36124 30756
rect 30423 30688 30696 30716
rect 30745 30719 30803 30725
rect 30423 30685 30435 30688
rect 30377 30679 30435 30685
rect 30745 30685 30757 30719
rect 30791 30685 30803 30719
rect 30745 30679 30803 30685
rect 30929 30719 30987 30725
rect 30929 30685 30941 30719
rect 30975 30716 30987 30719
rect 31754 30716 31760 30728
rect 30975 30688 31760 30716
rect 30975 30685 30987 30688
rect 30929 30679 30987 30685
rect 30760 30648 30788 30679
rect 31754 30676 31760 30688
rect 31812 30676 31818 30728
rect 35618 30676 35624 30728
rect 35676 30716 35682 30728
rect 35805 30719 35863 30725
rect 35805 30716 35817 30719
rect 35676 30688 35817 30716
rect 35676 30676 35682 30688
rect 35805 30685 35817 30688
rect 35851 30685 35863 30719
rect 35805 30679 35863 30685
rect 35894 30676 35900 30728
rect 35952 30716 35958 30728
rect 35952 30688 35997 30716
rect 35952 30676 35958 30688
rect 36078 30676 36084 30728
rect 36136 30716 36142 30728
rect 36136 30688 36181 30716
rect 36136 30676 36142 30688
rect 36262 30676 36268 30728
rect 36320 30725 36326 30728
rect 36320 30716 36328 30725
rect 36906 30716 36912 30728
rect 36320 30688 36365 30716
rect 36867 30688 36912 30716
rect 36320 30679 36328 30688
rect 36320 30676 36326 30679
rect 36906 30676 36912 30688
rect 36964 30676 36970 30728
rect 36998 30676 37004 30728
rect 37056 30716 37062 30728
rect 37200 30725 37228 30756
rect 37185 30719 37243 30725
rect 37056 30688 37101 30716
rect 37056 30676 37062 30688
rect 37185 30685 37197 30719
rect 37231 30685 37243 30719
rect 37185 30679 37243 30685
rect 37274 30676 37280 30728
rect 37332 30716 37338 30728
rect 37458 30725 37464 30728
rect 37415 30719 37464 30725
rect 37332 30688 37377 30716
rect 37332 30676 37338 30688
rect 37415 30685 37427 30719
rect 37461 30685 37464 30719
rect 37415 30679 37464 30685
rect 37458 30676 37464 30679
rect 37516 30676 37522 30728
rect 38197 30719 38255 30725
rect 38197 30685 38209 30719
rect 38243 30716 38255 30719
rect 38654 30716 38660 30728
rect 38243 30688 38660 30716
rect 38243 30685 38255 30688
rect 38197 30679 38255 30685
rect 38654 30676 38660 30688
rect 38712 30676 38718 30728
rect 57974 30716 57980 30728
rect 57935 30688 57980 30716
rect 57974 30676 57980 30688
rect 58032 30676 58038 30728
rect 36173 30651 36231 30657
rect 36173 30648 36185 30651
rect 29840 30620 30788 30648
rect 36004 30620 36185 30648
rect 22094 30580 22100 30592
rect 21048 30552 22100 30580
rect 21048 30540 21054 30552
rect 22094 30540 22100 30552
rect 22152 30540 22158 30592
rect 24854 30580 24860 30592
rect 24815 30552 24860 30580
rect 24854 30540 24860 30552
rect 24912 30540 24918 30592
rect 27430 30540 27436 30592
rect 27488 30580 27494 30592
rect 36004 30580 36032 30620
rect 36173 30617 36185 30620
rect 36219 30617 36231 30651
rect 38013 30651 38071 30657
rect 38013 30648 38025 30651
rect 36173 30611 36231 30617
rect 37384 30620 38025 30648
rect 27488 30552 36032 30580
rect 36449 30583 36507 30589
rect 27488 30540 27494 30552
rect 36449 30549 36461 30583
rect 36495 30580 36507 30583
rect 37384 30580 37412 30620
rect 38013 30617 38025 30620
rect 38059 30617 38071 30651
rect 38013 30611 38071 30617
rect 37550 30580 37556 30592
rect 36495 30552 37412 30580
rect 37511 30552 37556 30580
rect 36495 30549 36507 30552
rect 36449 30543 36507 30549
rect 37550 30540 37556 30552
rect 37608 30540 37614 30592
rect 58066 30580 58072 30592
rect 58027 30552 58072 30580
rect 58066 30540 58072 30552
rect 58124 30540 58130 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 19610 30376 19616 30388
rect 19523 30348 19616 30376
rect 19610 30336 19616 30348
rect 19668 30376 19674 30388
rect 20070 30376 20076 30388
rect 19668 30348 20076 30376
rect 19668 30336 19674 30348
rect 20070 30336 20076 30348
rect 20128 30336 20134 30388
rect 33778 30336 33784 30388
rect 33836 30376 33842 30388
rect 36262 30376 36268 30388
rect 33836 30348 36268 30376
rect 33836 30336 33842 30348
rect 36262 30336 36268 30348
rect 36320 30336 36326 30388
rect 36906 30376 36912 30388
rect 36372 30348 36912 30376
rect 17494 30268 17500 30320
rect 17552 30308 17558 30320
rect 17773 30311 17831 30317
rect 17773 30308 17785 30311
rect 17552 30280 17785 30308
rect 17552 30268 17558 30280
rect 17773 30277 17785 30280
rect 17819 30277 17831 30311
rect 17773 30271 17831 30277
rect 17862 30268 17868 30320
rect 17920 30308 17926 30320
rect 20622 30308 20628 30320
rect 17920 30280 20392 30308
rect 20583 30280 20628 30308
rect 17920 30268 17926 30280
rect 18233 30243 18291 30249
rect 18233 30209 18245 30243
rect 18279 30209 18291 30243
rect 18233 30203 18291 30209
rect 18248 30104 18276 30203
rect 18322 30200 18328 30252
rect 18380 30240 18386 30252
rect 19337 30243 19395 30249
rect 18380 30212 18425 30240
rect 18380 30200 18386 30212
rect 19337 30209 19349 30243
rect 19383 30240 19395 30243
rect 20070 30240 20076 30252
rect 19383 30212 20076 30240
rect 19383 30209 19395 30212
rect 19337 30203 19395 30209
rect 20070 30200 20076 30212
rect 20128 30200 20134 30252
rect 20257 30243 20315 30249
rect 20257 30209 20269 30243
rect 20303 30209 20315 30243
rect 20364 30240 20392 30280
rect 20622 30268 20628 30280
rect 20680 30268 20686 30320
rect 22557 30311 22615 30317
rect 22557 30277 22569 30311
rect 22603 30308 22615 30311
rect 23474 30308 23480 30320
rect 22603 30280 23480 30308
rect 22603 30277 22615 30280
rect 22557 30271 22615 30277
rect 23474 30268 23480 30280
rect 23532 30268 23538 30320
rect 35618 30268 35624 30320
rect 35676 30308 35682 30320
rect 36372 30308 36400 30348
rect 36906 30336 36912 30348
rect 36964 30376 36970 30388
rect 42886 30376 42892 30388
rect 36964 30348 42892 30376
rect 36964 30336 36970 30348
rect 42886 30336 42892 30348
rect 42944 30376 42950 30388
rect 43162 30376 43168 30388
rect 42944 30348 43168 30376
rect 42944 30336 42950 30348
rect 43162 30336 43168 30348
rect 43220 30336 43226 30388
rect 35676 30280 36400 30308
rect 37461 30311 37519 30317
rect 35676 30268 35682 30280
rect 37461 30277 37473 30311
rect 37507 30308 37519 30311
rect 37550 30308 37556 30320
rect 37507 30280 37556 30308
rect 37507 30277 37519 30280
rect 37461 30271 37519 30277
rect 37550 30268 37556 30280
rect 37608 30268 37614 30320
rect 22097 30243 22155 30249
rect 22097 30240 22109 30243
rect 20364 30212 22109 30240
rect 20257 30203 20315 30209
rect 22097 30209 22109 30212
rect 22143 30240 22155 30243
rect 22186 30240 22192 30252
rect 22143 30212 22192 30240
rect 22143 30209 22155 30212
rect 22097 30203 22155 30209
rect 18785 30175 18843 30181
rect 18785 30141 18797 30175
rect 18831 30172 18843 30175
rect 19426 30172 19432 30184
rect 18831 30144 19432 30172
rect 18831 30141 18843 30144
rect 18785 30135 18843 30141
rect 19426 30132 19432 30144
rect 19484 30172 19490 30184
rect 19978 30172 19984 30184
rect 19484 30144 19984 30172
rect 19484 30132 19490 30144
rect 19978 30132 19984 30144
rect 20036 30132 20042 30184
rect 19610 30104 19616 30116
rect 18248 30076 19616 30104
rect 19610 30064 19616 30076
rect 19668 30064 19674 30116
rect 20272 30104 20300 30203
rect 22186 30200 22192 30212
rect 22244 30200 22250 30252
rect 37645 30243 37703 30249
rect 37645 30209 37657 30243
rect 37691 30240 37703 30243
rect 42334 30240 42340 30252
rect 37691 30212 42340 30240
rect 37691 30209 37703 30212
rect 37645 30203 37703 30209
rect 42334 30200 42340 30212
rect 42392 30200 42398 30252
rect 21910 30132 21916 30184
rect 21968 30172 21974 30184
rect 22005 30175 22063 30181
rect 22005 30172 22017 30175
rect 21968 30144 22017 30172
rect 21968 30132 21974 30144
rect 22005 30141 22017 30144
rect 22051 30172 22063 30175
rect 23014 30172 23020 30184
rect 22051 30144 23020 30172
rect 22051 30141 22063 30144
rect 22005 30135 22063 30141
rect 23014 30132 23020 30144
rect 23072 30132 23078 30184
rect 20990 30104 20996 30116
rect 20272 30076 20996 30104
rect 20990 30064 20996 30076
rect 21048 30064 21054 30116
rect 37642 29996 37648 30048
rect 37700 30036 37706 30048
rect 37737 30039 37795 30045
rect 37737 30036 37749 30039
rect 37700 30008 37749 30036
rect 37700 29996 37706 30008
rect 37737 30005 37749 30008
rect 37783 30005 37795 30039
rect 37737 29999 37795 30005
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 20438 29792 20444 29844
rect 20496 29832 20502 29844
rect 21729 29835 21787 29841
rect 21729 29832 21741 29835
rect 20496 29804 21741 29832
rect 20496 29792 20502 29804
rect 21729 29801 21741 29804
rect 21775 29801 21787 29835
rect 21729 29795 21787 29801
rect 34790 29792 34796 29844
rect 34848 29832 34854 29844
rect 35437 29835 35495 29841
rect 35437 29832 35449 29835
rect 34848 29804 35449 29832
rect 34848 29792 34854 29804
rect 35437 29801 35449 29804
rect 35483 29801 35495 29835
rect 35437 29795 35495 29801
rect 36814 29792 36820 29844
rect 36872 29832 36878 29844
rect 43806 29832 43812 29844
rect 36872 29804 41414 29832
rect 43767 29804 43812 29832
rect 36872 29792 36878 29804
rect 41386 29764 41414 29804
rect 43806 29792 43812 29804
rect 43864 29792 43870 29844
rect 53466 29764 53472 29776
rect 41386 29736 53472 29764
rect 53466 29724 53472 29736
rect 53524 29724 53530 29776
rect 6178 29656 6184 29708
rect 6236 29696 6242 29708
rect 17678 29696 17684 29708
rect 6236 29668 17684 29696
rect 6236 29656 6242 29668
rect 17678 29656 17684 29668
rect 17736 29656 17742 29708
rect 22830 29656 22836 29708
rect 22888 29696 22894 29708
rect 34790 29696 34796 29708
rect 22888 29668 34796 29696
rect 22888 29656 22894 29668
rect 34790 29656 34796 29668
rect 34848 29656 34854 29708
rect 34974 29656 34980 29708
rect 35032 29696 35038 29708
rect 43070 29696 43076 29708
rect 35032 29668 43076 29696
rect 35032 29656 35038 29668
rect 43070 29656 43076 29668
rect 43128 29656 43134 29708
rect 47210 29696 47216 29708
rect 43364 29668 47216 29696
rect 1581 29631 1639 29637
rect 1581 29597 1593 29631
rect 1627 29628 1639 29631
rect 15194 29628 15200 29640
rect 1627 29600 6914 29628
rect 15155 29600 15200 29628
rect 1627 29597 1639 29600
rect 1581 29591 1639 29597
rect 1854 29560 1860 29572
rect 1815 29532 1860 29560
rect 1854 29520 1860 29532
rect 1912 29520 1918 29572
rect 6886 29560 6914 29600
rect 15194 29588 15200 29600
rect 15252 29588 15258 29640
rect 15351 29631 15409 29637
rect 15351 29597 15363 29631
rect 15397 29628 15409 29631
rect 17862 29628 17868 29640
rect 15397 29600 17868 29628
rect 15397 29597 15409 29600
rect 15351 29591 15409 29597
rect 17862 29588 17868 29600
rect 17920 29588 17926 29640
rect 19150 29588 19156 29640
rect 19208 29628 19214 29640
rect 19334 29628 19340 29640
rect 19208 29600 19340 29628
rect 19208 29588 19214 29600
rect 19334 29588 19340 29600
rect 19392 29628 19398 29640
rect 19521 29631 19579 29637
rect 19521 29628 19533 29631
rect 19392 29600 19533 29628
rect 19392 29588 19398 29600
rect 19521 29597 19533 29600
rect 19567 29597 19579 29631
rect 19521 29591 19579 29597
rect 19889 29631 19947 29637
rect 19889 29597 19901 29631
rect 19935 29597 19947 29631
rect 20438 29628 20444 29640
rect 20399 29600 20444 29628
rect 19889 29591 19947 29597
rect 15565 29563 15623 29569
rect 15565 29560 15577 29563
rect 6886 29532 15577 29560
rect 15565 29529 15577 29532
rect 15611 29529 15623 29563
rect 15565 29523 15623 29529
rect 18782 29520 18788 29572
rect 18840 29560 18846 29572
rect 19904 29560 19932 29591
rect 20438 29588 20444 29600
rect 20496 29588 20502 29640
rect 20990 29628 20996 29640
rect 20951 29600 20996 29628
rect 20990 29588 20996 29600
rect 21048 29588 21054 29640
rect 34882 29628 34888 29640
rect 34843 29600 34888 29628
rect 34882 29588 34888 29600
rect 34940 29588 34946 29640
rect 35161 29631 35219 29637
rect 35161 29628 35173 29631
rect 34992 29600 35173 29628
rect 18840 29532 19932 29560
rect 18840 29520 18846 29532
rect 20714 29520 20720 29572
rect 20772 29560 20778 29572
rect 21637 29563 21695 29569
rect 21637 29560 21649 29563
rect 20772 29532 21649 29560
rect 20772 29520 20778 29532
rect 21637 29529 21649 29532
rect 21683 29529 21695 29563
rect 21637 29523 21695 29529
rect 34238 29520 34244 29572
rect 34296 29560 34302 29572
rect 34992 29560 35020 29600
rect 35161 29597 35173 29600
rect 35207 29597 35219 29631
rect 35161 29591 35219 29597
rect 35253 29631 35311 29637
rect 35253 29597 35265 29631
rect 35299 29628 35311 29631
rect 36170 29628 36176 29640
rect 35299 29600 36176 29628
rect 35299 29597 35311 29600
rect 35253 29591 35311 29597
rect 36170 29588 36176 29600
rect 36228 29588 36234 29640
rect 43162 29628 43168 29640
rect 43123 29600 43168 29628
rect 43162 29588 43168 29600
rect 43220 29588 43226 29640
rect 43364 29637 43392 29668
rect 47210 29656 47216 29668
rect 47268 29656 47274 29708
rect 58158 29696 58164 29708
rect 58119 29668 58164 29696
rect 58158 29656 58164 29668
rect 58216 29656 58222 29708
rect 43313 29631 43392 29637
rect 43313 29597 43325 29631
rect 43359 29600 43392 29631
rect 43359 29597 43371 29600
rect 43313 29591 43371 29597
rect 43438 29588 43444 29640
rect 43496 29628 43502 29640
rect 43671 29631 43729 29637
rect 43496 29600 43541 29628
rect 43496 29588 43502 29600
rect 43671 29597 43683 29631
rect 43717 29628 43729 29631
rect 46106 29628 46112 29640
rect 43717 29600 46112 29628
rect 43717 29597 43729 29600
rect 43671 29591 43729 29597
rect 46106 29588 46112 29600
rect 46164 29588 46170 29640
rect 57885 29631 57943 29637
rect 57885 29628 57897 29631
rect 51046 29600 57897 29628
rect 34296 29532 35020 29560
rect 34296 29520 34302 29532
rect 35066 29520 35072 29572
rect 35124 29560 35130 29572
rect 43533 29563 43591 29569
rect 35124 29532 35169 29560
rect 35124 29520 35130 29532
rect 43533 29529 43545 29563
rect 43579 29560 43591 29563
rect 43579 29532 43668 29560
rect 43579 29529 43591 29532
rect 43533 29523 43591 29529
rect 43640 29504 43668 29532
rect 44634 29520 44640 29572
rect 44692 29560 44698 29572
rect 51046 29560 51074 29600
rect 57885 29597 57897 29600
rect 57931 29597 57943 29631
rect 57885 29591 57943 29597
rect 57054 29560 57060 29572
rect 44692 29532 51074 29560
rect 57015 29532 57060 29560
rect 44692 29520 44698 29532
rect 57054 29520 57060 29532
rect 57112 29520 57118 29572
rect 18874 29452 18880 29504
rect 18932 29492 18938 29504
rect 19521 29495 19579 29501
rect 19521 29492 19533 29495
rect 18932 29464 19533 29492
rect 18932 29452 18938 29464
rect 19521 29461 19533 29464
rect 19567 29461 19579 29495
rect 19521 29455 19579 29461
rect 43622 29452 43628 29504
rect 43680 29452 43686 29504
rect 57146 29492 57152 29504
rect 57107 29464 57152 29492
rect 57146 29452 57152 29464
rect 57204 29452 57210 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 19426 29248 19432 29300
rect 19484 29288 19490 29300
rect 19613 29291 19671 29297
rect 19613 29288 19625 29291
rect 19484 29260 19625 29288
rect 19484 29248 19490 29260
rect 19613 29257 19625 29260
rect 19659 29257 19671 29291
rect 24394 29288 24400 29300
rect 24355 29260 24400 29288
rect 19613 29251 19671 29257
rect 24394 29248 24400 29260
rect 24452 29248 24458 29300
rect 32858 29248 32864 29300
rect 32916 29288 32922 29300
rect 35066 29288 35072 29300
rect 32916 29260 35072 29288
rect 32916 29248 32922 29260
rect 35066 29248 35072 29260
rect 35124 29248 35130 29300
rect 43070 29248 43076 29300
rect 43128 29288 43134 29300
rect 49050 29288 49056 29300
rect 43128 29260 49056 29288
rect 43128 29248 43134 29260
rect 49050 29248 49056 29260
rect 49108 29248 49114 29300
rect 18601 29223 18659 29229
rect 18601 29189 18613 29223
rect 18647 29220 18659 29223
rect 20438 29220 20444 29232
rect 18647 29192 20444 29220
rect 18647 29189 18659 29192
rect 18601 29183 18659 29189
rect 20438 29180 20444 29192
rect 20496 29180 20502 29232
rect 34882 29180 34888 29232
rect 34940 29220 34946 29232
rect 37274 29220 37280 29232
rect 34940 29192 37280 29220
rect 34940 29180 34946 29192
rect 37274 29180 37280 29192
rect 37332 29180 37338 29232
rect 1581 29155 1639 29161
rect 1581 29121 1593 29155
rect 1627 29152 1639 29155
rect 2866 29152 2872 29164
rect 1627 29124 2872 29152
rect 1627 29121 1639 29124
rect 1581 29115 1639 29121
rect 2866 29112 2872 29124
rect 2924 29112 2930 29164
rect 18414 29112 18420 29164
rect 18472 29152 18478 29164
rect 18693 29155 18751 29161
rect 18693 29152 18705 29155
rect 18472 29124 18705 29152
rect 18472 29112 18478 29124
rect 18693 29121 18705 29124
rect 18739 29121 18751 29155
rect 18693 29115 18751 29121
rect 18782 29112 18788 29164
rect 18840 29152 18846 29164
rect 19429 29155 19487 29161
rect 19429 29152 19441 29155
rect 18840 29124 18885 29152
rect 18984 29124 19441 29152
rect 18840 29112 18846 29124
rect 1762 29084 1768 29096
rect 1723 29056 1768 29084
rect 1762 29044 1768 29056
rect 1820 29044 1826 29096
rect 18049 29087 18107 29093
rect 18049 29053 18061 29087
rect 18095 29053 18107 29087
rect 18049 29047 18107 29053
rect 18064 29016 18092 29047
rect 18138 29044 18144 29096
rect 18196 29084 18202 29096
rect 18233 29087 18291 29093
rect 18233 29084 18245 29087
rect 18196 29056 18245 29084
rect 18196 29044 18202 29056
rect 18233 29053 18245 29056
rect 18279 29053 18291 29087
rect 18233 29047 18291 29053
rect 18322 29044 18328 29096
rect 18380 29084 18386 29096
rect 18984 29084 19012 29124
rect 19429 29121 19441 29124
rect 19475 29121 19487 29155
rect 19429 29115 19487 29121
rect 19518 29112 19524 29164
rect 19576 29152 19582 29164
rect 20625 29155 20683 29161
rect 20625 29152 20637 29155
rect 19576 29124 20637 29152
rect 19576 29112 19582 29124
rect 20625 29121 20637 29124
rect 20671 29121 20683 29155
rect 20625 29115 20683 29121
rect 23753 29155 23811 29161
rect 23753 29121 23765 29155
rect 23799 29152 23811 29155
rect 24118 29152 24124 29164
rect 23799 29124 24124 29152
rect 23799 29121 23811 29124
rect 23753 29115 23811 29121
rect 24118 29112 24124 29124
rect 24176 29112 24182 29164
rect 24210 29112 24216 29164
rect 24268 29152 24274 29164
rect 25314 29152 25320 29164
rect 24268 29124 25320 29152
rect 24268 29112 24274 29124
rect 25314 29112 25320 29124
rect 25372 29112 25378 29164
rect 31294 29112 31300 29164
rect 31352 29152 31358 29164
rect 57146 29152 57152 29164
rect 31352 29124 57152 29152
rect 31352 29112 31358 29124
rect 57146 29112 57152 29124
rect 57204 29112 57210 29164
rect 19150 29084 19156 29096
rect 18380 29056 19012 29084
rect 19076 29056 19156 29084
rect 18380 29044 18386 29056
rect 19076 29016 19104 29056
rect 19150 29044 19156 29056
rect 19208 29084 19214 29096
rect 19610 29084 19616 29096
rect 19208 29056 19616 29084
rect 19208 29044 19214 29056
rect 19610 29044 19616 29056
rect 19668 29044 19674 29096
rect 26418 29044 26424 29096
rect 26476 29084 26482 29096
rect 31018 29084 31024 29096
rect 26476 29056 31024 29084
rect 26476 29044 26482 29056
rect 31018 29044 31024 29056
rect 31076 29044 31082 29096
rect 20809 29019 20867 29025
rect 20809 29016 20821 29019
rect 18064 28988 19104 29016
rect 19444 28988 20821 29016
rect 18414 28908 18420 28960
rect 18472 28948 18478 28960
rect 19058 28948 19064 28960
rect 18472 28920 19064 28948
rect 18472 28908 18478 28920
rect 19058 28908 19064 28920
rect 19116 28948 19122 28960
rect 19444 28948 19472 28988
rect 20809 28985 20821 28988
rect 20855 29016 20867 29019
rect 20990 29016 20996 29028
rect 20855 28988 20996 29016
rect 20855 28985 20867 28988
rect 20809 28979 20867 28985
rect 20990 28976 20996 28988
rect 21048 28976 21054 29028
rect 24302 28976 24308 29028
rect 24360 29016 24366 29028
rect 27706 29016 27712 29028
rect 24360 28988 27712 29016
rect 24360 28976 24366 28988
rect 27706 28976 27712 28988
rect 27764 28976 27770 29028
rect 32950 28976 32956 29028
rect 33008 29016 33014 29028
rect 39850 29016 39856 29028
rect 33008 28988 39856 29016
rect 33008 28976 33014 28988
rect 39850 28976 39856 28988
rect 39908 28976 39914 29028
rect 19116 28920 19472 28948
rect 19116 28908 19122 28920
rect 34146 28908 34152 28960
rect 34204 28948 34210 28960
rect 41690 28948 41696 28960
rect 34204 28920 41696 28948
rect 34204 28908 34210 28920
rect 41690 28908 41696 28920
rect 41748 28908 41754 28960
rect 47210 28908 47216 28960
rect 47268 28948 47274 28960
rect 52730 28948 52736 28960
rect 47268 28920 52736 28948
rect 47268 28908 47274 28920
rect 52730 28908 52736 28920
rect 52788 28908 52794 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 26142 28704 26148 28756
rect 26200 28744 26206 28756
rect 41138 28744 41144 28756
rect 26200 28716 41144 28744
rect 26200 28704 26206 28716
rect 41138 28704 41144 28716
rect 41196 28704 41202 28756
rect 2866 28676 2872 28688
rect 2827 28648 2872 28676
rect 2866 28636 2872 28648
rect 2924 28636 2930 28688
rect 16298 28636 16304 28688
rect 16356 28676 16362 28688
rect 27154 28676 27160 28688
rect 16356 28648 27160 28676
rect 16356 28636 16362 28648
rect 27154 28636 27160 28648
rect 27212 28636 27218 28688
rect 35710 28636 35716 28688
rect 35768 28676 35774 28688
rect 47578 28676 47584 28688
rect 35768 28648 47584 28676
rect 35768 28636 35774 28648
rect 47578 28636 47584 28648
rect 47636 28636 47642 28688
rect 36998 28568 37004 28620
rect 37056 28608 37062 28620
rect 47946 28608 47952 28620
rect 37056 28580 47952 28608
rect 37056 28568 37062 28580
rect 47946 28568 47952 28580
rect 48004 28568 48010 28620
rect 1578 28540 1584 28552
rect 1539 28512 1584 28540
rect 1578 28500 1584 28512
rect 1636 28500 1642 28552
rect 2498 28540 2504 28552
rect 2459 28512 2504 28540
rect 2498 28500 2504 28512
rect 2556 28500 2562 28552
rect 2655 28543 2713 28549
rect 2655 28509 2667 28543
rect 2701 28540 2713 28543
rect 18230 28540 18236 28552
rect 2701 28512 18236 28540
rect 2701 28509 2713 28512
rect 2655 28503 2713 28509
rect 18230 28500 18236 28512
rect 18288 28500 18294 28552
rect 25406 28500 25412 28552
rect 25464 28540 25470 28552
rect 42886 28540 42892 28552
rect 25464 28512 42892 28540
rect 25464 28500 25470 28512
rect 42886 28500 42892 28512
rect 42944 28500 42950 28552
rect 43990 28500 43996 28552
rect 44048 28540 44054 28552
rect 57885 28543 57943 28549
rect 57885 28540 57897 28543
rect 44048 28512 57897 28540
rect 44048 28500 44054 28512
rect 57885 28509 57897 28512
rect 57931 28509 57943 28543
rect 57885 28503 57943 28509
rect 1854 28472 1860 28484
rect 1815 28444 1860 28472
rect 1854 28432 1860 28444
rect 1912 28432 1918 28484
rect 24946 28432 24952 28484
rect 25004 28472 25010 28484
rect 31846 28472 31852 28484
rect 25004 28444 31852 28472
rect 25004 28432 25010 28444
rect 31846 28432 31852 28444
rect 31904 28432 31910 28484
rect 58158 28472 58164 28484
rect 58119 28444 58164 28472
rect 58158 28432 58164 28444
rect 58216 28432 58222 28484
rect 23014 28364 23020 28416
rect 23072 28404 23078 28416
rect 54754 28404 54760 28416
rect 23072 28376 54760 28404
rect 23072 28364 23078 28376
rect 54754 28364 54760 28376
rect 54812 28364 54818 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 1578 28160 1584 28212
rect 1636 28200 1642 28212
rect 2869 28203 2927 28209
rect 2869 28200 2881 28203
rect 1636 28172 2881 28200
rect 1636 28160 1642 28172
rect 2869 28169 2881 28172
rect 2915 28169 2927 28203
rect 2869 28163 2927 28169
rect 31846 28160 31852 28212
rect 31904 28200 31910 28212
rect 44174 28200 44180 28212
rect 31904 28172 44180 28200
rect 31904 28160 31910 28172
rect 44174 28160 44180 28172
rect 44232 28160 44238 28212
rect 55306 28160 55312 28212
rect 55364 28200 55370 28212
rect 56042 28200 56048 28212
rect 55364 28172 56048 28200
rect 55364 28160 55370 28172
rect 56042 28160 56048 28172
rect 56100 28160 56106 28212
rect 2225 28135 2283 28141
rect 2225 28101 2237 28135
rect 2271 28132 2283 28135
rect 2271 28104 6914 28132
rect 2271 28101 2283 28104
rect 2225 28095 2283 28101
rect 1394 28064 1400 28076
rect 1355 28036 1400 28064
rect 1394 28024 1400 28036
rect 1452 28024 1458 28076
rect 2498 28064 2504 28076
rect 2459 28036 2504 28064
rect 2498 28024 2504 28036
rect 2556 28024 2562 28076
rect 2700 28073 2728 28104
rect 2655 28067 2728 28073
rect 2655 28033 2667 28067
rect 2701 28036 2728 28067
rect 6886 28064 6914 28104
rect 17954 28064 17960 28076
rect 6886 28036 17960 28064
rect 2701 28033 2713 28036
rect 2655 28027 2713 28033
rect 17954 28024 17960 28036
rect 18012 28024 18018 28076
rect 1578 27996 1584 28008
rect 1539 27968 1584 27996
rect 1578 27956 1584 27968
rect 1636 27956 1642 28008
rect 30374 27820 30380 27872
rect 30432 27860 30438 27872
rect 33042 27860 33048 27872
rect 30432 27832 33048 27860
rect 30432 27820 30438 27832
rect 33042 27820 33048 27832
rect 33100 27820 33106 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 1394 27616 1400 27668
rect 1452 27656 1458 27668
rect 2225 27659 2283 27665
rect 2225 27656 2237 27659
rect 1452 27628 2237 27656
rect 1452 27616 1458 27628
rect 2225 27625 2237 27628
rect 2271 27625 2283 27659
rect 2225 27619 2283 27625
rect 18046 27616 18052 27668
rect 18104 27656 18110 27668
rect 22002 27656 22008 27668
rect 18104 27628 22008 27656
rect 18104 27616 18110 27628
rect 22002 27616 22008 27628
rect 22060 27616 22066 27668
rect 44818 27616 44824 27668
rect 44876 27656 44882 27668
rect 45646 27656 45652 27668
rect 44876 27628 45652 27656
rect 44876 27616 44882 27628
rect 45646 27616 45652 27628
rect 45704 27616 45710 27668
rect 17954 27548 17960 27600
rect 18012 27588 18018 27600
rect 18874 27588 18880 27600
rect 18012 27560 18880 27588
rect 18012 27548 18018 27560
rect 18874 27548 18880 27560
rect 18932 27588 18938 27600
rect 18932 27560 19472 27588
rect 18932 27548 18938 27560
rect 18049 27523 18107 27529
rect 18049 27489 18061 27523
rect 18095 27520 18107 27523
rect 18414 27520 18420 27532
rect 18095 27492 18420 27520
rect 18095 27489 18107 27492
rect 18049 27483 18107 27489
rect 18414 27480 18420 27492
rect 18472 27480 18478 27532
rect 19334 27520 19340 27532
rect 18524 27492 19340 27520
rect 2222 27461 2228 27464
rect 2041 27455 2099 27461
rect 2041 27421 2053 27455
rect 2087 27421 2099 27455
rect 2041 27415 2099 27421
rect 2195 27455 2228 27461
rect 2195 27421 2207 27455
rect 2195 27415 2228 27421
rect 2056 27384 2084 27415
rect 2222 27412 2228 27415
rect 2280 27412 2286 27464
rect 17954 27412 17960 27464
rect 18012 27452 18018 27464
rect 18524 27461 18552 27492
rect 19334 27480 19340 27492
rect 19392 27480 19398 27532
rect 19444 27520 19472 27560
rect 20530 27548 20536 27600
rect 20588 27588 20594 27600
rect 24026 27588 24032 27600
rect 20588 27560 24032 27588
rect 20588 27548 20594 27560
rect 24026 27548 24032 27560
rect 24084 27548 24090 27600
rect 31938 27520 31944 27532
rect 19444 27492 31944 27520
rect 31938 27480 31944 27492
rect 31996 27520 32002 27532
rect 32858 27520 32864 27532
rect 31996 27492 32864 27520
rect 31996 27480 32002 27492
rect 32858 27480 32864 27492
rect 32916 27480 32922 27532
rect 35894 27480 35900 27532
rect 35952 27520 35958 27532
rect 42058 27520 42064 27532
rect 35952 27492 42064 27520
rect 35952 27480 35958 27492
rect 42058 27480 42064 27492
rect 42116 27480 42122 27532
rect 18141 27455 18199 27461
rect 18141 27452 18153 27455
rect 18012 27424 18153 27452
rect 18012 27412 18018 27424
rect 18141 27421 18153 27424
rect 18187 27421 18199 27455
rect 18141 27415 18199 27421
rect 18509 27455 18567 27461
rect 18509 27421 18521 27455
rect 18555 27421 18567 27455
rect 18782 27452 18788 27464
rect 18509 27415 18567 27421
rect 18616 27424 18788 27452
rect 18616 27396 18644 27424
rect 18782 27412 18788 27424
rect 18840 27412 18846 27464
rect 57974 27452 57980 27464
rect 57935 27424 57980 27452
rect 57974 27412 57980 27424
rect 58032 27412 58038 27464
rect 2498 27384 2504 27396
rect 2056 27356 2504 27384
rect 2498 27344 2504 27356
rect 2556 27344 2562 27396
rect 18598 27384 18604 27396
rect 18559 27356 18604 27384
rect 18598 27344 18604 27356
rect 18656 27344 18662 27396
rect 18693 27387 18751 27393
rect 18693 27353 18705 27387
rect 18739 27384 18751 27387
rect 20714 27384 20720 27396
rect 18739 27356 20720 27384
rect 18739 27353 18751 27356
rect 18693 27347 18751 27353
rect 17862 27276 17868 27328
rect 17920 27316 17926 27328
rect 18708 27316 18736 27347
rect 20714 27344 20720 27356
rect 20772 27344 20778 27396
rect 17920 27288 18736 27316
rect 17920 27276 17926 27288
rect 25314 27276 25320 27328
rect 25372 27316 25378 27328
rect 58069 27319 58127 27325
rect 58069 27316 58081 27319
rect 25372 27288 58081 27316
rect 25372 27276 25378 27288
rect 58069 27285 58081 27288
rect 58115 27285 58127 27319
rect 58069 27279 58127 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 37274 27072 37280 27124
rect 37332 27112 37338 27124
rect 39574 27112 39580 27124
rect 37332 27084 39580 27112
rect 37332 27072 37338 27084
rect 39574 27072 39580 27084
rect 39632 27072 39638 27124
rect 2869 27047 2927 27053
rect 2869 27044 2881 27047
rect 1596 27016 2881 27044
rect 1596 26985 1624 27016
rect 2869 27013 2881 27016
rect 2915 27013 2927 27047
rect 18046 27044 18052 27056
rect 18007 27016 18052 27044
rect 2869 27007 2927 27013
rect 18046 27004 18052 27016
rect 18104 27004 18110 27056
rect 18598 27044 18604 27056
rect 18432 27016 18604 27044
rect 1581 26979 1639 26985
rect 1581 26945 1593 26979
rect 1627 26945 1639 26979
rect 2498 26976 2504 26988
rect 2459 26948 2504 26976
rect 1581 26939 1639 26945
rect 2498 26936 2504 26948
rect 2556 26936 2562 26988
rect 2655 26979 2713 26985
rect 2655 26945 2667 26979
rect 2701 26976 2713 26979
rect 2701 26948 6914 26976
rect 2701 26945 2713 26948
rect 2655 26939 2713 26945
rect 1762 26908 1768 26920
rect 1723 26880 1768 26908
rect 1762 26868 1768 26880
rect 1820 26868 1826 26920
rect 6886 26772 6914 26948
rect 17862 26936 17868 26988
rect 17920 26976 17926 26988
rect 18432 26985 18460 27016
rect 18598 27004 18604 27016
rect 18656 27044 18662 27056
rect 18656 27016 20024 27044
rect 18656 27004 18662 27016
rect 17957 26979 18015 26985
rect 17957 26976 17969 26979
rect 17920 26948 17969 26976
rect 17920 26936 17926 26948
rect 17957 26945 17969 26948
rect 18003 26945 18015 26979
rect 17957 26939 18015 26945
rect 18417 26979 18475 26985
rect 18417 26945 18429 26979
rect 18463 26945 18475 26979
rect 18417 26939 18475 26945
rect 18509 26979 18567 26985
rect 18509 26945 18521 26979
rect 18555 26945 18567 26979
rect 18509 26939 18567 26945
rect 18969 26979 19027 26985
rect 18969 26945 18981 26979
rect 19015 26976 19027 26979
rect 19334 26976 19340 26988
rect 19015 26948 19340 26976
rect 19015 26945 19027 26948
rect 18969 26939 19027 26945
rect 18230 26868 18236 26920
rect 18288 26908 18294 26920
rect 18524 26908 18552 26939
rect 19334 26936 19340 26948
rect 19392 26976 19398 26988
rect 19996 26985 20024 27016
rect 35710 27004 35716 27056
rect 35768 27044 35774 27056
rect 48038 27044 48044 27056
rect 35768 27016 48044 27044
rect 35768 27004 35774 27016
rect 48038 27004 48044 27016
rect 48096 27004 48102 27056
rect 19981 26979 20039 26985
rect 19392 26948 19739 26976
rect 19392 26936 19398 26948
rect 19242 26908 19248 26920
rect 18288 26880 19248 26908
rect 18288 26868 18294 26880
rect 19242 26868 19248 26880
rect 19300 26908 19306 26920
rect 19521 26911 19579 26917
rect 19521 26908 19533 26911
rect 19300 26880 19533 26908
rect 19300 26868 19306 26880
rect 19521 26877 19533 26880
rect 19567 26877 19579 26911
rect 19521 26871 19579 26877
rect 19613 26911 19671 26917
rect 19613 26877 19625 26911
rect 19659 26877 19671 26911
rect 19711 26908 19739 26948
rect 19981 26945 19993 26979
rect 20027 26945 20039 26979
rect 19981 26939 20039 26945
rect 20073 26979 20131 26985
rect 20073 26945 20085 26979
rect 20119 26976 20131 26979
rect 20162 26976 20168 26988
rect 20119 26948 20168 26976
rect 20119 26945 20131 26948
rect 20073 26939 20131 26945
rect 20088 26908 20116 26939
rect 20162 26936 20168 26948
rect 20220 26936 20226 26988
rect 20533 26979 20591 26985
rect 20533 26945 20545 26979
rect 20579 26976 20591 26979
rect 20714 26976 20720 26988
rect 20579 26948 20720 26976
rect 20579 26945 20591 26948
rect 20533 26939 20591 26945
rect 20714 26936 20720 26948
rect 20772 26936 20778 26988
rect 24670 26936 24676 26988
rect 24728 26976 24734 26988
rect 46474 26976 46480 26988
rect 24728 26948 46480 26976
rect 24728 26936 24734 26948
rect 46474 26936 46480 26948
rect 46532 26936 46538 26988
rect 19711 26880 20116 26908
rect 19613 26871 19671 26877
rect 17586 26800 17592 26852
rect 17644 26840 17650 26852
rect 19628 26840 19656 26871
rect 26602 26868 26608 26920
rect 26660 26908 26666 26920
rect 49786 26908 49792 26920
rect 26660 26880 49792 26908
rect 26660 26868 26666 26880
rect 49786 26868 49792 26880
rect 49844 26868 49850 26920
rect 21450 26840 21456 26852
rect 17644 26812 21456 26840
rect 17644 26800 17650 26812
rect 21450 26800 21456 26812
rect 21508 26800 21514 26852
rect 22186 26772 22192 26784
rect 6886 26744 22192 26772
rect 22186 26732 22192 26744
rect 22244 26732 22250 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 58710 26500 58716 26512
rect 26344 26472 58716 26500
rect 2869 26435 2927 26441
rect 2869 26432 2881 26435
rect 1596 26404 2881 26432
rect 1596 26373 1624 26404
rect 2869 26401 2881 26404
rect 2915 26401 2927 26435
rect 18598 26432 18604 26444
rect 18559 26404 18604 26432
rect 2869 26395 2927 26401
rect 18598 26392 18604 26404
rect 18656 26392 18662 26444
rect 20162 26432 20168 26444
rect 20123 26404 20168 26432
rect 20162 26392 20168 26404
rect 20220 26392 20226 26444
rect 25866 26392 25872 26444
rect 25924 26432 25930 26444
rect 26237 26435 26295 26441
rect 26237 26432 26249 26435
rect 25924 26404 26249 26432
rect 25924 26392 25930 26404
rect 26237 26401 26249 26404
rect 26283 26401 26295 26435
rect 26237 26395 26295 26401
rect 1581 26367 1639 26373
rect 1581 26333 1593 26367
rect 1627 26333 1639 26367
rect 2498 26364 2504 26376
rect 2459 26336 2504 26364
rect 1581 26327 1639 26333
rect 2498 26324 2504 26336
rect 2556 26324 2562 26376
rect 2590 26324 2596 26376
rect 2648 26364 2654 26376
rect 18233 26367 18291 26373
rect 2648 26336 2693 26364
rect 2648 26324 2654 26336
rect 18233 26333 18245 26367
rect 18279 26364 18291 26367
rect 18322 26364 18328 26376
rect 18279 26336 18328 26364
rect 18279 26333 18291 26336
rect 18233 26327 18291 26333
rect 18322 26324 18328 26336
rect 18380 26324 18386 26376
rect 19426 26364 19432 26376
rect 19339 26336 19432 26364
rect 19426 26324 19432 26336
rect 19484 26364 19490 26376
rect 20070 26364 20076 26376
rect 19484 26336 20076 26364
rect 19484 26324 19490 26336
rect 20070 26324 20076 26336
rect 20128 26324 20134 26376
rect 25409 26367 25467 26373
rect 25409 26333 25421 26367
rect 25455 26364 25467 26367
rect 26053 26367 26111 26373
rect 26053 26364 26065 26367
rect 25455 26336 26065 26364
rect 25455 26333 25467 26336
rect 25409 26327 25467 26333
rect 26053 26333 26065 26336
rect 26099 26364 26111 26367
rect 26344 26364 26372 26472
rect 58710 26460 58716 26472
rect 58768 26460 58774 26512
rect 28350 26432 28356 26444
rect 27172 26404 28356 26432
rect 27172 26373 27200 26404
rect 28350 26392 28356 26404
rect 28408 26392 28414 26444
rect 58158 26432 58164 26444
rect 58119 26404 58164 26432
rect 58158 26392 58164 26404
rect 58216 26392 58222 26444
rect 26099 26336 26372 26364
rect 27157 26367 27215 26373
rect 26099 26333 26111 26336
rect 26053 26327 26111 26333
rect 27157 26333 27169 26367
rect 27203 26333 27215 26367
rect 27157 26327 27215 26333
rect 27249 26367 27307 26373
rect 27249 26333 27261 26367
rect 27295 26333 27307 26367
rect 27249 26327 27307 26333
rect 1854 26296 1860 26308
rect 1815 26268 1860 26296
rect 1854 26256 1860 26268
rect 1912 26256 1918 26308
rect 26142 26296 26148 26308
rect 26103 26268 26148 26296
rect 26142 26256 26148 26268
rect 26200 26256 26206 26308
rect 26786 26256 26792 26308
rect 26844 26296 26850 26308
rect 27264 26296 27292 26327
rect 40402 26324 40408 26376
rect 40460 26364 40466 26376
rect 57885 26367 57943 26373
rect 57885 26364 57897 26367
rect 40460 26336 57897 26364
rect 40460 26324 40466 26336
rect 57885 26333 57897 26336
rect 57931 26333 57943 26367
rect 57885 26327 57943 26333
rect 27430 26296 27436 26308
rect 26844 26268 27292 26296
rect 27391 26268 27436 26296
rect 26844 26256 26850 26268
rect 27430 26256 27436 26268
rect 27488 26256 27494 26308
rect 25682 26228 25688 26240
rect 25643 26200 25688 26228
rect 25682 26188 25688 26200
rect 25740 26188 25746 26240
rect 26878 26188 26884 26240
rect 26936 26228 26942 26240
rect 58342 26228 58348 26240
rect 26936 26200 58348 26228
rect 26936 26188 26942 26200
rect 58342 26188 58348 26200
rect 58400 26188 58406 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 23382 25984 23388 26036
rect 23440 26024 23446 26036
rect 24854 26024 24860 26036
rect 23440 25996 24860 26024
rect 23440 25984 23446 25996
rect 24854 25984 24860 25996
rect 24912 26024 24918 26036
rect 28261 26027 28319 26033
rect 28261 26024 28273 26027
rect 24912 25996 28273 26024
rect 24912 25984 24918 25996
rect 28261 25993 28273 25996
rect 28307 25993 28319 26027
rect 28261 25987 28319 25993
rect 25866 25916 25872 25968
rect 25924 25956 25930 25968
rect 28353 25959 28411 25965
rect 25924 25928 26096 25956
rect 25924 25916 25930 25928
rect 1581 25891 1639 25897
rect 1581 25857 1593 25891
rect 1627 25888 1639 25891
rect 2682 25888 2688 25900
rect 1627 25860 2688 25888
rect 1627 25857 1639 25860
rect 1581 25851 1639 25857
rect 2682 25848 2688 25860
rect 2740 25848 2746 25900
rect 19889 25891 19947 25897
rect 19889 25857 19901 25891
rect 19935 25888 19947 25891
rect 20530 25888 20536 25900
rect 19935 25860 20536 25888
rect 19935 25857 19947 25860
rect 19889 25851 19947 25857
rect 20530 25848 20536 25860
rect 20588 25848 20594 25900
rect 20625 25891 20683 25897
rect 20625 25857 20637 25891
rect 20671 25888 20683 25891
rect 21082 25888 21088 25900
rect 20671 25860 21088 25888
rect 20671 25857 20683 25860
rect 20625 25851 20683 25857
rect 21082 25848 21088 25860
rect 21140 25848 21146 25900
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25857 26019 25891
rect 26068 25888 26096 25928
rect 28353 25925 28365 25959
rect 28399 25956 28411 25959
rect 28442 25956 28448 25968
rect 28399 25928 28448 25956
rect 28399 25925 28411 25928
rect 28353 25919 28411 25925
rect 28442 25916 28448 25928
rect 28500 25916 28506 25968
rect 29273 25959 29331 25965
rect 29273 25925 29285 25959
rect 29319 25956 29331 25959
rect 29822 25956 29828 25968
rect 29319 25928 29828 25956
rect 29319 25925 29331 25928
rect 29273 25919 29331 25925
rect 29822 25916 29828 25928
rect 29880 25916 29886 25968
rect 26068 25860 26280 25888
rect 25961 25851 26019 25857
rect 1762 25820 1768 25832
rect 1723 25792 1768 25820
rect 1762 25780 1768 25792
rect 1820 25780 1826 25832
rect 20438 25780 20444 25832
rect 20496 25820 20502 25832
rect 20717 25823 20775 25829
rect 20717 25820 20729 25823
rect 20496 25792 20729 25820
rect 20496 25780 20502 25792
rect 20717 25789 20729 25792
rect 20763 25820 20775 25823
rect 25866 25820 25872 25832
rect 20763 25792 25872 25820
rect 20763 25789 20775 25792
rect 20717 25783 20775 25789
rect 25866 25780 25872 25792
rect 25924 25780 25930 25832
rect 25317 25755 25375 25761
rect 25317 25721 25329 25755
rect 25363 25752 25375 25755
rect 25976 25752 26004 25851
rect 26050 25780 26056 25832
rect 26108 25820 26114 25832
rect 26252 25829 26280 25860
rect 27982 25848 27988 25900
rect 28040 25888 28046 25900
rect 29457 25891 29515 25897
rect 29457 25888 29469 25891
rect 28040 25860 29469 25888
rect 28040 25848 28046 25860
rect 29457 25857 29469 25860
rect 29503 25857 29515 25891
rect 58066 25888 58072 25900
rect 58027 25860 58072 25888
rect 29457 25851 29515 25857
rect 58066 25848 58072 25860
rect 58124 25848 58130 25900
rect 26237 25823 26295 25829
rect 26108 25792 26153 25820
rect 26108 25780 26114 25792
rect 26237 25789 26249 25823
rect 26283 25789 26295 25823
rect 26237 25783 26295 25789
rect 28261 25823 28319 25829
rect 28261 25789 28273 25823
rect 28307 25820 28319 25823
rect 29086 25820 29092 25832
rect 28307 25792 29092 25820
rect 28307 25789 28319 25792
rect 28261 25783 28319 25789
rect 29086 25780 29092 25792
rect 29144 25780 29150 25832
rect 58434 25752 58440 25764
rect 25363 25724 58440 25752
rect 25363 25721 25375 25724
rect 25317 25715 25375 25721
rect 58434 25712 58440 25724
rect 58492 25712 58498 25764
rect 20070 25644 20076 25696
rect 20128 25684 20134 25696
rect 20165 25687 20223 25693
rect 20165 25684 20177 25687
rect 20128 25656 20177 25684
rect 20128 25644 20134 25656
rect 20165 25653 20177 25656
rect 20211 25653 20223 25687
rect 25590 25684 25596 25696
rect 25551 25656 25596 25684
rect 20165 25647 20223 25653
rect 25590 25644 25596 25656
rect 25648 25644 25654 25696
rect 27798 25684 27804 25696
rect 27759 25656 27804 25684
rect 27798 25644 27804 25656
rect 27856 25644 27862 25696
rect 29641 25687 29699 25693
rect 29641 25653 29653 25687
rect 29687 25684 29699 25687
rect 31570 25684 31576 25696
rect 29687 25656 31576 25684
rect 29687 25653 29699 25656
rect 29641 25647 29699 25653
rect 31570 25644 31576 25656
rect 31628 25644 31634 25696
rect 58250 25684 58256 25696
rect 58211 25656 58256 25684
rect 58250 25644 58256 25656
rect 58308 25644 58314 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 2682 25480 2688 25492
rect 2643 25452 2688 25480
rect 2682 25440 2688 25452
rect 2740 25440 2746 25492
rect 19242 25440 19248 25492
rect 19300 25480 19306 25492
rect 19978 25480 19984 25492
rect 19300 25452 19984 25480
rect 19300 25440 19306 25452
rect 19978 25440 19984 25452
rect 20036 25440 20042 25492
rect 26878 25480 26884 25492
rect 22066 25452 26884 25480
rect 2498 25372 2504 25424
rect 2556 25372 2562 25424
rect 2516 25344 2544 25372
rect 15194 25344 15200 25356
rect 2516 25316 15200 25344
rect 1578 25276 1584 25288
rect 1539 25248 1584 25276
rect 1578 25236 1584 25248
rect 1636 25236 1642 25288
rect 2516 25285 2544 25316
rect 15194 25304 15200 25316
rect 15252 25304 15258 25356
rect 16482 25344 16488 25356
rect 16443 25316 16488 25344
rect 16482 25304 16488 25316
rect 16540 25304 16546 25356
rect 20438 25304 20444 25356
rect 20496 25344 20502 25356
rect 21913 25347 21971 25353
rect 21913 25344 21925 25347
rect 20496 25316 21925 25344
rect 20496 25304 20502 25316
rect 21913 25313 21925 25316
rect 21959 25313 21971 25347
rect 21913 25307 21971 25313
rect 2501 25279 2559 25285
rect 2501 25245 2513 25279
rect 2547 25245 2559 25279
rect 2501 25239 2559 25245
rect 2655 25279 2713 25285
rect 2655 25245 2667 25279
rect 2701 25276 2713 25279
rect 16117 25279 16175 25285
rect 2701 25248 9674 25276
rect 2701 25245 2713 25248
rect 2655 25239 2713 25245
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 9646 25140 9674 25248
rect 16117 25245 16129 25279
rect 16163 25276 16175 25279
rect 17218 25276 17224 25288
rect 16163 25248 17224 25276
rect 16163 25245 16175 25248
rect 16117 25239 16175 25245
rect 17218 25236 17224 25248
rect 17276 25236 17282 25288
rect 19337 25279 19395 25285
rect 19337 25245 19349 25279
rect 19383 25276 19395 25279
rect 20162 25276 20168 25288
rect 19383 25248 20168 25276
rect 19383 25245 19395 25248
rect 19337 25239 19395 25245
rect 20162 25236 20168 25248
rect 20220 25236 20226 25288
rect 21085 25279 21143 25285
rect 21085 25245 21097 25279
rect 21131 25276 21143 25279
rect 21729 25279 21787 25285
rect 21729 25276 21741 25279
rect 21131 25248 21741 25276
rect 21131 25245 21143 25248
rect 21085 25239 21143 25245
rect 21729 25245 21741 25248
rect 21775 25276 21787 25279
rect 22066 25276 22094 25452
rect 26878 25440 26884 25452
rect 26936 25440 26942 25492
rect 27798 25440 27804 25492
rect 27856 25480 27862 25492
rect 55490 25480 55496 25492
rect 27856 25452 55496 25480
rect 27856 25440 27862 25452
rect 55490 25440 55496 25452
rect 55548 25440 55554 25492
rect 55582 25440 55588 25492
rect 55640 25480 55646 25492
rect 58894 25480 58900 25492
rect 55640 25452 58900 25480
rect 55640 25440 55646 25452
rect 58894 25440 58900 25452
rect 58952 25440 58958 25492
rect 36630 25372 36636 25424
rect 36688 25412 36694 25424
rect 58250 25412 58256 25424
rect 36688 25384 58256 25412
rect 36688 25372 36694 25384
rect 58250 25372 58256 25384
rect 58308 25372 58314 25424
rect 29089 25347 29147 25353
rect 29089 25313 29101 25347
rect 29135 25344 29147 25347
rect 30190 25344 30196 25356
rect 29135 25316 30196 25344
rect 29135 25313 29147 25316
rect 29089 25307 29147 25313
rect 30190 25304 30196 25316
rect 30248 25304 30254 25356
rect 56689 25347 56747 25353
rect 56689 25344 56701 25347
rect 55876 25316 56701 25344
rect 24946 25276 24952 25288
rect 21775 25248 22094 25276
rect 24859 25248 24952 25276
rect 21775 25245 21787 25248
rect 21729 25239 21787 25245
rect 24946 25236 24952 25248
rect 25004 25276 25010 25288
rect 27157 25279 27215 25285
rect 27157 25276 27169 25279
rect 25004 25248 27169 25276
rect 25004 25236 25010 25248
rect 27157 25245 27169 25248
rect 27203 25276 27215 25279
rect 28994 25276 29000 25288
rect 27203 25248 27568 25276
rect 28955 25248 29000 25276
rect 27203 25245 27215 25248
rect 27157 25239 27215 25245
rect 27540 25220 27568 25248
rect 28994 25236 29000 25248
rect 29052 25236 29058 25288
rect 29181 25279 29239 25285
rect 29181 25245 29193 25279
rect 29227 25276 29239 25279
rect 29454 25276 29460 25288
rect 29227 25248 29460 25276
rect 29227 25245 29239 25248
rect 29181 25239 29239 25245
rect 29454 25236 29460 25248
rect 29512 25236 29518 25288
rect 29733 25279 29791 25285
rect 29733 25245 29745 25279
rect 29779 25276 29791 25279
rect 29822 25276 29828 25288
rect 29779 25248 29828 25276
rect 29779 25245 29791 25248
rect 29733 25239 29791 25245
rect 29822 25236 29828 25248
rect 29880 25236 29886 25288
rect 55766 25236 55772 25288
rect 55824 25276 55830 25288
rect 55876 25285 55904 25316
rect 56689 25313 56701 25316
rect 56735 25313 56747 25347
rect 56689 25307 56747 25313
rect 55861 25279 55919 25285
rect 55861 25276 55873 25279
rect 55824 25248 55873 25276
rect 55824 25236 55830 25248
rect 55861 25245 55873 25248
rect 55907 25245 55919 25279
rect 56042 25276 56048 25288
rect 56003 25248 56048 25276
rect 55861 25239 55919 25245
rect 56042 25236 56048 25248
rect 56100 25236 56106 25288
rect 56870 25276 56876 25288
rect 56831 25248 56876 25276
rect 56870 25236 56876 25248
rect 56928 25236 56934 25288
rect 57885 25279 57943 25285
rect 57885 25245 57897 25279
rect 57931 25245 57943 25279
rect 57885 25239 57943 25245
rect 19604 25211 19662 25217
rect 19604 25177 19616 25211
rect 19650 25208 19662 25211
rect 19978 25208 19984 25220
rect 19650 25180 19984 25208
rect 19650 25177 19662 25180
rect 19604 25171 19662 25177
rect 19978 25168 19984 25180
rect 20036 25168 20042 25220
rect 21266 25168 21272 25220
rect 21324 25208 21330 25220
rect 21821 25211 21879 25217
rect 21821 25208 21833 25211
rect 21324 25180 21833 25208
rect 21324 25168 21330 25180
rect 21821 25177 21833 25180
rect 21867 25177 21879 25211
rect 21821 25171 21879 25177
rect 25216 25211 25274 25217
rect 25216 25177 25228 25211
rect 25262 25208 25274 25211
rect 25682 25208 25688 25220
rect 25262 25180 25688 25208
rect 25262 25177 25274 25180
rect 25216 25171 25274 25177
rect 25682 25168 25688 25180
rect 25740 25168 25746 25220
rect 26234 25168 26240 25220
rect 26292 25208 26298 25220
rect 27402 25211 27460 25217
rect 27402 25208 27414 25211
rect 26292 25180 27414 25208
rect 26292 25168 26298 25180
rect 27402 25177 27414 25180
rect 27448 25177 27460 25211
rect 27402 25171 27460 25177
rect 27522 25168 27528 25220
rect 27580 25168 27586 25220
rect 29086 25168 29092 25220
rect 29144 25208 29150 25220
rect 29917 25211 29975 25217
rect 29917 25208 29929 25211
rect 29144 25180 29929 25208
rect 29144 25168 29150 25180
rect 29917 25177 29929 25180
rect 29963 25177 29975 25211
rect 29917 25171 29975 25177
rect 53834 25168 53840 25220
rect 53892 25208 53898 25220
rect 57900 25208 57928 25239
rect 58158 25208 58164 25220
rect 53892 25180 57928 25208
rect 58119 25180 58164 25208
rect 53892 25168 53898 25180
rect 58158 25168 58164 25180
rect 58216 25168 58222 25220
rect 19242 25140 19248 25152
rect 9646 25112 19248 25140
rect 19242 25100 19248 25112
rect 19300 25100 19306 25152
rect 20622 25100 20628 25152
rect 20680 25140 20686 25152
rect 20717 25143 20775 25149
rect 20717 25140 20729 25143
rect 20680 25112 20729 25140
rect 20680 25100 20686 25112
rect 20717 25109 20729 25112
rect 20763 25109 20775 25143
rect 21358 25140 21364 25152
rect 21319 25112 21364 25140
rect 20717 25103 20775 25109
rect 21358 25100 21364 25112
rect 21416 25100 21422 25152
rect 22830 25100 22836 25152
rect 22888 25140 22894 25152
rect 26142 25140 26148 25152
rect 22888 25112 26148 25140
rect 22888 25100 22894 25112
rect 26142 25100 26148 25112
rect 26200 25140 26206 25152
rect 26329 25143 26387 25149
rect 26329 25140 26341 25143
rect 26200 25112 26341 25140
rect 26200 25100 26206 25112
rect 26329 25109 26341 25112
rect 26375 25109 26387 25143
rect 28534 25140 28540 25152
rect 28495 25112 28540 25140
rect 26329 25103 26387 25109
rect 28534 25100 28540 25112
rect 28592 25100 28598 25152
rect 30098 25140 30104 25152
rect 30059 25112 30104 25140
rect 30098 25100 30104 25112
rect 30156 25100 30162 25152
rect 56229 25143 56287 25149
rect 56229 25109 56241 25143
rect 56275 25140 56287 25143
rect 56318 25140 56324 25152
rect 56275 25112 56324 25140
rect 56275 25109 56287 25112
rect 56229 25103 56287 25109
rect 56318 25100 56324 25112
rect 56376 25100 56382 25152
rect 57057 25143 57115 25149
rect 57057 25109 57069 25143
rect 57103 25140 57115 25143
rect 57146 25140 57152 25152
rect 57103 25112 57152 25140
rect 57103 25109 57115 25112
rect 57057 25103 57115 25109
rect 57146 25100 57152 25112
rect 57204 25100 57210 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 1578 24896 1584 24948
rect 1636 24936 1642 24948
rect 16209 24939 16267 24945
rect 16209 24936 16221 24939
rect 1636 24908 16221 24936
rect 1636 24896 1642 24908
rect 16209 24905 16221 24908
rect 16255 24905 16267 24939
rect 20346 24936 20352 24948
rect 16209 24899 16267 24905
rect 19628 24908 20352 24936
rect 15194 24760 15200 24812
rect 15252 24800 15258 24812
rect 15562 24800 15568 24812
rect 15252 24772 15568 24800
rect 15252 24760 15258 24772
rect 15562 24760 15568 24772
rect 15620 24800 15626 24812
rect 15841 24803 15899 24809
rect 15841 24800 15853 24803
rect 15620 24772 15853 24800
rect 15620 24760 15626 24772
rect 15841 24769 15853 24772
rect 15887 24769 15899 24803
rect 15841 24763 15899 24769
rect 15995 24803 16053 24809
rect 15995 24769 16007 24803
rect 16041 24800 16053 24803
rect 16114 24800 16120 24812
rect 16041 24772 16120 24800
rect 16041 24769 16053 24772
rect 15995 24763 16053 24769
rect 16114 24760 16120 24772
rect 16172 24800 16178 24812
rect 16482 24800 16488 24812
rect 16172 24772 16488 24800
rect 16172 24760 16178 24772
rect 16482 24760 16488 24772
rect 16540 24760 16546 24812
rect 19334 24800 19340 24812
rect 19295 24772 19340 24800
rect 19334 24760 19340 24772
rect 19392 24760 19398 24812
rect 19628 24809 19656 24908
rect 20346 24896 20352 24908
rect 20404 24896 20410 24948
rect 20530 24896 20536 24948
rect 20588 24936 20594 24948
rect 56042 24936 56048 24948
rect 20588 24908 41414 24936
rect 56003 24908 56048 24936
rect 20588 24896 20594 24908
rect 22296 24840 22600 24868
rect 19521 24803 19579 24809
rect 19521 24769 19533 24803
rect 19567 24769 19579 24803
rect 19521 24763 19579 24769
rect 19613 24803 19671 24809
rect 19613 24769 19625 24803
rect 19659 24769 19671 24803
rect 19613 24763 19671 24769
rect 20073 24803 20131 24809
rect 20073 24769 20085 24803
rect 20119 24800 20131 24803
rect 20162 24800 20168 24812
rect 20119 24772 20168 24800
rect 20119 24769 20131 24772
rect 20073 24763 20131 24769
rect 19536 24732 19564 24763
rect 20162 24760 20168 24772
rect 20220 24760 20226 24812
rect 20340 24803 20398 24809
rect 20340 24769 20352 24803
rect 20386 24800 20398 24803
rect 21358 24800 21364 24812
rect 20386 24772 21364 24800
rect 20386 24769 20398 24772
rect 20340 24763 20398 24769
rect 21358 24760 21364 24772
rect 21416 24760 21422 24812
rect 22296 24800 22324 24840
rect 22462 24800 22468 24812
rect 22066 24772 22324 24800
rect 22423 24772 22468 24800
rect 19702 24732 19708 24744
rect 19536 24704 19708 24732
rect 19702 24692 19708 24704
rect 19760 24692 19766 24744
rect 22066 24664 22094 24772
rect 22462 24760 22468 24772
rect 22520 24760 22526 24812
rect 22572 24800 22600 24840
rect 26528 24840 28120 24868
rect 23566 24800 23572 24812
rect 22572 24772 23336 24800
rect 23527 24772 23572 24800
rect 22281 24735 22339 24741
rect 22281 24701 22293 24735
rect 22327 24732 22339 24735
rect 23198 24732 23204 24744
rect 22327 24704 23204 24732
rect 22327 24701 22339 24704
rect 22281 24695 22339 24701
rect 23198 24692 23204 24704
rect 23256 24692 23262 24744
rect 23308 24732 23336 24772
rect 23566 24760 23572 24772
rect 23624 24760 23630 24812
rect 26418 24800 26424 24812
rect 26379 24772 26424 24800
rect 26418 24760 26424 24772
rect 26476 24760 26482 24812
rect 23934 24732 23940 24744
rect 23308 24704 23940 24732
rect 23934 24692 23940 24704
rect 23992 24732 23998 24744
rect 26528 24732 26556 24840
rect 26605 24803 26663 24809
rect 26605 24769 26617 24803
rect 26651 24769 26663 24803
rect 26605 24763 26663 24769
rect 23992 24704 26556 24732
rect 23992 24692 23998 24704
rect 21008 24636 22094 24664
rect 19150 24556 19156 24608
rect 19208 24596 19214 24608
rect 19337 24599 19395 24605
rect 19337 24596 19349 24599
rect 19208 24568 19349 24596
rect 19208 24556 19214 24568
rect 19337 24565 19349 24568
rect 19383 24565 19395 24599
rect 19337 24559 19395 24565
rect 19426 24556 19432 24608
rect 19484 24596 19490 24608
rect 21008 24596 21036 24636
rect 22554 24624 22560 24676
rect 22612 24664 22618 24676
rect 24210 24664 24216 24676
rect 22612 24636 24216 24664
rect 22612 24624 22618 24636
rect 24210 24624 24216 24636
rect 24268 24624 24274 24676
rect 24302 24624 24308 24676
rect 24360 24664 24366 24676
rect 26620 24664 26648 24763
rect 27246 24760 27252 24812
rect 27304 24800 27310 24812
rect 27965 24803 28023 24809
rect 27965 24800 27977 24803
rect 27304 24772 27977 24800
rect 27304 24760 27310 24772
rect 27965 24769 27977 24772
rect 28011 24769 28023 24803
rect 28092 24800 28120 24840
rect 29914 24828 29920 24880
rect 29972 24868 29978 24880
rect 31386 24868 31392 24880
rect 29972 24840 31392 24868
rect 29972 24828 29978 24840
rect 31386 24828 31392 24840
rect 31444 24828 31450 24880
rect 31757 24871 31815 24877
rect 31757 24837 31769 24871
rect 31803 24868 31815 24871
rect 41386 24868 41414 24908
rect 56042 24896 56048 24908
rect 56100 24896 56106 24948
rect 56870 24896 56876 24948
rect 56928 24936 56934 24948
rect 57057 24939 57115 24945
rect 57057 24936 57069 24939
rect 56928 24908 57069 24936
rect 56928 24896 56934 24908
rect 57057 24905 57069 24908
rect 57103 24905 57115 24939
rect 57057 24899 57115 24905
rect 55582 24868 55588 24880
rect 31803 24840 32812 24868
rect 41386 24840 55588 24868
rect 31803 24837 31815 24840
rect 31757 24831 31815 24837
rect 29822 24809 29828 24812
rect 28092 24772 28764 24800
rect 27965 24763 28023 24769
rect 27614 24692 27620 24744
rect 27672 24732 27678 24744
rect 27709 24735 27767 24741
rect 27709 24732 27721 24735
rect 27672 24704 27721 24732
rect 27672 24692 27678 24704
rect 27709 24701 27721 24704
rect 27755 24701 27767 24735
rect 27709 24695 27767 24701
rect 24360 24636 27660 24664
rect 24360 24624 24366 24636
rect 27632 24608 27660 24636
rect 19484 24568 21036 24596
rect 19484 24556 19490 24568
rect 21266 24556 21272 24608
rect 21324 24596 21330 24608
rect 21453 24599 21511 24605
rect 21453 24596 21465 24599
rect 21324 24568 21465 24596
rect 21324 24556 21330 24568
rect 21453 24565 21465 24568
rect 21499 24565 21511 24599
rect 21453 24559 21511 24565
rect 22649 24599 22707 24605
rect 22649 24565 22661 24599
rect 22695 24596 22707 24599
rect 22738 24596 22744 24608
rect 22695 24568 22744 24596
rect 22695 24565 22707 24568
rect 22649 24559 22707 24565
rect 22738 24556 22744 24568
rect 22796 24556 22802 24608
rect 24670 24556 24676 24608
rect 24728 24596 24734 24608
rect 24765 24599 24823 24605
rect 24765 24596 24777 24599
rect 24728 24568 24777 24596
rect 24728 24556 24734 24568
rect 24765 24565 24777 24568
rect 24811 24565 24823 24599
rect 24765 24559 24823 24565
rect 26050 24556 26056 24608
rect 26108 24596 26114 24608
rect 26513 24599 26571 24605
rect 26513 24596 26525 24599
rect 26108 24568 26525 24596
rect 26108 24556 26114 24568
rect 26513 24565 26525 24568
rect 26559 24565 26571 24599
rect 26513 24559 26571 24565
rect 27614 24556 27620 24608
rect 27672 24556 27678 24608
rect 27724 24596 27752 24695
rect 28736 24664 28764 24772
rect 29816 24763 29828 24809
rect 29880 24800 29886 24812
rect 31573 24803 31631 24809
rect 29880 24772 29916 24800
rect 29822 24760 29828 24763
rect 29880 24760 29886 24772
rect 31573 24769 31585 24803
rect 31619 24769 31631 24803
rect 32582 24800 32588 24812
rect 32543 24772 32588 24800
rect 31573 24763 31631 24769
rect 28902 24692 28908 24744
rect 28960 24732 28966 24744
rect 29549 24735 29607 24741
rect 29549 24732 29561 24735
rect 28960 24704 29561 24732
rect 28960 24692 28966 24704
rect 29549 24701 29561 24704
rect 29595 24701 29607 24735
rect 31588 24732 31616 24763
rect 32582 24760 32588 24772
rect 32640 24760 32646 24812
rect 32784 24809 32812 24840
rect 55582 24828 55588 24840
rect 55640 24828 55646 24880
rect 56781 24871 56839 24877
rect 55876 24840 56088 24868
rect 32677 24803 32735 24809
rect 32677 24769 32689 24803
rect 32723 24769 32735 24803
rect 32677 24763 32735 24769
rect 32769 24803 32827 24809
rect 32769 24769 32781 24803
rect 32815 24769 32827 24803
rect 32769 24763 32827 24769
rect 31662 24732 31668 24744
rect 31588 24704 31668 24732
rect 29549 24695 29607 24701
rect 31662 24692 31668 24704
rect 31720 24692 31726 24744
rect 31846 24692 31852 24744
rect 31904 24732 31910 24744
rect 32692 24732 32720 24763
rect 32858 24760 32864 24812
rect 32916 24800 32922 24812
rect 32953 24803 33011 24809
rect 32953 24800 32965 24803
rect 32916 24772 32965 24800
rect 32916 24760 32922 24772
rect 32953 24769 32965 24772
rect 32999 24800 33011 24803
rect 36078 24800 36084 24812
rect 32999 24772 36084 24800
rect 32999 24769 33011 24772
rect 32953 24763 33011 24769
rect 36078 24760 36084 24772
rect 36136 24760 36142 24812
rect 36998 24760 37004 24812
rect 37056 24800 37062 24812
rect 45278 24800 45284 24812
rect 37056 24772 45284 24800
rect 37056 24760 37062 24772
rect 45278 24760 45284 24772
rect 45336 24760 45342 24812
rect 45462 24800 45468 24812
rect 45423 24772 45468 24800
rect 45462 24760 45468 24772
rect 45520 24760 45526 24812
rect 45833 24803 45891 24809
rect 45833 24769 45845 24803
rect 45879 24800 45891 24803
rect 51166 24800 51172 24812
rect 45879 24772 51172 24800
rect 45879 24769 45891 24772
rect 45833 24763 45891 24769
rect 51166 24760 51172 24772
rect 51224 24760 51230 24812
rect 54297 24803 54355 24809
rect 54297 24769 54309 24803
rect 54343 24800 54355 24803
rect 55306 24800 55312 24812
rect 54343 24772 55312 24800
rect 54343 24769 54355 24772
rect 54297 24763 54355 24769
rect 55306 24760 55312 24772
rect 55364 24760 55370 24812
rect 55490 24800 55496 24812
rect 55451 24772 55496 24800
rect 55490 24760 55496 24772
rect 55548 24760 55554 24812
rect 55876 24809 55904 24840
rect 55677 24803 55735 24809
rect 55677 24769 55689 24803
rect 55723 24769 55735 24803
rect 55677 24763 55735 24769
rect 55769 24803 55827 24809
rect 55769 24769 55781 24803
rect 55815 24769 55827 24803
rect 55769 24763 55827 24769
rect 55861 24803 55919 24809
rect 55861 24769 55873 24803
rect 55907 24769 55919 24803
rect 56060 24800 56088 24840
rect 56781 24837 56793 24871
rect 56827 24868 56839 24871
rect 56827 24840 57008 24868
rect 56827 24837 56839 24840
rect 56781 24831 56839 24837
rect 56226 24800 56232 24812
rect 56060 24772 56232 24800
rect 55861 24763 55919 24769
rect 31904 24704 32720 24732
rect 31904 24692 31910 24704
rect 33042 24692 33048 24744
rect 33100 24732 33106 24744
rect 45373 24735 45431 24741
rect 45373 24732 45385 24735
rect 33100 24704 45385 24732
rect 33100 24692 33106 24704
rect 45373 24701 45385 24704
rect 45419 24701 45431 24735
rect 45373 24695 45431 24701
rect 45738 24692 45744 24744
rect 45796 24732 45802 24744
rect 45925 24735 45983 24741
rect 45925 24732 45937 24735
rect 45796 24704 45937 24732
rect 45796 24692 45802 24704
rect 45925 24701 45937 24704
rect 45971 24701 45983 24735
rect 51810 24732 51816 24744
rect 45925 24695 45983 24701
rect 46308 24704 51816 24732
rect 28736 24636 29224 24664
rect 28902 24596 28908 24608
rect 27724 24568 28908 24596
rect 28902 24556 28908 24568
rect 28960 24556 28966 24608
rect 29086 24596 29092 24608
rect 29047 24568 29092 24596
rect 29086 24556 29092 24568
rect 29144 24556 29150 24608
rect 29196 24596 29224 24636
rect 32582 24624 32588 24676
rect 32640 24664 32646 24676
rect 33229 24667 33287 24673
rect 33229 24664 33241 24667
rect 32640 24636 33241 24664
rect 32640 24624 32646 24636
rect 33229 24633 33241 24636
rect 33275 24664 33287 24667
rect 46198 24664 46204 24676
rect 33275 24636 38654 24664
rect 33275 24633 33287 24636
rect 33229 24627 33287 24633
rect 30466 24596 30472 24608
rect 29196 24568 30472 24596
rect 30466 24556 30472 24568
rect 30524 24556 30530 24608
rect 30834 24556 30840 24608
rect 30892 24596 30898 24608
rect 30929 24599 30987 24605
rect 30929 24596 30941 24599
rect 30892 24568 30941 24596
rect 30892 24556 30898 24568
rect 30929 24565 30941 24568
rect 30975 24565 30987 24599
rect 32306 24596 32312 24608
rect 32267 24568 32312 24596
rect 30929 24559 30987 24565
rect 32306 24556 32312 24568
rect 32364 24556 32370 24608
rect 38626 24596 38654 24636
rect 41386 24636 46204 24664
rect 41386 24596 41414 24636
rect 46198 24624 46204 24636
rect 46256 24624 46262 24676
rect 38626 24568 41414 24596
rect 44913 24599 44971 24605
rect 44913 24565 44925 24599
rect 44959 24596 44971 24599
rect 45002 24596 45008 24608
rect 44959 24568 45008 24596
rect 44959 24565 44971 24568
rect 44913 24559 44971 24565
rect 45002 24556 45008 24568
rect 45060 24556 45066 24608
rect 45278 24556 45284 24608
rect 45336 24596 45342 24608
rect 46308 24596 46336 24704
rect 51810 24692 51816 24704
rect 51868 24732 51874 24744
rect 54110 24732 54116 24744
rect 51868 24704 54116 24732
rect 51868 24692 51874 24704
rect 54110 24692 54116 24704
rect 54168 24732 54174 24744
rect 54573 24735 54631 24741
rect 54573 24732 54585 24735
rect 54168 24704 54585 24732
rect 54168 24692 54174 24704
rect 54573 24701 54585 24704
rect 54619 24701 54631 24735
rect 54573 24695 54631 24701
rect 55122 24692 55128 24744
rect 55180 24732 55186 24744
rect 55692 24732 55720 24763
rect 55180 24704 55720 24732
rect 55784 24732 55812 24763
rect 56226 24760 56232 24772
rect 56284 24760 56290 24812
rect 56502 24760 56508 24812
rect 56560 24800 56566 24812
rect 56560 24772 56605 24800
rect 56560 24760 56566 24772
rect 56686 24760 56692 24812
rect 56744 24800 56750 24812
rect 56870 24800 56876 24812
rect 56744 24772 56789 24800
rect 56831 24772 56876 24800
rect 56744 24760 56750 24772
rect 56870 24760 56876 24772
rect 56928 24760 56934 24812
rect 56980 24800 57008 24840
rect 58066 24800 58072 24812
rect 56980 24772 57836 24800
rect 58027 24772 58072 24800
rect 57422 24732 57428 24744
rect 55784 24704 57428 24732
rect 55180 24692 55186 24704
rect 46382 24624 46388 24676
rect 46440 24664 46446 24676
rect 55030 24664 55036 24676
rect 46440 24636 55036 24664
rect 46440 24624 46446 24636
rect 55030 24624 55036 24636
rect 55088 24624 55094 24676
rect 55692 24664 55720 24704
rect 57422 24692 57428 24704
rect 57480 24692 57486 24744
rect 57808 24732 57836 24772
rect 58066 24760 58072 24772
rect 58124 24760 58130 24812
rect 58342 24732 58348 24744
rect 57808 24704 58348 24732
rect 58342 24692 58348 24704
rect 58400 24692 58406 24744
rect 55692 24636 56180 24664
rect 45336 24568 46336 24596
rect 45336 24556 45342 24568
rect 50062 24556 50068 24608
rect 50120 24596 50126 24608
rect 54478 24596 54484 24608
rect 50120 24568 54484 24596
rect 50120 24556 50126 24568
rect 54478 24556 54484 24568
rect 54536 24596 54542 24608
rect 55766 24596 55772 24608
rect 54536 24568 55772 24596
rect 54536 24556 54542 24568
rect 55766 24556 55772 24568
rect 55824 24556 55830 24608
rect 56152 24596 56180 24636
rect 56226 24624 56232 24676
rect 56284 24664 56290 24676
rect 56870 24664 56876 24676
rect 56284 24636 56876 24664
rect 56284 24624 56290 24636
rect 56870 24624 56876 24636
rect 56928 24624 56934 24676
rect 56686 24596 56692 24608
rect 56152 24568 56692 24596
rect 56686 24556 56692 24568
rect 56744 24556 56750 24608
rect 58250 24596 58256 24608
rect 58211 24568 58256 24596
rect 58250 24556 58256 24568
rect 58308 24556 58314 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 20162 24392 20168 24404
rect 19536 24364 20168 24392
rect 17589 24259 17647 24265
rect 17589 24225 17601 24259
rect 17635 24256 17647 24259
rect 19426 24256 19432 24268
rect 17635 24228 19432 24256
rect 17635 24225 17647 24228
rect 17589 24219 17647 24225
rect 19426 24216 19432 24228
rect 19484 24216 19490 24268
rect 19536 24265 19564 24364
rect 20162 24352 20168 24364
rect 20220 24392 20226 24404
rect 24946 24392 24952 24404
rect 20220 24364 24952 24392
rect 20220 24352 20226 24364
rect 22554 24324 22560 24336
rect 20548 24296 22560 24324
rect 19521 24259 19579 24265
rect 19521 24225 19533 24259
rect 19567 24225 19579 24259
rect 19521 24219 19579 24225
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24188 1639 24191
rect 13078 24188 13084 24200
rect 1627 24160 13084 24188
rect 1627 24157 1639 24160
rect 1581 24151 1639 24157
rect 13078 24148 13084 24160
rect 13136 24148 13142 24200
rect 17494 24188 17500 24200
rect 17455 24160 17500 24188
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 17678 24148 17684 24200
rect 17736 24188 17742 24200
rect 17865 24191 17923 24197
rect 17865 24188 17877 24191
rect 17736 24160 17877 24188
rect 17736 24148 17742 24160
rect 17865 24157 17877 24160
rect 17911 24157 17923 24191
rect 17865 24151 17923 24157
rect 18049 24191 18107 24197
rect 18049 24157 18061 24191
rect 18095 24188 18107 24191
rect 19242 24188 19248 24200
rect 18095 24160 19248 24188
rect 18095 24157 18107 24160
rect 18049 24151 18107 24157
rect 19242 24148 19248 24160
rect 19300 24148 19306 24200
rect 19788 24191 19846 24197
rect 19788 24157 19800 24191
rect 19834 24188 19846 24191
rect 20070 24188 20076 24200
rect 19834 24160 20076 24188
rect 19834 24157 19846 24160
rect 19788 24151 19846 24157
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 1854 24120 1860 24132
rect 1815 24092 1860 24120
rect 1854 24080 1860 24092
rect 1912 24080 1918 24132
rect 16850 24120 16856 24132
rect 16811 24092 16856 24120
rect 16850 24080 16856 24092
rect 16908 24080 16914 24132
rect 17770 24080 17776 24132
rect 17828 24120 17834 24132
rect 20548 24120 20576 24296
rect 22554 24284 22560 24296
rect 22612 24284 22618 24336
rect 22646 24284 22652 24336
rect 22704 24324 22710 24336
rect 23017 24327 23075 24333
rect 23017 24324 23029 24327
rect 22704 24296 23029 24324
rect 22704 24284 22710 24296
rect 23017 24293 23029 24296
rect 23063 24324 23075 24327
rect 23063 24296 24440 24324
rect 23063 24293 23075 24296
rect 23017 24287 23075 24293
rect 21450 24216 21456 24268
rect 21508 24256 21514 24268
rect 21508 24228 21956 24256
rect 21508 24216 21514 24228
rect 21174 24148 21180 24200
rect 21232 24188 21238 24200
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 21232 24160 21373 24188
rect 21232 24148 21238 24160
rect 21361 24157 21373 24160
rect 21407 24157 21419 24191
rect 21542 24188 21548 24200
rect 21503 24160 21548 24188
rect 21361 24151 21419 24157
rect 21542 24148 21548 24160
rect 21600 24148 21606 24200
rect 21928 24120 21956 24228
rect 23014 24148 23020 24200
rect 23072 24188 23078 24200
rect 23569 24191 23627 24197
rect 23569 24188 23581 24191
rect 23072 24160 23581 24188
rect 23072 24148 23078 24160
rect 23569 24157 23581 24160
rect 23615 24157 23627 24191
rect 23569 24151 23627 24157
rect 23385 24123 23443 24129
rect 23385 24120 23397 24123
rect 17828 24092 20576 24120
rect 20640 24092 21772 24120
rect 21928 24092 23397 24120
rect 17828 24080 17834 24092
rect 19702 24012 19708 24064
rect 19760 24052 19766 24064
rect 20640 24052 20668 24092
rect 19760 24024 20668 24052
rect 20901 24055 20959 24061
rect 19760 24012 19766 24024
rect 20901 24021 20913 24055
rect 20947 24052 20959 24055
rect 21082 24052 21088 24064
rect 20947 24024 21088 24052
rect 20947 24021 20959 24024
rect 20901 24015 20959 24021
rect 21082 24012 21088 24024
rect 21140 24012 21146 24064
rect 21744 24061 21772 24092
rect 23385 24089 23397 24092
rect 23431 24120 23443 24123
rect 24412 24120 24440 24296
rect 24596 24265 24624 24364
rect 24946 24352 24952 24364
rect 25004 24352 25010 24404
rect 26418 24352 26424 24404
rect 26476 24392 26482 24404
rect 28994 24392 29000 24404
rect 26476 24364 29000 24392
rect 26476 24352 26482 24364
rect 28994 24352 29000 24364
rect 29052 24352 29058 24404
rect 30006 24352 30012 24404
rect 30064 24392 30070 24404
rect 30742 24392 30748 24404
rect 30064 24364 30748 24392
rect 30064 24352 30070 24364
rect 30742 24352 30748 24364
rect 30800 24352 30806 24404
rect 30926 24352 30932 24404
rect 30984 24392 30990 24404
rect 40034 24392 40040 24404
rect 30984 24364 40040 24392
rect 30984 24352 30990 24364
rect 40034 24352 40040 24364
rect 40092 24352 40098 24404
rect 58250 24392 58256 24404
rect 41386 24364 58256 24392
rect 27154 24284 27160 24336
rect 27212 24324 27218 24336
rect 29730 24324 29736 24336
rect 27212 24296 29736 24324
rect 27212 24284 27218 24296
rect 29730 24284 29736 24296
rect 29788 24324 29794 24336
rect 29914 24324 29920 24336
rect 29788 24296 29920 24324
rect 29788 24284 29794 24296
rect 29914 24284 29920 24296
rect 29972 24284 29978 24336
rect 35618 24284 35624 24336
rect 35676 24324 35682 24336
rect 41386 24324 41414 24364
rect 58250 24352 58256 24364
rect 58308 24352 58314 24404
rect 44634 24324 44640 24336
rect 35676 24296 41414 24324
rect 44595 24296 44640 24324
rect 35676 24284 35682 24296
rect 44634 24284 44640 24296
rect 44692 24284 44698 24336
rect 53929 24327 53987 24333
rect 53929 24293 53941 24327
rect 53975 24324 53987 24327
rect 55858 24324 55864 24336
rect 53975 24296 55864 24324
rect 53975 24293 53987 24296
rect 53929 24287 53987 24293
rect 24581 24259 24639 24265
rect 24581 24225 24593 24259
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 27062 24216 27068 24268
rect 27120 24256 27126 24268
rect 29638 24256 29644 24268
rect 27120 24228 29644 24256
rect 27120 24216 27126 24228
rect 29638 24216 29644 24228
rect 29696 24216 29702 24268
rect 44818 24216 44824 24268
rect 44876 24256 44882 24268
rect 45002 24256 45008 24268
rect 44876 24228 45008 24256
rect 44876 24216 44882 24228
rect 45002 24216 45008 24228
rect 45060 24256 45066 24268
rect 45060 24228 51074 24256
rect 45060 24216 45066 24228
rect 24848 24191 24906 24197
rect 24848 24157 24860 24191
rect 24894 24188 24906 24191
rect 25590 24188 25596 24200
rect 24894 24160 25596 24188
rect 24894 24157 24906 24160
rect 24848 24151 24906 24157
rect 25590 24148 25596 24160
rect 25648 24148 25654 24200
rect 26421 24191 26479 24197
rect 26421 24157 26433 24191
rect 26467 24188 26479 24191
rect 27522 24188 27528 24200
rect 26467 24160 27528 24188
rect 26467 24157 26479 24160
rect 26421 24151 26479 24157
rect 27522 24148 27528 24160
rect 27580 24148 27586 24200
rect 30009 24191 30067 24197
rect 30009 24157 30021 24191
rect 30055 24188 30067 24191
rect 31941 24191 31999 24197
rect 31941 24188 31953 24191
rect 30055 24160 31953 24188
rect 30055 24157 30067 24160
rect 30009 24151 30067 24157
rect 31941 24157 31953 24160
rect 31987 24188 31999 24191
rect 34790 24188 34796 24200
rect 31987 24160 34796 24188
rect 31987 24157 31999 24160
rect 31941 24151 31999 24157
rect 34790 24148 34796 24160
rect 34848 24148 34854 24200
rect 43257 24191 43315 24197
rect 43257 24157 43269 24191
rect 43303 24188 43315 24191
rect 44542 24188 44548 24200
rect 43303 24160 44548 24188
rect 43303 24157 43315 24160
rect 43257 24151 43315 24157
rect 44542 24148 44548 24160
rect 44600 24148 44606 24200
rect 50062 24148 50068 24200
rect 50120 24188 50126 24200
rect 50341 24191 50399 24197
rect 50341 24188 50353 24191
rect 50120 24160 50353 24188
rect 50120 24148 50126 24160
rect 50341 24157 50353 24160
rect 50387 24157 50399 24191
rect 50341 24151 50399 24157
rect 50525 24191 50583 24197
rect 50525 24157 50537 24191
rect 50571 24188 50583 24191
rect 50890 24188 50896 24200
rect 50571 24160 50896 24188
rect 50571 24157 50583 24160
rect 50525 24151 50583 24157
rect 50890 24148 50896 24160
rect 50948 24148 50954 24200
rect 51046 24188 51074 24228
rect 51534 24216 51540 24268
rect 51592 24256 51598 24268
rect 52089 24259 52147 24265
rect 51592 24228 51764 24256
rect 51592 24216 51598 24228
rect 51626 24188 51632 24200
rect 51046 24160 51488 24188
rect 51587 24160 51632 24188
rect 30276 24123 30334 24129
rect 23431 24092 23520 24120
rect 24412 24092 27660 24120
rect 23431 24089 23443 24092
rect 23385 24083 23443 24089
rect 21729 24055 21787 24061
rect 21729 24021 21741 24055
rect 21775 24052 21787 24055
rect 21818 24052 21824 24064
rect 21775 24024 21824 24052
rect 21775 24021 21787 24024
rect 21729 24015 21787 24021
rect 21818 24012 21824 24024
rect 21876 24012 21882 24064
rect 22278 24012 22284 24064
rect 22336 24052 22342 24064
rect 23014 24052 23020 24064
rect 22336 24024 23020 24052
rect 22336 24012 22342 24024
rect 23014 24012 23020 24024
rect 23072 24012 23078 24064
rect 23198 24052 23204 24064
rect 23159 24024 23204 24052
rect 23198 24012 23204 24024
rect 23256 24012 23262 24064
rect 23290 24012 23296 24064
rect 23348 24052 23354 24064
rect 23492 24052 23520 24092
rect 25130 24052 25136 24064
rect 23348 24024 23393 24052
rect 23492 24024 25136 24052
rect 23348 24012 23354 24024
rect 25130 24012 25136 24024
rect 25188 24012 25194 24064
rect 25222 24012 25228 24064
rect 25280 24052 25286 24064
rect 25958 24052 25964 24064
rect 25280 24024 25964 24052
rect 25280 24012 25286 24024
rect 25958 24012 25964 24024
rect 26016 24012 26022 24064
rect 27632 24061 27660 24092
rect 30276 24089 30288 24123
rect 30322 24120 30334 24123
rect 31110 24120 31116 24132
rect 30322 24092 31116 24120
rect 30322 24089 30334 24092
rect 30276 24083 30334 24089
rect 31110 24080 31116 24092
rect 31168 24080 31174 24132
rect 32208 24123 32266 24129
rect 32208 24089 32220 24123
rect 32254 24120 32266 24123
rect 32306 24120 32312 24132
rect 32254 24092 32312 24120
rect 32254 24089 32266 24092
rect 32208 24083 32266 24089
rect 32306 24080 32312 24092
rect 32364 24080 32370 24132
rect 43524 24123 43582 24129
rect 43524 24089 43536 24123
rect 43570 24120 43582 24123
rect 44450 24120 44456 24132
rect 43570 24092 44456 24120
rect 43570 24089 43582 24092
rect 43524 24083 43582 24089
rect 44450 24080 44456 24092
rect 44508 24080 44514 24132
rect 50798 24080 50804 24132
rect 50856 24120 50862 24132
rect 51350 24120 51356 24132
rect 50856 24092 51356 24120
rect 50856 24080 50862 24092
rect 51350 24080 51356 24092
rect 51408 24080 51414 24132
rect 51460 24120 51488 24160
rect 51626 24148 51632 24160
rect 51684 24148 51690 24200
rect 51736 24188 51764 24228
rect 52089 24225 52101 24259
rect 52135 24256 52147 24259
rect 52135 24228 52684 24256
rect 52135 24225 52147 24228
rect 52089 24219 52147 24225
rect 51931 24191 51989 24197
rect 51931 24188 51943 24191
rect 51736 24160 51943 24188
rect 51931 24157 51943 24160
rect 51977 24157 51989 24191
rect 52546 24188 52552 24200
rect 52507 24160 52552 24188
rect 51931 24151 51989 24157
rect 52546 24148 52552 24160
rect 52604 24148 52610 24200
rect 52656 24188 52684 24228
rect 53944 24188 53972 24287
rect 55858 24284 55864 24296
rect 55916 24284 55922 24336
rect 57422 24324 57428 24336
rect 57383 24296 57428 24324
rect 57422 24284 57428 24296
rect 57480 24284 57486 24336
rect 54478 24256 54484 24268
rect 54439 24228 54484 24256
rect 54478 24216 54484 24228
rect 54536 24216 54542 24268
rect 54662 24188 54668 24200
rect 52656 24160 53972 24188
rect 54623 24160 54668 24188
rect 54662 24148 54668 24160
rect 54720 24148 54726 24200
rect 56042 24188 56048 24200
rect 56003 24160 56048 24188
rect 56042 24148 56048 24160
rect 56100 24148 56106 24200
rect 56318 24197 56324 24200
rect 56312 24188 56324 24197
rect 56279 24160 56324 24188
rect 56312 24151 56324 24160
rect 56318 24148 56324 24151
rect 56376 24148 56382 24200
rect 57882 24188 57888 24200
rect 57843 24160 57888 24188
rect 57882 24148 57888 24160
rect 57940 24148 57946 24200
rect 59078 24188 59084 24200
rect 57992 24160 59084 24188
rect 51721 24123 51779 24129
rect 51721 24120 51733 24123
rect 51460 24092 51733 24120
rect 51721 24089 51733 24092
rect 51767 24089 51779 24123
rect 51721 24083 51779 24089
rect 51810 24080 51816 24132
rect 51868 24120 51874 24132
rect 52816 24123 52874 24129
rect 51868 24092 51913 24120
rect 51868 24080 51874 24092
rect 52816 24089 52828 24123
rect 52862 24120 52874 24123
rect 53282 24120 53288 24132
rect 52862 24092 53288 24120
rect 52862 24089 52874 24092
rect 52816 24083 52874 24089
rect 53282 24080 53288 24092
rect 53340 24080 53346 24132
rect 54018 24080 54024 24132
rect 54076 24120 54082 24132
rect 54076 24092 54984 24120
rect 54076 24080 54082 24092
rect 27617 24055 27675 24061
rect 27617 24021 27629 24055
rect 27663 24021 27675 24055
rect 27617 24015 27675 24021
rect 27982 24012 27988 24064
rect 28040 24052 28046 24064
rect 31389 24055 31447 24061
rect 31389 24052 31401 24055
rect 28040 24024 31401 24052
rect 28040 24012 28046 24024
rect 31389 24021 31401 24024
rect 31435 24021 31447 24055
rect 31389 24015 31447 24021
rect 32674 24012 32680 24064
rect 32732 24052 32738 24064
rect 33321 24055 33379 24061
rect 33321 24052 33333 24055
rect 32732 24024 33333 24052
rect 32732 24012 32738 24024
rect 33321 24021 33333 24024
rect 33367 24021 33379 24055
rect 33321 24015 33379 24021
rect 43346 24012 43352 24064
rect 43404 24052 43410 24064
rect 44634 24052 44640 24064
rect 43404 24024 44640 24052
rect 43404 24012 43410 24024
rect 44634 24012 44640 24024
rect 44692 24012 44698 24064
rect 50614 24012 50620 24064
rect 50672 24052 50678 24064
rect 50709 24055 50767 24061
rect 50709 24052 50721 24055
rect 50672 24024 50721 24052
rect 50672 24012 50678 24024
rect 50709 24021 50721 24024
rect 50755 24021 50767 24055
rect 50709 24015 50767 24021
rect 51445 24055 51503 24061
rect 51445 24021 51457 24055
rect 51491 24052 51503 24055
rect 53098 24052 53104 24064
rect 51491 24024 53104 24052
rect 51491 24021 51503 24024
rect 51445 24015 51503 24021
rect 53098 24012 53104 24024
rect 53156 24012 53162 24064
rect 54846 24052 54852 24064
rect 54807 24024 54852 24052
rect 54846 24012 54852 24024
rect 54904 24012 54910 24064
rect 54956 24052 54984 24092
rect 55030 24080 55036 24132
rect 55088 24120 55094 24132
rect 57992 24120 58020 24160
rect 59078 24148 59084 24160
rect 59136 24148 59142 24200
rect 58158 24120 58164 24132
rect 55088 24092 58020 24120
rect 58119 24092 58164 24120
rect 55088 24080 55094 24092
rect 58158 24080 58164 24092
rect 58216 24080 58222 24132
rect 57974 24052 57980 24064
rect 54956 24024 57980 24052
rect 57974 24012 57980 24024
rect 58032 24012 58038 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 19978 23808 19984 23860
rect 20036 23848 20042 23860
rect 20165 23851 20223 23857
rect 20165 23848 20177 23851
rect 20036 23820 20177 23848
rect 20036 23808 20042 23820
rect 20165 23817 20177 23820
rect 20211 23817 20223 23851
rect 20622 23848 20628 23860
rect 20583 23820 20628 23848
rect 20165 23811 20223 23817
rect 20622 23808 20628 23820
rect 20680 23808 20686 23860
rect 22278 23848 22284 23860
rect 22239 23820 22284 23848
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 27062 23848 27068 23860
rect 22388 23820 27068 23848
rect 15194 23780 15200 23792
rect 13556 23752 15200 23780
rect 13556 23721 13584 23752
rect 15194 23740 15200 23752
rect 15252 23740 15258 23792
rect 17586 23780 17592 23792
rect 15396 23752 17592 23780
rect 1581 23715 1639 23721
rect 1581 23681 1593 23715
rect 1627 23712 1639 23715
rect 13541 23715 13599 23721
rect 1627 23684 9674 23712
rect 1627 23681 1639 23684
rect 1581 23675 1639 23681
rect 1762 23644 1768 23656
rect 1723 23616 1768 23644
rect 1762 23604 1768 23616
rect 1820 23604 1826 23656
rect 9646 23508 9674 23684
rect 13541 23681 13553 23715
rect 13587 23681 13599 23715
rect 13541 23675 13599 23681
rect 13695 23715 13753 23721
rect 13695 23681 13707 23715
rect 13741 23712 13753 23715
rect 15396 23712 15424 23752
rect 17586 23740 17592 23752
rect 17644 23740 17650 23792
rect 19058 23740 19064 23792
rect 19116 23780 19122 23792
rect 19153 23783 19211 23789
rect 19153 23780 19165 23783
rect 19116 23752 19165 23780
rect 19116 23740 19122 23752
rect 19153 23749 19165 23752
rect 19199 23780 19211 23783
rect 19242 23780 19248 23792
rect 19199 23752 19248 23780
rect 19199 23749 19211 23752
rect 19153 23743 19211 23749
rect 19242 23740 19248 23752
rect 19300 23740 19306 23792
rect 20533 23783 20591 23789
rect 20533 23749 20545 23783
rect 20579 23780 20591 23783
rect 22388 23780 22416 23820
rect 27062 23808 27068 23820
rect 27120 23808 27126 23860
rect 27246 23848 27252 23860
rect 27207 23820 27252 23848
rect 27246 23808 27252 23820
rect 27304 23808 27310 23860
rect 27522 23808 27528 23860
rect 27580 23848 27586 23860
rect 29549 23851 29607 23857
rect 29549 23848 29561 23851
rect 27580 23820 29561 23848
rect 27580 23808 27586 23820
rect 29549 23817 29561 23820
rect 29595 23817 29607 23851
rect 29549 23811 29607 23817
rect 29914 23808 29920 23860
rect 29972 23848 29978 23860
rect 31110 23848 31116 23860
rect 29972 23820 30328 23848
rect 31071 23820 31116 23848
rect 29972 23808 29978 23820
rect 20579 23752 22416 23780
rect 22480 23752 23980 23780
rect 20579 23749 20591 23752
rect 20533 23743 20591 23749
rect 15562 23712 15568 23724
rect 13741 23684 15424 23712
rect 15523 23684 15568 23712
rect 13741 23681 13753 23684
rect 13695 23675 13753 23681
rect 15562 23672 15568 23684
rect 15620 23672 15626 23724
rect 15719 23715 15777 23721
rect 15719 23681 15731 23715
rect 15765 23712 15777 23715
rect 17770 23712 17776 23724
rect 15765 23684 17776 23712
rect 15765 23681 15777 23684
rect 15719 23675 15777 23681
rect 17770 23672 17776 23684
rect 17828 23672 17834 23724
rect 18138 23712 18144 23724
rect 18099 23684 18144 23712
rect 18138 23672 18144 23684
rect 18196 23672 18202 23724
rect 21818 23672 21824 23724
rect 21876 23712 21882 23724
rect 22222 23715 22280 23721
rect 22222 23712 22234 23715
rect 21876 23684 22234 23712
rect 21876 23672 21882 23684
rect 22222 23681 22234 23684
rect 22268 23681 22280 23715
rect 22222 23675 22280 23681
rect 13906 23644 13912 23656
rect 13867 23616 13912 23644
rect 13906 23604 13912 23616
rect 13964 23604 13970 23656
rect 20438 23604 20444 23656
rect 20496 23644 20502 23656
rect 20717 23647 20775 23653
rect 20717 23644 20729 23647
rect 20496 23616 20729 23644
rect 20496 23604 20502 23616
rect 20717 23613 20729 23616
rect 20763 23613 20775 23647
rect 20717 23607 20775 23613
rect 22094 23604 22100 23656
rect 22152 23644 22158 23656
rect 22480 23644 22508 23752
rect 22738 23712 22744 23724
rect 22699 23684 22744 23712
rect 22738 23672 22744 23684
rect 22796 23672 22802 23724
rect 23198 23672 23204 23724
rect 23256 23712 23262 23724
rect 23952 23721 23980 23752
rect 24210 23740 24216 23792
rect 24268 23780 24274 23792
rect 27154 23780 27160 23792
rect 24268 23752 27160 23780
rect 24268 23740 24274 23752
rect 27154 23740 27160 23752
rect 27212 23740 27218 23792
rect 30098 23780 30104 23792
rect 27724 23752 30104 23780
rect 27724 23721 27752 23752
rect 30098 23740 30104 23752
rect 30156 23740 30162 23792
rect 30300 23780 30328 23820
rect 31110 23808 31116 23820
rect 31168 23808 31174 23860
rect 32861 23851 32919 23857
rect 32861 23848 32873 23851
rect 31220 23820 32873 23848
rect 31220 23780 31248 23820
rect 32861 23817 32873 23820
rect 32907 23817 32919 23851
rect 36170 23848 36176 23860
rect 32861 23811 32919 23817
rect 33520 23820 36176 23848
rect 32674 23780 32680 23792
rect 30300 23752 31248 23780
rect 32635 23752 32680 23780
rect 32674 23740 32680 23752
rect 32732 23740 32738 23792
rect 23293 23715 23351 23721
rect 23293 23712 23305 23715
rect 23256 23684 23305 23712
rect 23256 23672 23262 23684
rect 23293 23681 23305 23684
rect 23339 23681 23351 23715
rect 23293 23675 23351 23681
rect 23937 23715 23995 23721
rect 23937 23681 23949 23715
rect 23983 23712 23995 23715
rect 27525 23715 27583 23721
rect 23983 23684 27476 23712
rect 23983 23681 23995 23684
rect 23937 23675 23995 23681
rect 22646 23644 22652 23656
rect 22152 23616 22508 23644
rect 22607 23616 22652 23644
rect 22152 23604 22158 23616
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 23308 23644 23336 23675
rect 25038 23644 25044 23656
rect 23308 23616 25044 23644
rect 25038 23604 25044 23616
rect 25096 23604 25102 23656
rect 15933 23579 15991 23585
rect 15933 23576 15945 23579
rect 12406 23548 15945 23576
rect 12406 23508 12434 23548
rect 15933 23545 15945 23548
rect 15979 23545 15991 23579
rect 15933 23539 15991 23545
rect 20530 23536 20536 23588
rect 20588 23576 20594 23588
rect 25133 23579 25191 23585
rect 25133 23576 25145 23579
rect 20588 23548 25145 23576
rect 20588 23536 20594 23548
rect 25133 23545 25145 23548
rect 25179 23545 25191 23579
rect 25133 23539 25191 23545
rect 9646 23480 12434 23508
rect 19794 23468 19800 23520
rect 19852 23508 19858 23520
rect 21450 23508 21456 23520
rect 19852 23480 21456 23508
rect 19852 23468 19858 23480
rect 21450 23468 21456 23480
rect 21508 23468 21514 23520
rect 21726 23468 21732 23520
rect 21784 23508 21790 23520
rect 22097 23511 22155 23517
rect 22097 23508 22109 23511
rect 21784 23480 22109 23508
rect 21784 23468 21790 23480
rect 22097 23477 22109 23480
rect 22143 23477 22155 23511
rect 22097 23471 22155 23477
rect 23385 23511 23443 23517
rect 23385 23477 23397 23511
rect 23431 23508 23443 23511
rect 24302 23508 24308 23520
rect 23431 23480 24308 23508
rect 23431 23477 23443 23480
rect 23385 23471 23443 23477
rect 24302 23468 24308 23480
rect 24360 23468 24366 23520
rect 27448 23508 27476 23684
rect 27525 23681 27537 23715
rect 27571 23681 27583 23715
rect 27525 23675 27583 23681
rect 27617 23715 27675 23721
rect 27617 23681 27629 23715
rect 27663 23681 27675 23715
rect 27617 23675 27675 23681
rect 27709 23715 27767 23721
rect 27709 23681 27721 23715
rect 27755 23681 27767 23715
rect 27890 23712 27896 23724
rect 27851 23684 27896 23712
rect 27709 23675 27767 23681
rect 27540 23576 27568 23675
rect 27632 23644 27660 23675
rect 27890 23672 27896 23684
rect 27948 23672 27954 23724
rect 27982 23672 27988 23724
rect 28040 23712 28046 23724
rect 28353 23715 28411 23721
rect 28353 23712 28365 23715
rect 28040 23684 28365 23712
rect 28040 23672 28046 23684
rect 28353 23681 28365 23684
rect 28399 23681 28411 23715
rect 28353 23675 28411 23681
rect 28994 23672 29000 23724
rect 29052 23712 29058 23724
rect 29052 23684 30144 23712
rect 29052 23672 29058 23684
rect 30116 23656 30144 23684
rect 31294 23672 31300 23724
rect 31352 23710 31358 23724
rect 31389 23715 31447 23721
rect 31389 23710 31401 23715
rect 31352 23682 31401 23710
rect 31352 23672 31358 23682
rect 31389 23681 31401 23682
rect 31435 23681 31447 23715
rect 31389 23675 31447 23681
rect 31478 23715 31536 23721
rect 31478 23681 31490 23715
rect 31524 23681 31536 23715
rect 31478 23675 31536 23681
rect 29730 23644 29736 23656
rect 27632 23616 29736 23644
rect 29730 23604 29736 23616
rect 29788 23604 29794 23656
rect 30098 23604 30104 23656
rect 30156 23644 30162 23656
rect 31493 23644 31521 23675
rect 31570 23672 31576 23724
rect 31628 23712 31634 23724
rect 31628 23684 31673 23712
rect 31628 23672 31634 23684
rect 31754 23672 31760 23724
rect 31812 23712 31818 23724
rect 32858 23712 32864 23724
rect 31812 23684 32864 23712
rect 31812 23672 31818 23684
rect 32858 23672 32864 23684
rect 32916 23672 32922 23724
rect 31846 23644 31852 23656
rect 30156 23616 31852 23644
rect 30156 23604 30162 23616
rect 31846 23604 31852 23616
rect 31904 23604 31910 23656
rect 32122 23604 32128 23656
rect 32180 23644 32186 23656
rect 32953 23647 33011 23653
rect 32953 23644 32965 23647
rect 32180 23616 32965 23644
rect 32180 23604 32186 23616
rect 32953 23613 32965 23616
rect 32999 23644 33011 23647
rect 33520 23644 33548 23820
rect 36170 23808 36176 23820
rect 36228 23808 36234 23860
rect 40402 23848 40408 23860
rect 40363 23820 40408 23848
rect 40402 23808 40408 23820
rect 40460 23808 40466 23860
rect 56502 23848 56508 23860
rect 41386 23820 56508 23848
rect 41386 23780 41414 23820
rect 56502 23808 56508 23820
rect 56560 23808 56566 23860
rect 57514 23848 57520 23860
rect 57475 23820 57520 23848
rect 57514 23808 57520 23820
rect 57572 23808 57578 23860
rect 32999 23616 33548 23644
rect 33612 23752 41414 23780
rect 41969 23783 42027 23789
rect 32999 23613 33011 23616
rect 32953 23607 33011 23613
rect 28258 23576 28264 23588
rect 27540 23548 28264 23576
rect 28258 23536 28264 23548
rect 28316 23576 28322 23588
rect 30926 23576 30932 23588
rect 28316 23548 30932 23576
rect 28316 23536 28322 23548
rect 30926 23536 30932 23548
rect 30984 23536 30990 23588
rect 32674 23576 32680 23588
rect 32324 23548 32680 23576
rect 29086 23508 29092 23520
rect 27448 23480 29092 23508
rect 29086 23468 29092 23480
rect 29144 23468 29150 23520
rect 31662 23468 31668 23520
rect 31720 23508 31726 23520
rect 32324 23508 32352 23548
rect 32674 23536 32680 23548
rect 32732 23536 32738 23588
rect 31720 23480 32352 23508
rect 32401 23511 32459 23517
rect 31720 23468 31726 23480
rect 32401 23477 32413 23511
rect 32447 23508 32459 23511
rect 33612 23508 33640 23752
rect 41969 23749 41981 23783
rect 42015 23780 42027 23783
rect 42858 23783 42916 23789
rect 42858 23780 42870 23783
rect 42015 23752 42870 23780
rect 42015 23749 42027 23752
rect 41969 23743 42027 23749
rect 42858 23749 42870 23752
rect 42904 23749 42916 23783
rect 52546 23780 52552 23792
rect 42858 23743 42916 23749
rect 43732 23752 44680 23780
rect 33956 23715 34014 23721
rect 33956 23681 33968 23715
rect 34002 23712 34014 23715
rect 34698 23712 34704 23724
rect 34002 23684 34704 23712
rect 34002 23681 34014 23684
rect 33956 23675 34014 23681
rect 34698 23672 34704 23684
rect 34756 23672 34762 23724
rect 36446 23712 36452 23724
rect 36407 23684 36452 23712
rect 36446 23672 36452 23684
rect 36504 23672 36510 23724
rect 36633 23715 36691 23721
rect 36633 23681 36645 23715
rect 36679 23681 36691 23715
rect 38378 23712 38384 23724
rect 38339 23684 38384 23712
rect 36633 23675 36691 23681
rect 33689 23647 33747 23653
rect 33689 23613 33701 23647
rect 33735 23613 33747 23647
rect 33689 23607 33747 23613
rect 32447 23480 33640 23508
rect 33704 23508 33732 23607
rect 35894 23604 35900 23656
rect 35952 23644 35958 23656
rect 36648 23644 36676 23675
rect 38378 23672 38384 23684
rect 38436 23672 38442 23724
rect 39114 23672 39120 23724
rect 39172 23712 39178 23724
rect 39281 23715 39339 23721
rect 39281 23712 39293 23715
rect 39172 23684 39293 23712
rect 39172 23672 39178 23684
rect 39281 23681 39293 23684
rect 39327 23681 39339 23715
rect 41874 23712 41880 23724
rect 41835 23684 41880 23712
rect 39281 23675 39339 23681
rect 41874 23672 41880 23684
rect 41932 23672 41938 23724
rect 42061 23715 42119 23721
rect 42061 23681 42073 23715
rect 42107 23712 42119 23715
rect 43732 23712 43760 23752
rect 44652 23724 44680 23752
rect 50356 23752 52552 23780
rect 42107 23684 43760 23712
rect 42107 23681 42119 23684
rect 42061 23675 42119 23681
rect 44358 23672 44364 23724
rect 44416 23712 44422 23724
rect 44453 23715 44511 23721
rect 44453 23712 44465 23715
rect 44416 23684 44465 23712
rect 44416 23672 44422 23684
rect 44453 23681 44465 23684
rect 44499 23681 44511 23715
rect 44634 23712 44640 23724
rect 44595 23684 44640 23712
rect 44453 23675 44511 23681
rect 44634 23672 44640 23684
rect 44692 23672 44698 23724
rect 50356 23721 50384 23752
rect 52546 23740 52552 23752
rect 52604 23780 52610 23792
rect 56042 23780 56048 23792
rect 52604 23752 56048 23780
rect 52604 23740 52610 23752
rect 50614 23721 50620 23724
rect 50341 23715 50399 23721
rect 50341 23681 50353 23715
rect 50387 23681 50399 23715
rect 50608 23712 50620 23721
rect 50575 23684 50620 23712
rect 50341 23675 50399 23681
rect 50608 23675 50620 23684
rect 37826 23644 37832 23656
rect 35952 23616 37832 23644
rect 35952 23604 35958 23616
rect 37826 23604 37832 23616
rect 37884 23604 37890 23656
rect 38197 23647 38255 23653
rect 38197 23613 38209 23647
rect 38243 23644 38255 23647
rect 38746 23644 38752 23656
rect 38243 23616 38752 23644
rect 38243 23613 38255 23616
rect 38197 23607 38255 23613
rect 38746 23604 38752 23616
rect 38804 23604 38810 23656
rect 38930 23604 38936 23656
rect 38988 23644 38994 23656
rect 39025 23647 39083 23653
rect 39025 23644 39037 23647
rect 38988 23616 39037 23644
rect 38988 23604 38994 23616
rect 39025 23613 39037 23616
rect 39071 23613 39083 23647
rect 39025 23607 39083 23613
rect 40402 23604 40408 23656
rect 40460 23644 40466 23656
rect 42613 23647 42671 23653
rect 42613 23644 42625 23647
rect 40460 23616 42625 23644
rect 40460 23604 40466 23616
rect 42613 23613 42625 23616
rect 42659 23613 42671 23647
rect 42613 23607 42671 23613
rect 44542 23604 44548 23656
rect 44600 23644 44606 23656
rect 50356 23644 50384 23675
rect 50614 23672 50620 23675
rect 50672 23672 50678 23724
rect 53098 23712 53104 23724
rect 53059 23684 53104 23712
rect 53098 23672 53104 23684
rect 53156 23672 53162 23724
rect 53282 23712 53288 23724
rect 53243 23684 53288 23712
rect 53282 23672 53288 23684
rect 53340 23672 53346 23724
rect 53760 23721 53788 23752
rect 56042 23740 56048 23752
rect 56100 23780 56106 23792
rect 56870 23780 56876 23792
rect 56100 23752 56876 23780
rect 56100 23740 56106 23752
rect 53745 23715 53803 23721
rect 53745 23681 53757 23715
rect 53791 23681 53803 23715
rect 53745 23675 53803 23681
rect 54012 23715 54070 23721
rect 54012 23681 54024 23715
rect 54058 23712 54070 23715
rect 54846 23712 54852 23724
rect 54058 23684 54852 23712
rect 54058 23681 54070 23684
rect 54012 23675 54070 23681
rect 54846 23672 54852 23684
rect 54904 23672 54910 23724
rect 56152 23721 56180 23752
rect 56870 23740 56876 23752
rect 56928 23740 56934 23792
rect 56410 23721 56416 23724
rect 56137 23715 56195 23721
rect 56137 23681 56149 23715
rect 56183 23681 56195 23715
rect 56137 23675 56195 23681
rect 56404 23675 56416 23721
rect 56468 23712 56474 23724
rect 56468 23684 56504 23712
rect 56410 23672 56416 23675
rect 56468 23672 56474 23684
rect 44600 23616 50384 23644
rect 44600 23604 44606 23616
rect 51994 23604 52000 23656
rect 52052 23644 52058 23656
rect 52917 23647 52975 23653
rect 52917 23644 52929 23647
rect 52052 23616 52929 23644
rect 52052 23604 52058 23616
rect 52917 23613 52929 23616
rect 52963 23613 52975 23647
rect 52917 23607 52975 23613
rect 35066 23576 35072 23588
rect 35027 23548 35072 23576
rect 35066 23536 35072 23548
rect 35124 23536 35130 23588
rect 35434 23536 35440 23588
rect 35492 23576 35498 23588
rect 35802 23576 35808 23588
rect 35492 23548 35808 23576
rect 35492 23536 35498 23548
rect 35802 23536 35808 23548
rect 35860 23536 35866 23588
rect 40034 23536 40040 23588
rect 40092 23576 40098 23588
rect 51718 23576 51724 23588
rect 40092 23548 41414 23576
rect 40092 23536 40098 23548
rect 34790 23508 34796 23520
rect 33704 23480 34796 23508
rect 32447 23477 32459 23480
rect 32401 23471 32459 23477
rect 34790 23468 34796 23480
rect 34848 23468 34854 23520
rect 36722 23468 36728 23520
rect 36780 23508 36786 23520
rect 36817 23511 36875 23517
rect 36817 23508 36829 23511
rect 36780 23480 36829 23508
rect 36780 23468 36786 23480
rect 36817 23477 36829 23480
rect 36863 23477 36875 23511
rect 36817 23471 36875 23477
rect 38565 23511 38623 23517
rect 38565 23477 38577 23511
rect 38611 23508 38623 23511
rect 39022 23508 39028 23520
rect 38611 23480 39028 23508
rect 38611 23477 38623 23480
rect 38565 23471 38623 23477
rect 39022 23468 39028 23480
rect 39080 23468 39086 23520
rect 41386 23508 41414 23548
rect 43548 23548 46244 23576
rect 51679 23548 51724 23576
rect 43548 23508 43576 23548
rect 43990 23508 43996 23520
rect 41386 23480 43576 23508
rect 43951 23480 43996 23508
rect 43990 23468 43996 23480
rect 44048 23468 44054 23520
rect 44450 23508 44456 23520
rect 44411 23480 44456 23508
rect 44450 23468 44456 23480
rect 44508 23468 44514 23520
rect 46216 23508 46244 23548
rect 51718 23536 51724 23548
rect 51776 23536 51782 23588
rect 54018 23508 54024 23520
rect 46216 23480 54024 23508
rect 54018 23468 54024 23480
rect 54076 23468 54082 23520
rect 54386 23468 54392 23520
rect 54444 23508 54450 23520
rect 55125 23511 55183 23517
rect 55125 23508 55137 23511
rect 54444 23480 55137 23508
rect 54444 23468 54450 23480
rect 55125 23477 55137 23480
rect 55171 23508 55183 23511
rect 57790 23508 57796 23520
rect 55171 23480 57796 23508
rect 55171 23477 55183 23480
rect 55125 23471 55183 23477
rect 57790 23468 57796 23480
rect 57848 23468 57854 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 19794 23304 19800 23316
rect 19755 23276 19800 23304
rect 19794 23264 19800 23276
rect 19852 23264 19858 23316
rect 19981 23307 20039 23313
rect 19981 23273 19993 23307
rect 20027 23304 20039 23307
rect 22462 23304 22468 23316
rect 20027 23276 22468 23304
rect 20027 23273 20039 23276
rect 19981 23267 20039 23273
rect 22462 23264 22468 23276
rect 22520 23304 22526 23316
rect 24762 23304 24768 23316
rect 22520 23276 24768 23304
rect 22520 23264 22526 23276
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 25593 23307 25651 23313
rect 25593 23273 25605 23307
rect 25639 23304 25651 23307
rect 26234 23304 26240 23316
rect 25639 23276 26240 23304
rect 25639 23273 25651 23276
rect 25593 23267 25651 23273
rect 26234 23264 26240 23276
rect 26292 23264 26298 23316
rect 28077 23307 28135 23313
rect 28077 23304 28089 23307
rect 26344 23276 28089 23304
rect 19334 23196 19340 23248
rect 19392 23236 19398 23248
rect 20441 23239 20499 23245
rect 20441 23236 20453 23239
rect 19392 23208 20453 23236
rect 19392 23196 19398 23208
rect 20441 23205 20453 23208
rect 20487 23236 20499 23239
rect 20530 23236 20536 23248
rect 20487 23208 20536 23236
rect 20487 23205 20499 23208
rect 20441 23199 20499 23205
rect 20530 23196 20536 23208
rect 20588 23196 20594 23248
rect 24949 23239 25007 23245
rect 24949 23236 24961 23239
rect 22066 23208 24961 23236
rect 17586 23128 17592 23180
rect 17644 23168 17650 23180
rect 18417 23171 18475 23177
rect 18417 23168 18429 23171
rect 17644 23140 18429 23168
rect 17644 23128 17650 23140
rect 18417 23137 18429 23140
rect 18463 23137 18475 23171
rect 18874 23168 18880 23180
rect 18835 23140 18880 23168
rect 18417 23131 18475 23137
rect 1581 23103 1639 23109
rect 1581 23069 1593 23103
rect 1627 23100 1639 23103
rect 13906 23100 13912 23112
rect 1627 23072 13912 23100
rect 1627 23069 1639 23072
rect 1581 23063 1639 23069
rect 13906 23060 13912 23072
rect 13964 23060 13970 23112
rect 15930 23100 15936 23112
rect 15891 23072 15936 23100
rect 15930 23060 15936 23072
rect 15988 23060 15994 23112
rect 1854 23032 1860 23044
rect 1815 23004 1860 23032
rect 1854 22992 1860 23004
rect 1912 22992 1918 23044
rect 16200 23035 16258 23041
rect 16200 23001 16212 23035
rect 16246 23032 16258 23035
rect 17770 23032 17776 23044
rect 16246 23004 17776 23032
rect 16246 23001 16258 23004
rect 16200 22995 16258 23001
rect 17770 22992 17776 23004
rect 17828 22992 17834 23044
rect 18432 23032 18460 23131
rect 18874 23128 18880 23140
rect 18932 23128 18938 23180
rect 21174 23168 21180 23180
rect 20640 23140 21180 23168
rect 18509 23103 18567 23109
rect 18509 23069 18521 23103
rect 18555 23100 18567 23103
rect 19794 23100 19800 23112
rect 18555 23072 19800 23100
rect 18555 23069 18567 23072
rect 18509 23063 18567 23069
rect 19794 23060 19800 23072
rect 19852 23060 19858 23112
rect 20640 23109 20668 23140
rect 21174 23128 21180 23140
rect 21232 23128 21238 23180
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23069 20683 23103
rect 20625 23063 20683 23069
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 20993 23103 21051 23109
rect 20993 23100 21005 23103
rect 20864 23072 21005 23100
rect 20864 23060 20870 23072
rect 20993 23069 21005 23072
rect 21039 23069 21051 23103
rect 20993 23063 21051 23069
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23100 21787 23103
rect 22066 23100 22094 23208
rect 24949 23205 24961 23208
rect 24995 23205 25007 23239
rect 24949 23199 25007 23205
rect 25038 23196 25044 23248
rect 25096 23236 25102 23248
rect 26344 23236 26372 23276
rect 28077 23273 28089 23276
rect 28123 23273 28135 23307
rect 28077 23267 28135 23273
rect 29733 23307 29791 23313
rect 29733 23273 29745 23307
rect 29779 23304 29791 23307
rect 29822 23304 29828 23316
rect 29779 23276 29828 23304
rect 29779 23273 29791 23276
rect 29733 23267 29791 23273
rect 29822 23264 29828 23276
rect 29880 23264 29886 23316
rect 35345 23307 35403 23313
rect 35345 23273 35357 23307
rect 35391 23304 35403 23307
rect 35391 23276 38332 23304
rect 35391 23273 35403 23276
rect 35345 23267 35403 23273
rect 27890 23236 27896 23248
rect 25096 23208 26372 23236
rect 26528 23208 27896 23236
rect 25096 23196 25102 23208
rect 24673 23171 24731 23177
rect 24673 23137 24685 23171
rect 24719 23168 24731 23171
rect 24762 23168 24768 23180
rect 24719 23140 24768 23168
rect 24719 23137 24731 23140
rect 24673 23131 24731 23137
rect 24762 23128 24768 23140
rect 24820 23128 24826 23180
rect 26142 23168 26148 23180
rect 25976 23140 26148 23168
rect 24578 23100 24584 23112
rect 21775 23072 22094 23100
rect 24539 23072 24584 23100
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 24578 23060 24584 23072
rect 24636 23060 24642 23112
rect 25314 23100 25320 23112
rect 25275 23072 25320 23100
rect 25314 23060 25320 23072
rect 25372 23100 25378 23112
rect 25682 23100 25688 23112
rect 25372 23072 25688 23100
rect 25372 23060 25378 23072
rect 25682 23060 25688 23072
rect 25740 23100 25746 23112
rect 25976 23109 26004 23140
rect 26142 23128 26148 23140
rect 26200 23128 26206 23180
rect 25823 23103 25881 23109
rect 25823 23100 25835 23103
rect 25740 23072 25835 23100
rect 25740 23060 25746 23072
rect 25823 23069 25835 23072
rect 25869 23069 25881 23103
rect 25823 23063 25881 23069
rect 25961 23103 26019 23109
rect 25961 23069 25973 23103
rect 26007 23069 26019 23103
rect 25961 23063 26019 23069
rect 26050 23060 26056 23112
rect 26108 23100 26114 23112
rect 26237 23103 26295 23109
rect 26108 23072 26153 23100
rect 26108 23060 26114 23072
rect 26237 23069 26249 23103
rect 26283 23100 26295 23103
rect 26528 23100 26556 23208
rect 27890 23196 27896 23208
rect 27948 23236 27954 23248
rect 29914 23236 29920 23248
rect 27948 23208 29920 23236
rect 27948 23196 27954 23208
rect 29914 23196 29920 23208
rect 29972 23196 29978 23248
rect 30098 23196 30104 23248
rect 30156 23196 30162 23248
rect 37826 23196 37832 23248
rect 37884 23236 37890 23248
rect 37921 23239 37979 23245
rect 37921 23236 37933 23239
rect 37884 23208 37933 23236
rect 37884 23196 37890 23208
rect 37921 23205 37933 23208
rect 37967 23236 37979 23239
rect 38102 23236 38108 23248
rect 37967 23208 38108 23236
rect 37967 23205 37979 23208
rect 37921 23199 37979 23205
rect 38102 23196 38108 23208
rect 38160 23196 38166 23248
rect 38304 23236 38332 23276
rect 38378 23264 38384 23316
rect 38436 23304 38442 23316
rect 38473 23307 38531 23313
rect 38473 23304 38485 23307
rect 38436 23276 38485 23304
rect 38436 23264 38442 23276
rect 38473 23273 38485 23276
rect 38519 23273 38531 23307
rect 40586 23304 40592 23316
rect 38473 23267 38531 23273
rect 39040 23276 40592 23304
rect 39040 23236 39068 23276
rect 40586 23264 40592 23276
rect 40644 23264 40650 23316
rect 41874 23264 41880 23316
rect 41932 23304 41938 23316
rect 41969 23307 42027 23313
rect 41969 23304 41981 23307
rect 41932 23276 41981 23304
rect 41932 23264 41938 23276
rect 41969 23273 41981 23276
rect 42015 23273 42027 23307
rect 42518 23304 42524 23316
rect 42479 23276 42524 23304
rect 41969 23267 42027 23273
rect 42518 23264 42524 23276
rect 42576 23264 42582 23316
rect 43257 23307 43315 23313
rect 43257 23273 43269 23307
rect 43303 23304 43315 23307
rect 44358 23304 44364 23316
rect 43303 23276 44364 23304
rect 43303 23273 43315 23276
rect 43257 23267 43315 23273
rect 44358 23264 44364 23276
rect 44416 23264 44422 23316
rect 50890 23304 50896 23316
rect 50851 23276 50896 23304
rect 50890 23264 50896 23276
rect 50948 23264 50954 23316
rect 53745 23307 53803 23313
rect 53745 23273 53757 23307
rect 53791 23304 53803 23307
rect 54662 23304 54668 23316
rect 53791 23276 54668 23304
rect 53791 23273 53803 23276
rect 53745 23267 53803 23273
rect 54662 23264 54668 23276
rect 54720 23264 54726 23316
rect 58253 23307 58311 23313
rect 58253 23273 58265 23307
rect 58299 23304 58311 23307
rect 58342 23304 58348 23316
rect 58299 23276 58348 23304
rect 58299 23273 58311 23276
rect 58253 23267 58311 23273
rect 58342 23264 58348 23276
rect 58400 23264 58406 23316
rect 40310 23236 40316 23248
rect 38304 23208 39068 23236
rect 39132 23208 40316 23236
rect 26283 23072 26556 23100
rect 26697 23103 26755 23109
rect 26283 23069 26295 23072
rect 26237 23063 26295 23069
rect 26697 23069 26709 23103
rect 26743 23100 26755 23103
rect 28534 23100 28540 23112
rect 26743 23072 28540 23100
rect 26743 23069 26755 23072
rect 26697 23063 26755 23069
rect 19613 23035 19671 23041
rect 18432 23004 19564 23032
rect 17313 22967 17371 22973
rect 17313 22933 17325 22967
rect 17359 22964 17371 22967
rect 19426 22964 19432 22976
rect 17359 22936 19432 22964
rect 17359 22933 17371 22936
rect 17313 22927 17371 22933
rect 19426 22924 19432 22936
rect 19484 22924 19490 22976
rect 19536 22964 19564 23004
rect 19613 23001 19625 23035
rect 19659 23032 19671 23035
rect 20346 23032 20352 23044
rect 19659 23004 20352 23032
rect 19659 23001 19671 23004
rect 19613 22995 19671 23001
rect 20346 22992 20352 23004
rect 20404 22992 20410 23044
rect 20438 22992 20444 23044
rect 20496 23032 20502 23044
rect 20717 23035 20775 23041
rect 20496 23004 20668 23032
rect 20496 22992 20502 23004
rect 19813 22967 19871 22973
rect 19813 22964 19825 22967
rect 19536 22936 19825 22964
rect 19813 22933 19825 22936
rect 19859 22964 19871 22967
rect 20530 22964 20536 22976
rect 19859 22936 20536 22964
rect 19859 22933 19871 22936
rect 19813 22927 19871 22933
rect 20530 22924 20536 22936
rect 20588 22924 20594 22976
rect 20640 22964 20668 23004
rect 20717 23001 20729 23035
rect 20763 23032 20775 23035
rect 20898 23032 20904 23044
rect 20763 23004 20904 23032
rect 20763 23001 20775 23004
rect 20717 22995 20775 23001
rect 20898 22992 20904 23004
rect 20956 23032 20962 23044
rect 21542 23032 21548 23044
rect 20956 23004 21548 23032
rect 20956 22992 20962 23004
rect 21542 22992 21548 23004
rect 21600 22992 21606 23044
rect 23842 22992 23848 23044
rect 23900 23032 23906 23044
rect 26712 23032 26740 23063
rect 28534 23060 28540 23072
rect 28592 23060 28598 23112
rect 29638 23060 29644 23112
rect 29696 23100 29702 23112
rect 30113 23109 30141 23196
rect 31754 23168 31760 23180
rect 30852 23140 31760 23168
rect 30009 23103 30067 23109
rect 29696 23094 29868 23100
rect 30009 23094 30021 23103
rect 29696 23072 30021 23094
rect 29696 23060 29702 23072
rect 29840 23069 30021 23072
rect 30055 23069 30067 23103
rect 29840 23066 30067 23069
rect 30009 23063 30067 23066
rect 30098 23103 30156 23109
rect 30098 23069 30110 23103
rect 30144 23069 30156 23103
rect 30098 23063 30156 23069
rect 30190 23060 30196 23112
rect 30248 23109 30254 23112
rect 30248 23100 30256 23109
rect 30248 23072 30293 23100
rect 30248 23063 30256 23072
rect 30248 23060 30254 23063
rect 30374 23060 30380 23112
rect 30432 23100 30438 23112
rect 30852 23100 30880 23140
rect 31754 23128 31760 23140
rect 31812 23128 31818 23180
rect 36170 23168 36176 23180
rect 33520 23140 35480 23168
rect 31018 23100 31024 23112
rect 30432 23072 30880 23100
rect 30979 23072 31024 23100
rect 30432 23060 30438 23072
rect 31018 23060 31024 23072
rect 31076 23060 31082 23112
rect 33520 23032 33548 23140
rect 35452 23112 35480 23140
rect 35912 23140 36176 23168
rect 35434 23060 35440 23112
rect 35492 23100 35498 23112
rect 35912 23109 35940 23140
rect 36170 23128 36176 23140
rect 36228 23168 36234 23180
rect 39132 23177 39160 23208
rect 40310 23196 40316 23208
rect 40368 23236 40374 23248
rect 53834 23236 53840 23248
rect 40368 23208 53840 23236
rect 40368 23196 40374 23208
rect 53834 23196 53840 23208
rect 53892 23196 53898 23248
rect 39117 23171 39175 23177
rect 36228 23140 36676 23168
rect 36228 23128 36234 23140
rect 35897 23103 35955 23109
rect 35492 23072 35756 23100
rect 35492 23060 35498 23072
rect 23900 23004 26740 23032
rect 26804 23004 33548 23032
rect 33781 23035 33839 23041
rect 23900 22992 23906 23004
rect 20809 22967 20867 22973
rect 20809 22964 20821 22967
rect 20640 22936 20821 22964
rect 20809 22933 20821 22936
rect 20855 22964 20867 22967
rect 22278 22964 22284 22976
rect 20855 22936 22284 22964
rect 20855 22933 20867 22936
rect 20809 22927 20867 22933
rect 22278 22924 22284 22936
rect 22336 22924 22342 22976
rect 22922 22964 22928 22976
rect 22883 22936 22928 22964
rect 22922 22924 22928 22936
rect 22980 22924 22986 22976
rect 25590 22924 25596 22976
rect 25648 22964 25654 22976
rect 26804 22964 26832 23004
rect 33781 23001 33793 23035
rect 33827 23032 33839 23035
rect 33870 23032 33876 23044
rect 33827 23004 33876 23032
rect 33827 23001 33839 23004
rect 33781 22995 33839 23001
rect 33870 22992 33876 23004
rect 33928 22992 33934 23044
rect 33965 23035 34023 23041
rect 33965 23001 33977 23035
rect 34011 23032 34023 23035
rect 34330 23032 34336 23044
rect 34011 23004 34336 23032
rect 34011 23001 34023 23004
rect 33965 22995 34023 23001
rect 34330 22992 34336 23004
rect 34388 22992 34394 23044
rect 34606 22992 34612 23044
rect 34664 23032 34670 23044
rect 35621 23035 35679 23041
rect 34664 23004 35342 23032
rect 34664 22992 34670 23004
rect 25648 22936 26832 22964
rect 25648 22924 25654 22936
rect 26878 22924 26884 22976
rect 26936 22964 26942 22976
rect 32217 22967 32275 22973
rect 32217 22964 32229 22967
rect 26936 22936 32229 22964
rect 26936 22924 26942 22936
rect 32217 22933 32229 22936
rect 32263 22933 32275 22967
rect 34146 22964 34152 22976
rect 34107 22936 34152 22964
rect 32217 22927 32275 22933
rect 34146 22924 34152 22936
rect 34204 22924 34210 22976
rect 35314 22964 35342 23004
rect 35621 23001 35633 23035
rect 35667 23001 35679 23035
rect 35728 23032 35756 23072
rect 35897 23069 35909 23103
rect 35943 23069 35955 23103
rect 36538 23100 36544 23112
rect 36499 23072 36544 23100
rect 35897 23063 35955 23069
rect 36538 23060 36544 23072
rect 36596 23060 36602 23112
rect 36648 23100 36676 23140
rect 39117 23137 39129 23171
rect 39163 23137 39175 23171
rect 39117 23131 39175 23137
rect 39408 23140 40448 23168
rect 36648 23072 37044 23100
rect 37016 23044 37044 23072
rect 37826 23060 37832 23112
rect 37884 23100 37890 23112
rect 38657 23103 38715 23109
rect 38657 23100 38669 23103
rect 37884 23072 38669 23100
rect 37884 23060 37890 23072
rect 38657 23069 38669 23072
rect 38703 23069 38715 23103
rect 38657 23063 38715 23069
rect 38979 23103 39037 23109
rect 38979 23069 38991 23103
rect 39025 23100 39037 23103
rect 39408 23100 39436 23140
rect 39025 23072 39436 23100
rect 39025 23069 39037 23072
rect 38979 23063 39037 23069
rect 39482 23060 39488 23112
rect 39540 23100 39546 23112
rect 40313 23103 40371 23109
rect 39540 23094 40172 23100
rect 40221 23097 40279 23103
rect 40221 23094 40233 23097
rect 39540 23072 40233 23094
rect 39540 23060 39546 23072
rect 40144 23066 40233 23072
rect 40221 23063 40233 23066
rect 40267 23063 40279 23097
rect 40313 23069 40325 23103
rect 40359 23069 40371 23103
rect 40420 23100 40448 23140
rect 40494 23128 40500 23180
rect 40552 23168 40558 23180
rect 40681 23171 40739 23177
rect 40681 23168 40693 23171
rect 40552 23140 40693 23168
rect 40552 23128 40558 23140
rect 40681 23137 40693 23140
rect 40727 23137 40739 23171
rect 43990 23168 43996 23180
rect 40681 23131 40739 23137
rect 42536 23140 43996 23168
rect 42150 23103 42208 23109
rect 40420 23072 40540 23100
rect 40313 23063 40371 23069
rect 40221 23057 40279 23063
rect 35805 23035 35863 23041
rect 35805 23032 35817 23035
rect 35728 23004 35817 23032
rect 35621 22995 35679 23001
rect 35805 23001 35817 23004
rect 35851 23001 35863 23035
rect 35805 22995 35863 23001
rect 35636 22964 35664 22995
rect 36262 22992 36268 23044
rect 36320 23032 36326 23044
rect 36786 23035 36844 23041
rect 36786 23032 36798 23035
rect 36320 23004 36798 23032
rect 36320 22992 36326 23004
rect 36786 23001 36798 23004
rect 36832 23001 36844 23035
rect 36786 22995 36844 23001
rect 36998 22992 37004 23044
rect 37056 22992 37062 23044
rect 37274 22992 37280 23044
rect 37332 23032 37338 23044
rect 38749 23035 38807 23041
rect 38749 23032 38761 23035
rect 37332 23004 38761 23032
rect 37332 22992 37338 23004
rect 38749 23001 38761 23004
rect 38795 23001 38807 23035
rect 38749 22995 38807 23001
rect 38838 22992 38844 23044
rect 38896 23032 38902 23044
rect 40037 23035 40095 23041
rect 40037 23032 40049 23035
rect 38896 23004 38941 23032
rect 39960 23004 40049 23032
rect 38896 22992 38902 23004
rect 35314 22936 35664 22964
rect 36170 22924 36176 22976
rect 36228 22964 36234 22976
rect 39666 22964 39672 22976
rect 36228 22936 39672 22964
rect 36228 22924 36234 22936
rect 39666 22924 39672 22936
rect 39724 22924 39730 22976
rect 39758 22924 39764 22976
rect 39816 22964 39822 22976
rect 39960 22964 39988 23004
rect 40037 23001 40049 23004
rect 40083 23001 40095 23035
rect 40037 22995 40095 23001
rect 39816 22936 39988 22964
rect 39816 22924 39822 22936
rect 40218 22924 40224 22976
rect 40276 22964 40282 22976
rect 40328 22964 40356 23063
rect 40512 23044 40540 23072
rect 42150 23069 42162 23103
rect 42196 23100 42208 23103
rect 42536 23100 42564 23140
rect 43990 23128 43996 23140
rect 44048 23128 44054 23180
rect 54386 23168 54392 23180
rect 47964 23140 54248 23168
rect 54347 23140 54392 23168
rect 42196 23072 42564 23100
rect 42613 23103 42671 23109
rect 42196 23069 42208 23072
rect 42150 23063 42208 23069
rect 42613 23069 42625 23103
rect 42659 23100 42671 23103
rect 42794 23100 42800 23112
rect 42659 23072 42800 23100
rect 42659 23069 42671 23072
rect 42613 23063 42671 23069
rect 42794 23060 42800 23072
rect 42852 23060 42858 23112
rect 43346 23060 43352 23112
rect 43404 23109 43410 23112
rect 43404 23103 43440 23109
rect 43428 23069 43440 23103
rect 43404 23063 43440 23069
rect 43404 23060 43410 23063
rect 43714 23060 43720 23112
rect 43772 23100 43778 23112
rect 43809 23103 43867 23109
rect 43809 23100 43821 23103
rect 43772 23072 43821 23100
rect 43772 23060 43778 23072
rect 43809 23069 43821 23072
rect 43855 23069 43867 23103
rect 43809 23063 43867 23069
rect 43898 23060 43904 23112
rect 43956 23100 43962 23112
rect 44358 23100 44364 23112
rect 43956 23072 44364 23100
rect 43956 23060 43962 23072
rect 44358 23060 44364 23072
rect 44416 23060 44422 23112
rect 47964 23109 47992 23140
rect 47949 23103 48007 23109
rect 47949 23069 47961 23103
rect 47995 23069 48007 23103
rect 47949 23063 48007 23069
rect 48130 23060 48136 23112
rect 48188 23100 48194 23112
rect 50341 23103 50399 23109
rect 50341 23100 50353 23103
rect 48188 23072 50353 23100
rect 48188 23060 48194 23072
rect 50341 23069 50353 23072
rect 50387 23069 50399 23103
rect 50706 23100 50712 23112
rect 50667 23072 50712 23100
rect 50341 23063 50399 23069
rect 50706 23060 50712 23072
rect 50764 23060 50770 23112
rect 53926 23100 53932 23112
rect 53887 23072 53932 23100
rect 53926 23060 53932 23072
rect 53984 23060 53990 23112
rect 54110 23100 54116 23112
rect 54071 23072 54116 23100
rect 54110 23060 54116 23072
rect 54168 23060 54174 23112
rect 54220 23109 54248 23140
rect 54386 23128 54392 23140
rect 54444 23128 54450 23180
rect 56229 23171 56287 23177
rect 56229 23137 56241 23171
rect 56275 23168 56287 23171
rect 56502 23168 56508 23180
rect 56275 23140 56508 23168
rect 56275 23137 56287 23140
rect 56229 23131 56287 23137
rect 56502 23128 56508 23140
rect 56560 23128 56566 23180
rect 56870 23168 56876 23180
rect 56831 23140 56876 23168
rect 56870 23128 56876 23140
rect 56928 23128 56934 23180
rect 54220 23103 54289 23109
rect 54220 23072 54243 23103
rect 54231 23069 54243 23072
rect 54277 23100 54289 23103
rect 56042 23100 56048 23112
rect 54277 23072 56048 23100
rect 54277 23069 54289 23072
rect 54231 23063 54289 23069
rect 56042 23060 56048 23072
rect 56100 23060 56106 23112
rect 56137 23103 56195 23109
rect 56137 23069 56149 23103
rect 56183 23069 56195 23103
rect 56137 23063 56195 23069
rect 40405 23035 40463 23041
rect 40405 23001 40417 23035
rect 40451 23001 40463 23035
rect 40405 22995 40463 23001
rect 40276 22936 40356 22964
rect 40420 22964 40448 22995
rect 40494 22992 40500 23044
rect 40552 23041 40558 23044
rect 40552 23035 40581 23041
rect 40569 23032 40581 23035
rect 40569 23004 40645 23032
rect 40569 23001 40581 23004
rect 40552 22995 40581 23001
rect 40552 22992 40558 22995
rect 47854 22992 47860 23044
rect 47912 23032 47918 23044
rect 48225 23035 48283 23041
rect 48225 23032 48237 23035
rect 47912 23004 48237 23032
rect 47912 22992 47918 23004
rect 48225 23001 48237 23004
rect 48271 23001 48283 23035
rect 48225 22995 48283 23001
rect 40678 22964 40684 22976
rect 40420 22936 40684 22964
rect 40276 22924 40282 22936
rect 40678 22924 40684 22936
rect 40736 22924 40742 22976
rect 41414 22924 41420 22976
rect 41472 22964 41478 22976
rect 42153 22967 42211 22973
rect 42153 22964 42165 22967
rect 41472 22936 42165 22964
rect 41472 22924 41478 22936
rect 42153 22933 42165 22936
rect 42199 22964 42211 22967
rect 43441 22967 43499 22973
rect 43441 22964 43453 22967
rect 42199 22936 43453 22964
rect 42199 22933 42211 22936
rect 42153 22927 42211 22933
rect 43441 22933 43453 22936
rect 43487 22933 43499 22967
rect 48240 22964 48268 22995
rect 49970 22992 49976 23044
rect 50028 23032 50034 23044
rect 50525 23035 50583 23041
rect 50525 23032 50537 23035
rect 50028 23004 50537 23032
rect 50028 22992 50034 23004
rect 50525 23001 50537 23004
rect 50571 23001 50583 23035
rect 50525 22995 50583 23001
rect 50617 23035 50675 23041
rect 50617 23001 50629 23035
rect 50663 23032 50675 23035
rect 51718 23032 51724 23044
rect 50663 23004 51724 23032
rect 50663 23001 50675 23004
rect 50617 22995 50675 23001
rect 51718 22992 51724 23004
rect 51776 22992 51782 23044
rect 54021 23035 54079 23041
rect 54021 23032 54033 23035
rect 53392 23004 54033 23032
rect 53392 22976 53420 23004
rect 54021 23001 54033 23004
rect 54067 23001 54079 23035
rect 55950 23032 55956 23044
rect 55911 23004 55956 23032
rect 54021 22995 54079 23001
rect 55950 22992 55956 23004
rect 56008 22992 56014 23044
rect 50706 22964 50712 22976
rect 48240 22936 50712 22964
rect 43441 22927 43499 22933
rect 50706 22924 50712 22936
rect 50764 22924 50770 22976
rect 53374 22964 53380 22976
rect 53335 22936 53380 22964
rect 53374 22924 53380 22936
rect 53432 22924 53438 22976
rect 53926 22924 53932 22976
rect 53984 22964 53990 22976
rect 55122 22964 55128 22976
rect 53984 22936 55128 22964
rect 53984 22924 53990 22936
rect 55122 22924 55128 22936
rect 55180 22964 55186 22976
rect 56152 22964 56180 23063
rect 56318 23060 56324 23112
rect 56376 23109 56382 23112
rect 57146 23109 57152 23112
rect 56376 23100 56384 23109
rect 57140 23100 57152 23109
rect 56376 23072 56421 23100
rect 57107 23072 57152 23100
rect 56376 23063 56384 23072
rect 57140 23063 57152 23072
rect 56376 23060 56382 23063
rect 57146 23060 57152 23063
rect 57204 23060 57210 23112
rect 56229 23035 56287 23041
rect 56229 23001 56241 23035
rect 56275 23032 56287 23035
rect 57514 23032 57520 23044
rect 56275 23004 57520 23032
rect 56275 23001 56287 23004
rect 56229 22995 56287 23001
rect 57514 22992 57520 23004
rect 57572 22992 57578 23044
rect 55180 22936 56180 22964
rect 55180 22924 55186 22936
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 17310 22720 17316 22772
rect 17368 22760 17374 22772
rect 17494 22760 17500 22772
rect 17368 22732 17500 22760
rect 17368 22720 17374 22732
rect 17494 22720 17500 22732
rect 17552 22720 17558 22772
rect 19426 22720 19432 22772
rect 19484 22760 19490 22772
rect 23842 22760 23848 22772
rect 19484 22732 23704 22760
rect 23803 22732 23848 22760
rect 19484 22720 19490 22732
rect 19334 22692 19340 22704
rect 17052 22664 19340 22692
rect 1581 22627 1639 22633
rect 1581 22593 1593 22627
rect 1627 22624 1639 22627
rect 13538 22624 13544 22636
rect 1627 22596 13544 22624
rect 1627 22593 1639 22596
rect 1581 22587 1639 22593
rect 13538 22584 13544 22596
rect 13596 22584 13602 22636
rect 17052 22633 17080 22664
rect 17512 22636 17540 22664
rect 19334 22652 19340 22664
rect 19392 22652 19398 22704
rect 20346 22652 20352 22704
rect 20404 22692 20410 22704
rect 21177 22695 21235 22701
rect 21177 22692 21189 22695
rect 20404 22664 21189 22692
rect 20404 22652 20410 22664
rect 21177 22661 21189 22664
rect 21223 22692 21235 22695
rect 22732 22695 22790 22701
rect 21223 22664 22094 22692
rect 21223 22661 21235 22664
rect 21177 22655 21235 22661
rect 17037 22627 17095 22633
rect 17037 22593 17049 22627
rect 17083 22593 17095 22627
rect 17037 22587 17095 22593
rect 17405 22627 17463 22633
rect 17405 22593 17417 22627
rect 17451 22593 17463 22627
rect 17405 22587 17463 22593
rect 1762 22556 1768 22568
rect 1723 22528 1768 22556
rect 1762 22516 1768 22528
rect 1820 22516 1826 22568
rect 17420 22556 17448 22587
rect 17494 22584 17500 22636
rect 17552 22584 17558 22636
rect 17678 22584 17684 22636
rect 17736 22624 17742 22636
rect 17773 22627 17831 22633
rect 17773 22624 17785 22627
rect 17736 22596 17785 22624
rect 17736 22584 17742 22596
rect 17773 22593 17785 22596
rect 17819 22624 17831 22627
rect 17862 22624 17868 22636
rect 17819 22596 17868 22624
rect 17819 22593 17831 22596
rect 17773 22587 17831 22593
rect 17862 22584 17868 22596
rect 17920 22584 17926 22636
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22624 18475 22627
rect 18874 22624 18880 22636
rect 18463 22596 18880 22624
rect 18463 22593 18475 22596
rect 18417 22587 18475 22593
rect 18874 22584 18880 22596
rect 18932 22584 18938 22636
rect 21358 22624 21364 22636
rect 21319 22596 21364 22624
rect 21358 22584 21364 22596
rect 21416 22584 21422 22636
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22624 21511 22627
rect 21818 22624 21824 22636
rect 21499 22596 21824 22624
rect 21499 22593 21511 22596
rect 21453 22587 21511 22593
rect 18230 22556 18236 22568
rect 17420 22528 18236 22556
rect 18230 22516 18236 22528
rect 18288 22516 18294 22568
rect 20530 22516 20536 22568
rect 20588 22556 20594 22568
rect 21468 22556 21496 22587
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 22066 22624 22094 22664
rect 22732 22661 22744 22695
rect 22778 22692 22790 22695
rect 22922 22692 22928 22704
rect 22778 22664 22928 22692
rect 22778 22661 22790 22664
rect 22732 22655 22790 22661
rect 22922 22652 22928 22664
rect 22980 22652 22986 22704
rect 23676 22692 23704 22732
rect 23842 22720 23848 22732
rect 23900 22720 23906 22772
rect 24578 22720 24584 22772
rect 24636 22760 24642 22772
rect 25501 22763 25559 22769
rect 25501 22760 25513 22763
rect 24636 22732 25513 22760
rect 24636 22720 24642 22732
rect 25501 22729 25513 22732
rect 25547 22729 25559 22763
rect 25501 22723 25559 22729
rect 26234 22720 26240 22772
rect 26292 22760 26298 22772
rect 26418 22760 26424 22772
rect 26292 22732 26424 22760
rect 26292 22720 26298 22732
rect 26418 22720 26424 22732
rect 26476 22760 26482 22772
rect 27062 22760 27068 22772
rect 26476 22732 27068 22760
rect 26476 22720 26482 22732
rect 27062 22720 27068 22732
rect 27120 22720 27126 22772
rect 29362 22720 29368 22772
rect 29420 22760 29426 22772
rect 31018 22760 31024 22772
rect 29420 22732 31024 22760
rect 29420 22720 29426 22732
rect 31018 22720 31024 22732
rect 31076 22720 31082 22772
rect 34698 22720 34704 22772
rect 34756 22760 34762 22772
rect 35069 22763 35127 22769
rect 35069 22760 35081 22763
rect 34756 22732 35081 22760
rect 34756 22720 34762 22732
rect 35069 22729 35081 22732
rect 35115 22729 35127 22763
rect 35618 22760 35624 22772
rect 35069 22723 35127 22729
rect 35314 22732 35624 22760
rect 28994 22692 29000 22704
rect 23676 22664 29000 22692
rect 28994 22652 29000 22664
rect 29052 22652 29058 22704
rect 23290 22624 23296 22636
rect 22066 22596 23296 22624
rect 23290 22584 23296 22596
rect 23348 22624 23354 22636
rect 24302 22624 24308 22636
rect 23348 22596 23888 22624
rect 24263 22596 24308 22624
rect 23348 22584 23354 22596
rect 20588 22528 21496 22556
rect 20588 22516 20594 22528
rect 22370 22516 22376 22568
rect 22428 22556 22434 22568
rect 22465 22559 22523 22565
rect 22465 22556 22477 22559
rect 22428 22528 22477 22556
rect 22428 22516 22434 22528
rect 22465 22525 22477 22528
rect 22511 22525 22523 22559
rect 22465 22519 22523 22525
rect 17954 22380 17960 22432
rect 18012 22420 18018 22432
rect 19613 22423 19671 22429
rect 19613 22420 19625 22423
rect 18012 22392 19625 22420
rect 18012 22380 18018 22392
rect 19613 22389 19625 22392
rect 19659 22389 19671 22423
rect 19613 22383 19671 22389
rect 21177 22423 21235 22429
rect 21177 22389 21189 22423
rect 21223 22420 21235 22423
rect 23566 22420 23572 22432
rect 21223 22392 23572 22420
rect 21223 22389 21235 22392
rect 21177 22383 21235 22389
rect 23566 22380 23572 22392
rect 23624 22380 23630 22432
rect 23860 22420 23888 22596
rect 24302 22584 24308 22596
rect 24360 22584 24366 22636
rect 27430 22624 27436 22636
rect 27391 22596 27436 22624
rect 27430 22584 27436 22596
rect 27488 22584 27494 22636
rect 27706 22624 27712 22636
rect 27667 22596 27712 22624
rect 27706 22584 27712 22596
rect 27764 22584 27770 22636
rect 27982 22624 27988 22636
rect 27943 22596 27988 22624
rect 27982 22584 27988 22596
rect 28040 22584 28046 22636
rect 28350 22624 28356 22636
rect 28311 22596 28356 22624
rect 28350 22584 28356 22596
rect 28408 22624 28414 22636
rect 28534 22624 28540 22636
rect 28408 22596 28540 22624
rect 28408 22584 28414 22596
rect 28534 22584 28540 22596
rect 28592 22584 28598 22636
rect 29457 22627 29515 22633
rect 29457 22593 29469 22627
rect 29503 22624 29515 22627
rect 29638 22624 29644 22636
rect 29503 22596 29644 22624
rect 29503 22593 29515 22596
rect 29457 22587 29515 22593
rect 29638 22584 29644 22596
rect 29696 22584 29702 22636
rect 30374 22584 30380 22636
rect 30432 22624 30438 22636
rect 30834 22624 30840 22636
rect 30432 22596 30840 22624
rect 30432 22584 30438 22596
rect 30834 22584 30840 22596
rect 30892 22624 30898 22636
rect 32309 22627 32367 22633
rect 32309 22624 32321 22627
rect 30892 22596 32321 22624
rect 30892 22584 30898 22596
rect 32309 22593 32321 22596
rect 32355 22593 32367 22627
rect 32309 22587 32367 22593
rect 34054 22584 34060 22636
rect 34112 22624 34118 22636
rect 35314 22633 35342 22732
rect 35618 22720 35624 22732
rect 35676 22720 35682 22772
rect 35710 22720 35716 22772
rect 35768 22760 35774 22772
rect 35894 22760 35900 22772
rect 35768 22732 35900 22760
rect 35768 22720 35774 22732
rect 35894 22720 35900 22732
rect 35952 22720 35958 22772
rect 36262 22760 36268 22772
rect 36223 22732 36268 22760
rect 36262 22720 36268 22732
rect 36320 22720 36326 22772
rect 36630 22720 36636 22772
rect 36688 22720 36694 22772
rect 36722 22720 36728 22772
rect 36780 22760 36786 22772
rect 37826 22760 37832 22772
rect 36780 22720 36789 22760
rect 37787 22732 37832 22760
rect 37826 22720 37832 22732
rect 37884 22720 37890 22772
rect 40310 22760 40316 22772
rect 40271 22732 40316 22760
rect 40310 22720 40316 22732
rect 40368 22720 40374 22772
rect 43254 22720 43260 22772
rect 43312 22760 43318 22772
rect 44726 22760 44732 22772
rect 43312 22732 44732 22760
rect 43312 22720 43318 22732
rect 44726 22720 44732 22732
rect 44784 22720 44790 22772
rect 45554 22720 45560 22772
rect 45612 22760 45618 22772
rect 45830 22760 45836 22772
rect 45612 22732 45836 22760
rect 45612 22720 45618 22732
rect 45830 22720 45836 22732
rect 45888 22720 45894 22772
rect 49142 22760 49148 22772
rect 49103 22732 49148 22760
rect 49142 22720 49148 22732
rect 49200 22720 49206 22772
rect 36648 22692 36676 22720
rect 36510 22664 36676 22692
rect 35299 22627 35357 22633
rect 35299 22624 35311 22627
rect 34112 22596 35311 22624
rect 34112 22584 34118 22596
rect 35299 22593 35311 22596
rect 35345 22593 35357 22627
rect 35299 22587 35357 22593
rect 35437 22627 35495 22633
rect 35437 22593 35449 22627
rect 35483 22593 35495 22627
rect 35437 22587 35495 22593
rect 35529 22627 35587 22633
rect 35529 22593 35541 22627
rect 35575 22624 35587 22627
rect 35618 22624 35624 22636
rect 35575 22596 35624 22624
rect 35575 22593 35587 22596
rect 35529 22587 35587 22593
rect 27617 22559 27675 22565
rect 27617 22525 27629 22559
rect 27663 22556 27675 22559
rect 33594 22556 33600 22568
rect 27663 22528 33600 22556
rect 27663 22525 27675 22528
rect 27617 22519 27675 22525
rect 33594 22516 33600 22528
rect 33652 22516 33658 22568
rect 35452 22556 35480 22587
rect 35618 22584 35624 22596
rect 35676 22584 35682 22636
rect 35713 22627 35771 22633
rect 35713 22593 35725 22627
rect 35759 22624 35771 22627
rect 36078 22624 36084 22636
rect 35759 22596 36084 22624
rect 35759 22593 35771 22596
rect 35713 22587 35771 22593
rect 36078 22584 36084 22596
rect 36136 22584 36142 22636
rect 36262 22584 36268 22636
rect 36320 22624 36326 22636
rect 36510 22633 36538 22664
rect 36761 22639 36789 22720
rect 37550 22652 37556 22704
rect 37608 22692 37614 22704
rect 37645 22695 37703 22701
rect 37645 22692 37657 22695
rect 37608 22664 37657 22692
rect 37608 22652 37614 22664
rect 37645 22661 37657 22664
rect 37691 22661 37703 22695
rect 37645 22655 37703 22661
rect 38930 22652 38936 22704
rect 38988 22692 38994 22704
rect 40402 22692 40408 22704
rect 38988 22664 40408 22692
rect 38988 22652 38994 22664
rect 40402 22652 40408 22664
rect 40460 22652 40466 22704
rect 40586 22652 40592 22704
rect 40644 22692 40650 22704
rect 48130 22692 48136 22704
rect 40644 22664 48136 22692
rect 40644 22652 40650 22664
rect 48130 22652 48136 22664
rect 48188 22652 48194 22704
rect 36746 22633 36804 22639
rect 36510 22627 36579 22633
rect 36510 22624 36533 22627
rect 36320 22596 36533 22624
rect 36320 22584 36326 22596
rect 36521 22593 36533 22596
rect 36567 22593 36579 22627
rect 36521 22587 36579 22593
rect 36633 22627 36691 22633
rect 36633 22593 36645 22627
rect 36679 22593 36691 22627
rect 36746 22599 36758 22633
rect 36792 22599 36804 22633
rect 36746 22593 36804 22599
rect 36633 22587 36691 22593
rect 35433 22528 35480 22556
rect 27246 22448 27252 22500
rect 27304 22488 27310 22500
rect 30374 22488 30380 22500
rect 27304 22460 30380 22488
rect 27304 22448 27310 22460
rect 30374 22448 30380 22460
rect 30432 22448 30438 22500
rect 30466 22448 30472 22500
rect 30524 22488 30530 22500
rect 30524 22460 30788 22488
rect 30524 22448 30530 22460
rect 30653 22423 30711 22429
rect 30653 22420 30665 22423
rect 23860 22392 30665 22420
rect 30653 22389 30665 22392
rect 30699 22389 30711 22423
rect 30760 22420 30788 22460
rect 33134 22448 33140 22500
rect 33192 22488 33198 22500
rect 35433 22488 35461 22528
rect 36648 22488 36676 22587
rect 36906 22584 36912 22636
rect 36964 22624 36970 22636
rect 37458 22624 37464 22636
rect 36964 22596 37009 22624
rect 37419 22596 37464 22624
rect 36964 22584 36970 22596
rect 37458 22584 37464 22596
rect 37516 22584 37522 22636
rect 39022 22584 39028 22636
rect 39080 22624 39086 22636
rect 39189 22627 39247 22633
rect 39189 22624 39201 22627
rect 39080 22596 39201 22624
rect 39080 22584 39086 22596
rect 39189 22593 39201 22596
rect 39235 22593 39247 22627
rect 43806 22624 43812 22636
rect 43767 22596 43812 22624
rect 39189 22587 39247 22593
rect 43806 22584 43812 22596
rect 43864 22584 43870 22636
rect 43993 22627 44051 22633
rect 43993 22593 44005 22627
rect 44039 22593 44051 22627
rect 43993 22587 44051 22593
rect 44453 22627 44511 22633
rect 44453 22593 44465 22627
rect 44499 22624 44511 22627
rect 44542 22624 44548 22636
rect 44499 22596 44548 22624
rect 44499 22593 44511 22596
rect 44453 22587 44511 22593
rect 37182 22516 37188 22568
rect 37240 22556 37246 22568
rect 38930 22556 38936 22568
rect 37240 22528 38936 22556
rect 37240 22516 37246 22528
rect 38930 22516 38936 22528
rect 38988 22516 38994 22568
rect 43162 22516 43168 22568
rect 43220 22556 43226 22568
rect 44008 22556 44036 22587
rect 44542 22584 44548 22596
rect 44600 22584 44606 22636
rect 44726 22633 44732 22636
rect 44720 22587 44732 22633
rect 44784 22624 44790 22636
rect 48032 22627 48090 22633
rect 44784 22596 44820 22624
rect 44726 22584 44732 22587
rect 44784 22584 44790 22596
rect 48032 22593 48044 22627
rect 48078 22624 48090 22627
rect 48866 22624 48872 22636
rect 48078 22596 48872 22624
rect 48078 22593 48090 22596
rect 48032 22587 48090 22593
rect 48866 22584 48872 22596
rect 48924 22584 48930 22636
rect 56502 22624 56508 22636
rect 56463 22596 56508 22624
rect 56502 22584 56508 22596
rect 56560 22584 56566 22636
rect 56689 22627 56747 22633
rect 56689 22593 56701 22627
rect 56735 22624 56747 22627
rect 56778 22624 56784 22636
rect 56735 22596 56784 22624
rect 56735 22593 56747 22596
rect 56689 22587 56747 22593
rect 56778 22584 56784 22596
rect 56836 22584 56842 22636
rect 58066 22624 58072 22636
rect 58027 22596 58072 22624
rect 58066 22584 58072 22596
rect 58124 22584 58130 22636
rect 43220 22528 44036 22556
rect 47765 22559 47823 22565
rect 43220 22516 43226 22528
rect 47765 22525 47777 22559
rect 47811 22525 47823 22559
rect 47765 22519 47823 22525
rect 43714 22488 43720 22500
rect 33192 22460 36676 22488
rect 39868 22460 43720 22488
rect 33192 22448 33198 22460
rect 34624 22432 34652 22460
rect 33505 22423 33563 22429
rect 33505 22420 33517 22423
rect 30760 22392 33517 22420
rect 30653 22383 30711 22389
rect 33505 22389 33517 22392
rect 33551 22389 33563 22423
rect 33505 22383 33563 22389
rect 34606 22380 34612 22432
rect 34664 22380 34670 22432
rect 35894 22380 35900 22432
rect 35952 22420 35958 22432
rect 36170 22420 36176 22432
rect 35952 22392 36176 22420
rect 35952 22380 35958 22392
rect 36170 22380 36176 22392
rect 36228 22380 36234 22432
rect 36446 22380 36452 22432
rect 36504 22420 36510 22432
rect 39868 22420 39896 22460
rect 43714 22448 43720 22460
rect 43772 22448 43778 22500
rect 36504 22392 39896 22420
rect 43809 22423 43867 22429
rect 36504 22380 36510 22392
rect 43809 22389 43821 22423
rect 43855 22420 43867 22423
rect 44266 22420 44272 22432
rect 43855 22392 44272 22420
rect 43855 22389 43867 22392
rect 43809 22383 43867 22389
rect 44266 22380 44272 22392
rect 44324 22380 44330 22432
rect 47780 22420 47808 22519
rect 56410 22448 56416 22500
rect 56468 22488 56474 22500
rect 56505 22491 56563 22497
rect 56505 22488 56517 22491
rect 56468 22460 56517 22488
rect 56468 22448 56474 22460
rect 56505 22457 56517 22460
rect 56551 22457 56563 22491
rect 56505 22451 56563 22457
rect 48130 22420 48136 22432
rect 47780 22392 48136 22420
rect 48130 22380 48136 22392
rect 48188 22380 48194 22432
rect 56318 22380 56324 22432
rect 56376 22420 56382 22432
rect 58253 22423 58311 22429
rect 58253 22420 58265 22423
rect 56376 22392 58265 22420
rect 56376 22380 56382 22392
rect 58253 22389 58265 22392
rect 58299 22389 58311 22423
rect 58253 22383 58311 22389
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 13538 22216 13544 22228
rect 13499 22188 13544 22216
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 14274 22176 14280 22228
rect 14332 22216 14338 22228
rect 16850 22216 16856 22228
rect 14332 22188 16856 22216
rect 14332 22176 14338 22188
rect 16850 22176 16856 22188
rect 16908 22216 16914 22228
rect 53374 22216 53380 22228
rect 16908 22188 53380 22216
rect 16908 22176 16914 22188
rect 53374 22176 53380 22188
rect 53432 22176 53438 22228
rect 26970 22108 26976 22160
rect 27028 22148 27034 22160
rect 27982 22148 27988 22160
rect 27028 22120 27988 22148
rect 27028 22108 27034 22120
rect 27982 22108 27988 22120
rect 28040 22108 28046 22160
rect 31478 22148 31484 22160
rect 30208 22120 31484 22148
rect 24394 22080 24400 22092
rect 20456 22052 24400 22080
rect 13354 22012 13360 22024
rect 13315 21984 13360 22012
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 13511 22015 13569 22021
rect 13511 21981 13523 22015
rect 13557 22012 13569 22015
rect 14366 22012 14372 22024
rect 13557 21984 14228 22012
rect 14327 21984 14372 22012
rect 13557 21981 13569 21984
rect 13511 21975 13569 21981
rect 14200 21944 14228 21984
rect 14366 21972 14372 21984
rect 14424 21972 14430 22024
rect 16577 22015 16635 22021
rect 16577 21981 16589 22015
rect 16623 22012 16635 22015
rect 16666 22012 16672 22024
rect 16623 21984 16672 22012
rect 16623 21981 16635 21984
rect 16577 21975 16635 21981
rect 16666 21972 16672 21984
rect 16724 21972 16730 22024
rect 19426 22012 19432 22024
rect 19387 21984 19432 22012
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 20456 22012 20484 22052
rect 24394 22040 24400 22052
rect 24452 22040 24458 22092
rect 29730 22040 29736 22092
rect 29788 22080 29794 22092
rect 30208 22080 30236 22120
rect 31478 22108 31484 22120
rect 31536 22148 31542 22160
rect 33134 22148 33140 22160
rect 31536 22120 33140 22148
rect 31536 22108 31542 22120
rect 33134 22108 33140 22120
rect 33192 22108 33198 22160
rect 34146 22148 34152 22160
rect 34107 22120 34152 22148
rect 34146 22108 34152 22120
rect 34204 22108 34210 22160
rect 37090 22148 37096 22160
rect 37051 22120 37096 22148
rect 37090 22108 37096 22120
rect 37148 22108 37154 22160
rect 40034 22108 40040 22160
rect 40092 22148 40098 22160
rect 44361 22151 44419 22157
rect 44361 22148 44373 22151
rect 40092 22120 44373 22148
rect 40092 22108 40098 22120
rect 44361 22117 44373 22120
rect 44407 22117 44419 22151
rect 44361 22111 44419 22117
rect 45189 22151 45247 22157
rect 45189 22117 45201 22151
rect 45235 22117 45247 22151
rect 45189 22111 45247 22117
rect 30650 22080 30656 22092
rect 29788 22052 30236 22080
rect 29788 22040 29794 22052
rect 19536 21984 20484 22012
rect 21729 22015 21787 22021
rect 14921 21947 14979 21953
rect 14921 21944 14933 21947
rect 14200 21916 14933 21944
rect 14921 21913 14933 21916
rect 14967 21944 14979 21947
rect 19536 21944 19564 21984
rect 21729 21981 21741 22015
rect 21775 22012 21787 22015
rect 22278 22012 22284 22024
rect 21775 21984 22284 22012
rect 21775 21981 21787 21984
rect 21729 21975 21787 21981
rect 22278 21972 22284 21984
rect 22336 21972 22342 22024
rect 22370 21972 22376 22024
rect 22428 22012 22434 22024
rect 24581 22015 24639 22021
rect 24581 22012 24593 22015
rect 22428 21984 24593 22012
rect 22428 21972 22434 21984
rect 24581 21981 24593 21984
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 25130 21972 25136 22024
rect 25188 22012 25194 22024
rect 25188 21984 26832 22012
rect 25188 21972 25194 21984
rect 14967 21916 19564 21944
rect 19696 21947 19754 21953
rect 14967 21913 14979 21916
rect 14921 21907 14979 21913
rect 19696 21913 19708 21947
rect 19742 21944 19754 21947
rect 20714 21944 20720 21956
rect 19742 21916 20720 21944
rect 19742 21913 19754 21916
rect 19696 21907 19754 21913
rect 20714 21904 20720 21916
rect 20772 21904 20778 21956
rect 24848 21947 24906 21953
rect 24848 21913 24860 21947
rect 24894 21944 24906 21947
rect 26510 21944 26516 21956
rect 24894 21916 26516 21944
rect 24894 21913 24906 21916
rect 24848 21907 24906 21913
rect 26510 21904 26516 21916
rect 26568 21904 26574 21956
rect 26804 21944 26832 21984
rect 26878 21972 26884 22024
rect 26936 22012 26942 22024
rect 26936 21984 26981 22012
rect 26936 21972 26942 21984
rect 29270 21972 29276 22024
rect 29328 22012 29334 22024
rect 30006 22012 30012 22024
rect 29328 21984 30012 22012
rect 29328 21972 29334 21984
rect 30006 21972 30012 21984
rect 30064 22021 30070 22024
rect 30208 22021 30236 22052
rect 30392 22052 30656 22080
rect 30064 22015 30113 22021
rect 30064 21981 30067 22015
rect 30101 21981 30113 22015
rect 30064 21975 30113 21981
rect 30193 22015 30251 22021
rect 30193 21981 30205 22015
rect 30239 21981 30251 22015
rect 30193 21975 30251 21981
rect 30306 22015 30364 22021
rect 30306 21981 30318 22015
rect 30352 22012 30364 22015
rect 30392 22012 30420 22052
rect 30650 22040 30656 22052
rect 30708 22040 30714 22092
rect 31110 22040 31116 22092
rect 31168 22080 31174 22092
rect 34885 22083 34943 22089
rect 31168 22052 33364 22080
rect 31168 22040 31174 22052
rect 30352 21984 30420 22012
rect 30469 22015 30527 22021
rect 30352 21981 30364 21984
rect 30306 21975 30364 21981
rect 30469 21981 30481 22015
rect 30515 21981 30527 22015
rect 30469 21975 30527 21981
rect 30064 21972 30070 21975
rect 30484 21944 30512 21975
rect 30926 21972 30932 22024
rect 30984 22012 30990 22024
rect 31021 22015 31079 22021
rect 31021 22012 31033 22015
rect 30984 21984 31033 22012
rect 30984 21972 30990 21984
rect 31021 21981 31033 21984
rect 31067 22012 31079 22015
rect 31570 22012 31576 22024
rect 31067 21984 31576 22012
rect 31067 21981 31079 21984
rect 31021 21975 31079 21981
rect 31570 21972 31576 21984
rect 31628 21972 31634 22024
rect 33336 22012 33364 22052
rect 34885 22049 34897 22083
rect 34931 22080 34943 22083
rect 36538 22080 36544 22092
rect 34931 22052 36544 22080
rect 34931 22049 34943 22052
rect 34885 22043 34943 22049
rect 36538 22040 36544 22052
rect 36596 22080 36602 22092
rect 37182 22080 37188 22092
rect 36596 22052 37188 22080
rect 36596 22040 36602 22052
rect 37182 22040 37188 22052
rect 37240 22040 37246 22092
rect 37277 22083 37335 22089
rect 37277 22049 37289 22083
rect 37323 22049 37335 22083
rect 39114 22080 39120 22092
rect 39075 22052 39120 22080
rect 37277 22043 37335 22049
rect 33962 22021 33968 22024
rect 33954 22015 33968 22021
rect 33954 22012 33966 22015
rect 33336 21984 33966 22012
rect 33954 21981 33966 21984
rect 33954 21975 33968 21981
rect 33962 21972 33968 21975
rect 34020 21972 34026 22024
rect 35161 22015 35219 22021
rect 35161 21981 35173 22015
rect 35207 22012 35219 22015
rect 35434 22012 35440 22024
rect 35207 21984 35440 22012
rect 35207 21981 35219 21984
rect 35161 21975 35219 21981
rect 35434 21972 35440 21984
rect 35492 21972 35498 22024
rect 35618 21972 35624 22024
rect 35676 22012 35682 22024
rect 37001 22015 37059 22021
rect 37001 22012 37013 22015
rect 35676 21984 37013 22012
rect 35676 21972 35682 21984
rect 37001 21981 37013 21984
rect 37047 21981 37059 22015
rect 37292 22012 37320 22043
rect 39114 22040 39120 22052
rect 39172 22040 39178 22092
rect 45204 22080 45232 22111
rect 45370 22108 45376 22160
rect 45428 22148 45434 22160
rect 45741 22151 45799 22157
rect 45741 22148 45753 22151
rect 45428 22120 45753 22148
rect 45428 22108 45434 22120
rect 45741 22117 45753 22120
rect 45787 22148 45799 22151
rect 46109 22151 46167 22157
rect 46109 22148 46121 22151
rect 45787 22120 46121 22148
rect 45787 22117 45799 22120
rect 45741 22111 45799 22117
rect 46109 22117 46121 22120
rect 46155 22117 46167 22151
rect 49142 22148 49148 22160
rect 46109 22111 46167 22117
rect 48286 22120 49148 22148
rect 43180 22052 45232 22080
rect 37458 22012 37464 22024
rect 37001 21975 37059 21981
rect 37108 21984 37464 22012
rect 31754 21944 31760 21956
rect 26804 21916 28120 21944
rect 30484 21916 31760 21944
rect 15930 21836 15936 21888
rect 15988 21876 15994 21888
rect 16206 21876 16212 21888
rect 15988 21848 16212 21876
rect 15988 21836 15994 21848
rect 16206 21836 16212 21848
rect 16264 21836 16270 21888
rect 16574 21836 16580 21888
rect 16632 21876 16638 21888
rect 17773 21879 17831 21885
rect 17773 21876 17785 21879
rect 16632 21848 17785 21876
rect 16632 21836 16638 21848
rect 17773 21845 17785 21848
rect 17819 21845 17831 21879
rect 17773 21839 17831 21845
rect 20809 21879 20867 21885
rect 20809 21845 20821 21879
rect 20855 21876 20867 21879
rect 22002 21876 22008 21888
rect 20855 21848 22008 21876
rect 20855 21845 20867 21848
rect 20809 21839 20867 21845
rect 22002 21836 22008 21848
rect 22060 21836 22066 21888
rect 22922 21876 22928 21888
rect 22883 21848 22928 21876
rect 22922 21836 22928 21848
rect 22980 21836 22986 21888
rect 25961 21879 26019 21885
rect 25961 21845 25973 21879
rect 26007 21876 26019 21879
rect 27246 21876 27252 21888
rect 26007 21848 27252 21876
rect 26007 21845 26019 21848
rect 25961 21839 26019 21845
rect 27246 21836 27252 21848
rect 27304 21836 27310 21888
rect 28092 21885 28120 21916
rect 31754 21904 31760 21916
rect 31812 21904 31818 21956
rect 33781 21947 33839 21953
rect 33781 21913 33793 21947
rect 33827 21944 33839 21947
rect 34146 21944 34152 21956
rect 33827 21916 34152 21944
rect 33827 21913 33839 21916
rect 33781 21907 33839 21913
rect 33888 21888 33916 21916
rect 34146 21904 34152 21916
rect 34204 21904 34210 21956
rect 36538 21904 36544 21956
rect 36596 21944 36602 21956
rect 37108 21944 37136 21984
rect 37458 21972 37464 21984
rect 37516 22012 37522 22024
rect 37921 22015 37979 22021
rect 37921 22012 37933 22015
rect 37516 21984 37933 22012
rect 37516 21972 37522 21984
rect 37921 21981 37933 21984
rect 37967 21981 37979 22015
rect 38102 22012 38108 22024
rect 38063 21984 38108 22012
rect 37921 21975 37979 21981
rect 38102 21972 38108 21984
rect 38160 21972 38166 22024
rect 38838 22012 38844 22024
rect 38799 21984 38844 22012
rect 38838 21972 38844 21984
rect 38896 21972 38902 22024
rect 38933 22015 38991 22021
rect 38933 21981 38945 22015
rect 38979 22012 38991 22015
rect 39666 22012 39672 22024
rect 38979 21984 39672 22012
rect 38979 21981 38991 21984
rect 38933 21975 38991 21981
rect 39666 21972 39672 21984
rect 39724 21972 39730 22024
rect 40034 21972 40040 22024
rect 40092 22012 40098 22024
rect 40310 22012 40316 22024
rect 40092 21984 40137 22012
rect 40271 21984 40316 22012
rect 40092 21972 40098 21984
rect 40310 21972 40316 21984
rect 40368 22012 40374 22024
rect 40586 22012 40592 22024
rect 40368 21984 40592 22012
rect 40368 21972 40374 21984
rect 40586 21972 40592 21984
rect 40644 21972 40650 22024
rect 43180 22021 43208 22052
rect 43165 22015 43223 22021
rect 43165 21981 43177 22015
rect 43211 21981 43223 22015
rect 43165 21975 43223 21981
rect 43346 21972 43352 22024
rect 43404 22012 43410 22024
rect 43404 21984 43449 22012
rect 43404 21972 43410 21984
rect 43990 21972 43996 22024
rect 44048 22012 44054 22024
rect 44048 21984 44090 22012
rect 44048 21972 44054 21984
rect 44358 21972 44364 22024
rect 44416 22012 44422 22024
rect 44453 22015 44511 22021
rect 44453 22012 44465 22015
rect 44416 21984 44465 22012
rect 44416 21972 44422 21984
rect 44453 21981 44465 21984
rect 44499 21981 44511 22015
rect 44453 21975 44511 21981
rect 45370 22015 45428 22021
rect 45370 21981 45382 22015
rect 45416 22012 45428 22015
rect 45554 22012 45560 22024
rect 45416 21984 45560 22012
rect 45416 21981 45428 21984
rect 45370 21975 45428 21981
rect 37274 21944 37280 21956
rect 36596 21916 37136 21944
rect 37235 21916 37280 21944
rect 36596 21904 36602 21916
rect 37274 21904 37280 21916
rect 37332 21904 37338 21956
rect 38289 21947 38347 21953
rect 38289 21913 38301 21947
rect 38335 21944 38347 21947
rect 39482 21944 39488 21956
rect 38335 21916 39488 21944
rect 38335 21913 38347 21916
rect 38289 21907 38347 21913
rect 39482 21904 39488 21916
rect 39540 21904 39546 21956
rect 43254 21944 43260 21956
rect 43215 21916 43260 21944
rect 43254 21904 43260 21916
rect 43312 21904 43318 21956
rect 44468 21944 44496 21975
rect 45554 21972 45560 21984
rect 45612 21972 45618 22024
rect 45833 22015 45891 22021
rect 45833 21981 45845 22015
rect 45879 21981 45891 22015
rect 47486 22012 47492 22024
rect 47447 21984 47492 22012
rect 45833 21975 45891 21981
rect 45848 21944 45876 21975
rect 47486 21972 47492 21984
rect 47544 21972 47550 22024
rect 47854 22012 47860 22024
rect 47815 21984 47860 22012
rect 47854 21972 47860 21984
rect 47912 21972 47918 22024
rect 44468 21916 45876 21944
rect 47673 21947 47731 21953
rect 47673 21913 47685 21947
rect 47719 21913 47731 21947
rect 47673 21907 47731 21913
rect 47765 21947 47823 21953
rect 47765 21913 47777 21947
rect 47811 21944 47823 21947
rect 48286 21944 48314 22120
rect 49142 22108 49148 22120
rect 49200 22108 49206 22160
rect 48866 22080 48872 22092
rect 48827 22052 48872 22080
rect 48866 22040 48872 22052
rect 48924 22040 48930 22092
rect 51626 22040 51632 22092
rect 51684 22080 51690 22092
rect 53926 22080 53932 22092
rect 51684 22052 53932 22080
rect 51684 22040 51690 22052
rect 53926 22040 53932 22052
rect 53984 22040 53990 22092
rect 48498 22012 48504 22024
rect 48459 21984 48504 22012
rect 48498 21972 48504 21984
rect 48556 21972 48562 22024
rect 48685 22015 48743 22021
rect 48685 21981 48697 22015
rect 48731 21981 48743 22015
rect 48685 21975 48743 21981
rect 47811 21916 48314 21944
rect 47811 21913 47823 21916
rect 47765 21907 47823 21913
rect 28077 21879 28135 21885
rect 28077 21845 28089 21879
rect 28123 21845 28135 21879
rect 29822 21876 29828 21888
rect 29783 21848 29828 21876
rect 28077 21839 28135 21845
rect 29822 21836 29828 21848
rect 29880 21836 29886 21888
rect 30190 21836 30196 21888
rect 30248 21876 30254 21888
rect 32217 21879 32275 21885
rect 32217 21876 32229 21879
rect 30248 21848 32229 21876
rect 30248 21836 30254 21848
rect 32217 21845 32229 21848
rect 32263 21845 32275 21879
rect 32217 21839 32275 21845
rect 33870 21836 33876 21888
rect 33928 21836 33934 21888
rect 34330 21836 34336 21888
rect 34388 21876 34394 21888
rect 36265 21879 36323 21885
rect 36265 21876 36277 21879
rect 34388 21848 36277 21876
rect 34388 21836 34394 21848
rect 36265 21845 36277 21848
rect 36311 21845 36323 21879
rect 43806 21876 43812 21888
rect 43767 21848 43812 21876
rect 36265 21839 36323 21845
rect 43806 21836 43812 21848
rect 43864 21836 43870 21888
rect 43898 21836 43904 21888
rect 43956 21876 43962 21888
rect 43993 21879 44051 21885
rect 43993 21876 44005 21879
rect 43956 21848 44005 21876
rect 43956 21836 43962 21848
rect 43993 21845 44005 21848
rect 44039 21876 44051 21879
rect 45373 21879 45431 21885
rect 45373 21876 45385 21879
rect 44039 21848 45385 21876
rect 44039 21845 44051 21848
rect 43993 21839 44051 21845
rect 45373 21845 45385 21848
rect 45419 21845 45431 21879
rect 47688 21876 47716 21907
rect 47854 21876 47860 21888
rect 47688 21848 47860 21876
rect 45373 21839 45431 21845
rect 47854 21836 47860 21848
rect 47912 21836 47918 21888
rect 48041 21879 48099 21885
rect 48041 21845 48053 21879
rect 48087 21876 48099 21879
rect 48700 21876 48728 21975
rect 51718 21972 51724 22024
rect 51776 22012 51782 22024
rect 57885 22015 57943 22021
rect 57885 22012 57897 22015
rect 51776 21984 57897 22012
rect 51776 21972 51782 21984
rect 57885 21981 57897 21984
rect 57931 21981 57943 22015
rect 57885 21975 57943 21981
rect 58158 21944 58164 21956
rect 58119 21916 58164 21944
rect 58158 21904 58164 21916
rect 58216 21904 58222 21956
rect 48087 21848 48728 21876
rect 48087 21845 48099 21848
rect 48041 21839 48099 21845
rect 48774 21836 48780 21888
rect 48832 21876 48838 21888
rect 57882 21876 57888 21888
rect 48832 21848 57888 21876
rect 48832 21836 48838 21848
rect 57882 21836 57888 21848
rect 57940 21836 57946 21888
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 13354 21632 13360 21684
rect 13412 21672 13418 21684
rect 14185 21675 14243 21681
rect 14185 21672 14197 21675
rect 13412 21644 14197 21672
rect 13412 21632 13418 21644
rect 14185 21641 14197 21644
rect 14231 21672 14243 21675
rect 15562 21672 15568 21684
rect 14231 21644 15568 21672
rect 14231 21641 14243 21644
rect 14185 21635 14243 21641
rect 15562 21632 15568 21644
rect 15620 21632 15626 21684
rect 20349 21675 20407 21681
rect 20349 21672 20361 21675
rect 16132 21644 20361 21672
rect 7650 21564 7656 21616
rect 7708 21604 7714 21616
rect 13722 21604 13728 21616
rect 7708 21576 13728 21604
rect 7708 21564 7714 21576
rect 13722 21564 13728 21576
rect 13780 21564 13786 21616
rect 15930 21604 15936 21616
rect 13832 21576 15936 21604
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 13832 21536 13860 21576
rect 15930 21564 15936 21576
rect 15988 21564 15994 21616
rect 1719 21508 13860 21536
rect 13909 21539 13967 21545
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 13909 21505 13921 21539
rect 13955 21536 13967 21539
rect 15194 21536 15200 21548
rect 13955 21508 15200 21536
rect 13955 21505 13967 21508
rect 13909 21499 13967 21505
rect 15194 21496 15200 21508
rect 15252 21496 15258 21548
rect 15473 21539 15531 21545
rect 15473 21505 15485 21539
rect 15519 21505 15531 21539
rect 15654 21536 15660 21548
rect 15615 21508 15660 21536
rect 15473 21499 15531 21505
rect 1854 21468 1860 21480
rect 1815 21440 1860 21468
rect 1854 21428 1860 21440
rect 1912 21428 1918 21480
rect 15488 21468 15516 21499
rect 15654 21496 15660 21508
rect 15712 21496 15718 21548
rect 16132 21545 16160 21644
rect 20349 21641 20361 21644
rect 20395 21641 20407 21675
rect 20349 21635 20407 21641
rect 20438 21632 20444 21684
rect 20496 21672 20502 21684
rect 21174 21672 21180 21684
rect 20496 21644 21180 21672
rect 20496 21632 20502 21644
rect 21174 21632 21180 21644
rect 21232 21672 21238 21684
rect 25501 21675 25559 21681
rect 25501 21672 25513 21675
rect 21232 21644 25513 21672
rect 21232 21632 21238 21644
rect 25501 21641 25513 21644
rect 25547 21641 25559 21675
rect 27154 21672 27160 21684
rect 27115 21644 27160 21672
rect 25501 21635 25559 21641
rect 27154 21632 27160 21644
rect 27212 21632 27218 21684
rect 27341 21675 27399 21681
rect 27341 21641 27353 21675
rect 27387 21672 27399 21675
rect 27430 21672 27436 21684
rect 27387 21644 27436 21672
rect 27387 21641 27399 21644
rect 27341 21635 27399 21641
rect 27430 21632 27436 21644
rect 27488 21632 27494 21684
rect 30650 21632 30656 21684
rect 30708 21672 30714 21684
rect 31757 21675 31815 21681
rect 31757 21672 31769 21675
rect 30708 21644 31769 21672
rect 30708 21632 30714 21644
rect 31757 21641 31769 21644
rect 31803 21641 31815 21675
rect 31757 21635 31815 21641
rect 34606 21632 34612 21684
rect 34664 21672 34670 21684
rect 35434 21672 35440 21684
rect 34664 21644 35342 21672
rect 35395 21644 35440 21672
rect 34664 21632 34670 21644
rect 16206 21564 16212 21616
rect 16264 21604 16270 21616
rect 19426 21604 19432 21616
rect 16264 21576 19432 21604
rect 16264 21564 16270 21576
rect 17236 21545 17264 21576
rect 19426 21564 19432 21576
rect 19484 21564 19490 21616
rect 22640 21607 22698 21613
rect 22640 21573 22652 21607
rect 22686 21604 22698 21607
rect 22922 21604 22928 21616
rect 22686 21576 22928 21604
rect 22686 21573 22698 21576
rect 22640 21567 22698 21573
rect 22922 21564 22928 21576
rect 22980 21564 22986 21616
rect 29730 21604 29736 21616
rect 24320 21576 29736 21604
rect 24320 21548 24348 21576
rect 29730 21564 29736 21576
rect 29788 21564 29794 21616
rect 29822 21564 29828 21616
rect 29880 21604 29886 21616
rect 32554 21607 32612 21613
rect 32554 21604 32566 21607
rect 29880 21576 32566 21604
rect 29880 21564 29886 21576
rect 32554 21573 32566 21576
rect 32600 21573 32612 21607
rect 32554 21567 32612 21573
rect 33410 21564 33416 21616
rect 33468 21604 33474 21616
rect 34793 21607 34851 21613
rect 34793 21604 34805 21607
rect 33468 21576 34805 21604
rect 33468 21564 33474 21576
rect 34793 21573 34805 21576
rect 34839 21573 34851 21607
rect 35314 21604 35342 21644
rect 35434 21632 35440 21644
rect 35492 21632 35498 21684
rect 35710 21632 35716 21684
rect 35768 21672 35774 21684
rect 35768 21644 35940 21672
rect 35768 21632 35774 21644
rect 35314 21576 35848 21604
rect 34793 21567 34851 21573
rect 35452 21548 35480 21576
rect 16117 21539 16175 21545
rect 16117 21505 16129 21539
rect 16163 21505 16175 21539
rect 16117 21499 16175 21505
rect 16301 21539 16359 21545
rect 16301 21505 16313 21539
rect 16347 21505 16359 21539
rect 16301 21499 16359 21505
rect 17221 21539 17279 21545
rect 17221 21505 17233 21539
rect 17267 21505 17279 21539
rect 17221 21499 17279 21505
rect 17488 21539 17546 21545
rect 17488 21505 17500 21539
rect 17534 21536 17546 21539
rect 17954 21536 17960 21548
rect 17534 21508 17960 21536
rect 17534 21505 17546 21508
rect 17488 21499 17546 21505
rect 16022 21468 16028 21480
rect 15488 21440 16028 21468
rect 16022 21428 16028 21440
rect 16080 21468 16086 21480
rect 16316 21468 16344 21499
rect 17954 21496 17960 21508
rect 18012 21496 18018 21548
rect 19150 21536 19156 21548
rect 19111 21508 19156 21536
rect 19150 21496 19156 21508
rect 19208 21496 19214 21548
rect 22370 21536 22376 21548
rect 22331 21508 22376 21536
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 24302 21496 24308 21548
rect 24360 21536 24366 21548
rect 27338 21536 27344 21548
rect 24360 21508 24405 21536
rect 27299 21508 27344 21536
rect 24360 21496 24366 21508
rect 27338 21496 27344 21508
rect 27396 21496 27402 21548
rect 27614 21496 27620 21548
rect 27672 21536 27678 21548
rect 27801 21539 27859 21545
rect 27801 21536 27813 21539
rect 27672 21508 27813 21536
rect 27672 21496 27678 21508
rect 27801 21505 27813 21508
rect 27847 21505 27859 21539
rect 27801 21499 27859 21505
rect 28629 21539 28687 21545
rect 28629 21505 28641 21539
rect 28675 21536 28687 21539
rect 30190 21536 30196 21548
rect 28675 21508 30196 21536
rect 28675 21505 28687 21508
rect 28629 21499 28687 21505
rect 30190 21496 30196 21508
rect 30248 21496 30254 21548
rect 31386 21536 31392 21548
rect 31347 21508 31392 21536
rect 31386 21496 31392 21508
rect 31444 21496 31450 21548
rect 31570 21536 31576 21548
rect 31531 21508 31576 21536
rect 31570 21496 31576 21508
rect 31628 21536 31634 21548
rect 34330 21536 34336 21548
rect 31628 21508 33732 21536
rect 31628 21496 31634 21508
rect 16080 21440 16344 21468
rect 16080 21428 16086 21440
rect 24394 21428 24400 21480
rect 24452 21468 24458 21480
rect 26142 21468 26148 21480
rect 24452 21440 26148 21468
rect 24452 21428 24458 21440
rect 26142 21428 26148 21440
rect 26200 21428 26206 21480
rect 26252 21440 27384 21468
rect 15565 21403 15623 21409
rect 15565 21369 15577 21403
rect 15611 21400 15623 21403
rect 16942 21400 16948 21412
rect 15611 21372 16948 21400
rect 15611 21369 15623 21372
rect 15565 21363 15623 21369
rect 16942 21360 16948 21372
rect 17000 21360 17006 21412
rect 19150 21400 19156 21412
rect 18432 21372 19156 21400
rect 16117 21335 16175 21341
rect 16117 21301 16129 21335
rect 16163 21332 16175 21335
rect 18432 21332 18460 21372
rect 19150 21360 19156 21372
rect 19208 21360 19214 21412
rect 19334 21360 19340 21412
rect 19392 21400 19398 21412
rect 26252 21400 26280 21440
rect 19392 21372 21404 21400
rect 19392 21360 19398 21372
rect 18598 21332 18604 21344
rect 16163 21304 18460 21332
rect 18559 21304 18604 21332
rect 16163 21301 16175 21304
rect 16117 21295 16175 21301
rect 18598 21292 18604 21304
rect 18656 21292 18662 21344
rect 20898 21292 20904 21344
rect 20956 21332 20962 21344
rect 21266 21332 21272 21344
rect 20956 21304 21272 21332
rect 20956 21292 20962 21304
rect 21266 21292 21272 21304
rect 21324 21292 21330 21344
rect 21376 21332 21404 21372
rect 23308 21372 26280 21400
rect 27356 21400 27384 21440
rect 28902 21428 28908 21480
rect 28960 21468 28966 21480
rect 32309 21471 32367 21477
rect 32309 21468 32321 21471
rect 28960 21440 32321 21468
rect 28960 21428 28966 21440
rect 32309 21437 32321 21440
rect 32355 21437 32367 21471
rect 32309 21431 32367 21437
rect 30374 21400 30380 21412
rect 27356 21372 30380 21400
rect 23308 21332 23336 21372
rect 30374 21360 30380 21372
rect 30432 21360 30438 21412
rect 31294 21360 31300 21412
rect 31352 21400 31358 21412
rect 31570 21400 31576 21412
rect 31352 21372 31576 21400
rect 31352 21360 31358 21372
rect 31570 21360 31576 21372
rect 31628 21360 31634 21412
rect 33704 21409 33732 21508
rect 33796 21508 34336 21536
rect 33689 21403 33747 21409
rect 33689 21369 33701 21403
rect 33735 21369 33747 21403
rect 33689 21363 33747 21369
rect 21376 21304 23336 21332
rect 23753 21335 23811 21341
rect 23753 21301 23765 21335
rect 23799 21332 23811 21335
rect 26694 21332 26700 21344
rect 23799 21304 26700 21332
rect 23799 21301 23811 21304
rect 23753 21295 23811 21301
rect 26694 21292 26700 21304
rect 26752 21292 26758 21344
rect 27706 21332 27712 21344
rect 27667 21304 27712 21332
rect 27706 21292 27712 21304
rect 27764 21292 27770 21344
rect 27798 21292 27804 21344
rect 27856 21332 27862 21344
rect 29825 21335 29883 21341
rect 29825 21332 29837 21335
rect 27856 21304 29837 21332
rect 27856 21292 27862 21304
rect 29825 21301 29837 21304
rect 29871 21301 29883 21335
rect 30392 21332 30420 21360
rect 33796 21332 33824 21508
rect 34330 21496 34336 21508
rect 34388 21536 34394 21548
rect 34609 21539 34667 21545
rect 34609 21536 34621 21539
rect 34388 21508 34621 21536
rect 34388 21496 34394 21508
rect 34609 21505 34621 21508
rect 34655 21505 34667 21539
rect 34609 21499 34667 21505
rect 35434 21496 35440 21548
rect 35492 21496 35498 21548
rect 35710 21536 35716 21548
rect 35671 21508 35716 21536
rect 35710 21496 35716 21508
rect 35768 21496 35774 21548
rect 35820 21545 35848 21576
rect 35912 21545 35940 21644
rect 36446 21632 36452 21684
rect 36504 21672 36510 21684
rect 36504 21644 46244 21672
rect 36504 21632 36510 21644
rect 36998 21564 37004 21616
rect 37056 21604 37062 21616
rect 37056 21576 38056 21604
rect 37056 21564 37062 21576
rect 35805 21539 35863 21545
rect 35805 21505 35817 21539
rect 35851 21505 35863 21539
rect 35805 21499 35863 21505
rect 35897 21539 35955 21545
rect 35897 21505 35909 21539
rect 35943 21505 35955 21539
rect 35897 21499 35955 21505
rect 36078 21496 36084 21548
rect 36136 21536 36142 21548
rect 36136 21508 36229 21536
rect 36136 21496 36142 21508
rect 36262 21496 36268 21548
rect 36320 21536 36326 21548
rect 36541 21539 36599 21545
rect 36541 21536 36553 21539
rect 36320 21508 36553 21536
rect 36320 21496 36326 21508
rect 36541 21505 36553 21508
rect 36587 21505 36599 21539
rect 36541 21499 36599 21505
rect 36725 21539 36783 21545
rect 36725 21505 36737 21539
rect 36771 21536 36783 21539
rect 37366 21536 37372 21548
rect 36771 21508 37372 21536
rect 36771 21505 36783 21508
rect 36725 21499 36783 21505
rect 37366 21496 37372 21508
rect 37424 21536 37430 21548
rect 37829 21539 37887 21545
rect 37829 21536 37841 21539
rect 37424 21508 37841 21536
rect 37424 21496 37430 21508
rect 37829 21505 37841 21508
rect 37875 21505 37887 21539
rect 37829 21499 37887 21505
rect 33962 21428 33968 21480
rect 34020 21468 34026 21480
rect 34885 21471 34943 21477
rect 34885 21468 34897 21471
rect 34020 21440 34897 21468
rect 34020 21428 34026 21440
rect 34885 21437 34897 21440
rect 34931 21437 34943 21471
rect 36096 21468 36124 21496
rect 36906 21468 36912 21480
rect 36096 21440 36912 21468
rect 34885 21431 34943 21437
rect 36906 21428 36912 21440
rect 36964 21428 36970 21480
rect 37642 21428 37648 21480
rect 37700 21468 37706 21480
rect 38028 21477 38056 21576
rect 38838 21564 38844 21616
rect 38896 21604 38902 21616
rect 46216 21604 46244 21644
rect 47854 21632 47860 21684
rect 47912 21672 47918 21684
rect 51626 21672 51632 21684
rect 47912 21644 51632 21672
rect 47912 21632 47918 21644
rect 51626 21632 51632 21644
rect 51684 21632 51690 21684
rect 58802 21604 58808 21616
rect 38896 21576 45554 21604
rect 46216 21576 58808 21604
rect 38896 21564 38902 21576
rect 40402 21536 40408 21548
rect 40363 21508 40408 21536
rect 40402 21496 40408 21508
rect 40460 21496 40466 21548
rect 40494 21496 40500 21548
rect 40552 21536 40558 21548
rect 44266 21545 44272 21548
rect 40661 21539 40719 21545
rect 40661 21536 40673 21539
rect 40552 21508 40673 21536
rect 40552 21496 40558 21508
rect 40661 21505 40673 21508
rect 40707 21505 40719 21539
rect 40661 21499 40719 21505
rect 44260 21499 44272 21545
rect 44324 21536 44330 21548
rect 45526 21536 45554 21576
rect 58802 21564 58808 21576
rect 58860 21564 58866 21616
rect 48498 21536 48504 21548
rect 44324 21508 44360 21536
rect 45526 21508 48504 21536
rect 44266 21496 44272 21499
rect 44324 21496 44330 21508
rect 48498 21496 48504 21508
rect 48556 21536 48562 21548
rect 48556 21508 50108 21536
rect 48556 21496 48562 21508
rect 37921 21471 37979 21477
rect 37921 21468 37933 21471
rect 37700 21440 37933 21468
rect 37700 21428 37706 21440
rect 37921 21437 37933 21440
rect 37967 21437 37979 21471
rect 37921 21431 37979 21437
rect 38013 21471 38071 21477
rect 38013 21437 38025 21471
rect 38059 21437 38071 21471
rect 38013 21431 38071 21437
rect 37936 21400 37964 21431
rect 43346 21428 43352 21480
rect 43404 21468 43410 21480
rect 50080 21477 50108 21508
rect 50154 21496 50160 21548
rect 50212 21536 50218 21548
rect 50249 21539 50307 21545
rect 50249 21536 50261 21539
rect 50212 21508 50261 21536
rect 50212 21496 50218 21508
rect 50249 21505 50261 21508
rect 50295 21505 50307 21539
rect 50249 21499 50307 21505
rect 56226 21496 56232 21548
rect 56284 21536 56290 21548
rect 56413 21539 56471 21545
rect 56413 21536 56425 21539
rect 56284 21508 56425 21536
rect 56284 21496 56290 21508
rect 56413 21505 56425 21508
rect 56459 21505 56471 21539
rect 56413 21499 56471 21505
rect 56597 21539 56655 21545
rect 56597 21505 56609 21539
rect 56643 21536 56655 21539
rect 56778 21536 56784 21548
rect 56643 21508 56784 21536
rect 56643 21505 56655 21508
rect 56597 21499 56655 21505
rect 56778 21496 56784 21508
rect 56836 21496 56842 21548
rect 57146 21536 57152 21548
rect 57107 21508 57152 21536
rect 57146 21496 57152 21508
rect 57204 21496 57210 21548
rect 43993 21471 44051 21477
rect 43993 21468 44005 21471
rect 43404 21440 44005 21468
rect 43404 21428 43410 21440
rect 43993 21437 44005 21440
rect 44039 21437 44051 21471
rect 43993 21431 44051 21437
rect 50065 21471 50123 21477
rect 50065 21437 50077 21471
rect 50111 21468 50123 21471
rect 51994 21468 52000 21480
rect 50111 21440 52000 21468
rect 50111 21437 50123 21440
rect 50065 21431 50123 21437
rect 51994 21428 52000 21440
rect 52052 21428 52058 21480
rect 38286 21400 38292 21412
rect 35820 21372 37596 21400
rect 37936 21372 38292 21400
rect 30392 21304 33824 21332
rect 34333 21335 34391 21341
rect 29825 21295 29883 21301
rect 34333 21301 34345 21335
rect 34379 21332 34391 21335
rect 35820 21332 35848 21372
rect 34379 21304 35848 21332
rect 36909 21335 36967 21341
rect 34379 21301 34391 21304
rect 34333 21295 34391 21301
rect 36909 21301 36921 21335
rect 36955 21332 36967 21335
rect 36998 21332 37004 21344
rect 36955 21304 37004 21332
rect 36955 21301 36967 21304
rect 36909 21295 36967 21301
rect 36998 21292 37004 21304
rect 37056 21292 37062 21344
rect 37458 21332 37464 21344
rect 37419 21304 37464 21332
rect 37458 21292 37464 21304
rect 37516 21292 37522 21344
rect 37568 21332 37596 21372
rect 38286 21360 38292 21372
rect 38344 21360 38350 21412
rect 55950 21400 55956 21412
rect 41386 21372 41920 21400
rect 41386 21332 41414 21372
rect 41782 21332 41788 21344
rect 37568 21304 41414 21332
rect 41743 21304 41788 21332
rect 41782 21292 41788 21304
rect 41840 21292 41846 21344
rect 41892 21332 41920 21372
rect 45296 21372 55956 21400
rect 45296 21332 45324 21372
rect 55950 21360 55956 21372
rect 56008 21360 56014 21412
rect 41892 21304 45324 21332
rect 45370 21292 45376 21344
rect 45428 21332 45434 21344
rect 48774 21332 48780 21344
rect 45428 21304 48780 21332
rect 45428 21292 45434 21304
rect 48774 21292 48780 21304
rect 48832 21292 48838 21344
rect 50430 21332 50436 21344
rect 50391 21304 50436 21332
rect 50430 21292 50436 21304
rect 50488 21292 50494 21344
rect 56413 21335 56471 21341
rect 56413 21301 56425 21335
rect 56459 21332 56471 21335
rect 56962 21332 56968 21344
rect 56459 21304 56968 21332
rect 56459 21301 56471 21304
rect 56413 21295 56471 21301
rect 56962 21292 56968 21304
rect 57020 21292 57026 21344
rect 57238 21332 57244 21344
rect 57199 21304 57244 21332
rect 57238 21292 57244 21304
rect 57296 21292 57302 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 17770 21128 17776 21140
rect 17731 21100 17776 21128
rect 17770 21088 17776 21100
rect 17828 21088 17834 21140
rect 18598 21088 18604 21140
rect 18656 21128 18662 21140
rect 29362 21128 29368 21140
rect 18656 21100 29368 21128
rect 18656 21088 18662 21100
rect 29362 21088 29368 21100
rect 29420 21088 29426 21140
rect 29454 21088 29460 21140
rect 29512 21128 29518 21140
rect 29825 21131 29883 21137
rect 29825 21128 29837 21131
rect 29512 21100 29837 21128
rect 29512 21088 29518 21100
rect 29825 21097 29837 21100
rect 29871 21097 29883 21131
rect 29825 21091 29883 21097
rect 29914 21088 29920 21140
rect 29972 21128 29978 21140
rect 31018 21128 31024 21140
rect 29972 21100 31024 21128
rect 29972 21088 29978 21100
rect 31018 21088 31024 21100
rect 31076 21128 31082 21140
rect 31294 21128 31300 21140
rect 31076 21100 31300 21128
rect 31076 21088 31082 21100
rect 31294 21088 31300 21100
rect 31352 21088 31358 21140
rect 31386 21088 31392 21140
rect 31444 21128 31450 21140
rect 31754 21128 31760 21140
rect 31444 21100 31760 21128
rect 31444 21088 31450 21100
rect 31754 21088 31760 21100
rect 31812 21128 31818 21140
rect 36262 21128 36268 21140
rect 31812 21100 36268 21128
rect 31812 21088 31818 21100
rect 36262 21088 36268 21100
rect 36320 21088 36326 21140
rect 36354 21088 36360 21140
rect 36412 21128 36418 21140
rect 40957 21131 41015 21137
rect 40957 21128 40969 21131
rect 36412 21100 40969 21128
rect 36412 21088 36418 21100
rect 40957 21097 40969 21100
rect 41003 21097 41015 21131
rect 40957 21091 41015 21097
rect 44450 21088 44456 21140
rect 44508 21128 44514 21140
rect 48133 21131 48191 21137
rect 48133 21128 48145 21131
rect 44508 21100 48145 21128
rect 44508 21088 44514 21100
rect 48133 21097 48145 21100
rect 48179 21097 48191 21131
rect 51718 21128 51724 21140
rect 51679 21100 51724 21128
rect 48133 21091 48191 21097
rect 51718 21088 51724 21100
rect 51776 21088 51782 21140
rect 57790 21088 57796 21140
rect 57848 21128 57854 21140
rect 58253 21131 58311 21137
rect 58253 21128 58265 21131
rect 57848 21100 58265 21128
rect 57848 21088 57854 21100
rect 58253 21097 58265 21100
rect 58299 21097 58311 21131
rect 58253 21091 58311 21097
rect 16025 21063 16083 21069
rect 16025 21029 16037 21063
rect 16071 21060 16083 21063
rect 19334 21060 19340 21072
rect 16071 21032 19340 21060
rect 16071 21029 16083 21032
rect 16025 21023 16083 21029
rect 19334 21020 19340 21032
rect 19392 21020 19398 21072
rect 20809 21063 20867 21069
rect 20809 21029 20821 21063
rect 20855 21060 20867 21063
rect 24302 21060 24308 21072
rect 20855 21032 24308 21060
rect 20855 21029 20867 21032
rect 20809 21023 20867 21029
rect 24302 21020 24308 21032
rect 24360 21020 24366 21072
rect 26789 21063 26847 21069
rect 26789 21060 26801 21063
rect 24412 21032 26801 21060
rect 14461 20995 14519 21001
rect 14461 20961 14473 20995
rect 14507 20992 14519 20995
rect 15930 20992 15936 21004
rect 14507 20964 15936 20992
rect 14507 20961 14519 20964
rect 14461 20955 14519 20961
rect 15930 20952 15936 20964
rect 15988 20952 15994 21004
rect 24412 20992 24440 21032
rect 26789 21029 26801 21032
rect 26835 21029 26847 21063
rect 26789 21023 26847 21029
rect 27246 21020 27252 21072
rect 27304 21060 27310 21072
rect 27798 21060 27804 21072
rect 27304 21032 27804 21060
rect 27304 21020 27310 21032
rect 27798 21020 27804 21032
rect 27856 21020 27862 21072
rect 28353 21063 28411 21069
rect 28353 21029 28365 21063
rect 28399 21060 28411 21063
rect 35802 21060 35808 21072
rect 28399 21032 35808 21060
rect 28399 21029 28411 21032
rect 28353 21023 28411 21029
rect 35802 21020 35808 21032
rect 35860 21020 35866 21072
rect 37458 21020 37464 21072
rect 37516 21060 37522 21072
rect 47486 21060 47492 21072
rect 37516 21032 47492 21060
rect 37516 21020 37522 21032
rect 47486 21020 47492 21032
rect 47544 21020 47550 21072
rect 20456 20964 24440 20992
rect 24673 20995 24731 21001
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20924 1639 20927
rect 10778 20924 10784 20936
rect 1627 20896 10784 20924
rect 1627 20893 1639 20896
rect 1581 20887 1639 20893
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 14737 20927 14795 20933
rect 14737 20893 14749 20927
rect 14783 20924 14795 20927
rect 15194 20924 15200 20936
rect 14783 20896 15200 20924
rect 14783 20893 14795 20896
rect 14737 20887 14795 20893
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 16574 20924 16580 20936
rect 16535 20896 16580 20924
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 19426 20924 19432 20936
rect 19387 20896 19432 20924
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 20456 20924 20484 20964
rect 24673 20961 24685 20995
rect 24719 20961 24731 20995
rect 31481 20995 31539 21001
rect 31481 20992 31493 20995
rect 24673 20955 24731 20961
rect 25608 20964 31493 20992
rect 21726 20924 21732 20936
rect 19536 20896 20484 20924
rect 21687 20896 21732 20924
rect 1854 20856 1860 20868
rect 1815 20828 1860 20856
rect 1854 20816 1860 20828
rect 1912 20816 1918 20868
rect 18138 20856 18144 20868
rect 16960 20828 18144 20856
rect 13722 20748 13728 20800
rect 13780 20788 13786 20800
rect 16960 20788 16988 20828
rect 18138 20816 18144 20828
rect 18196 20816 18202 20868
rect 18414 20816 18420 20868
rect 18472 20856 18478 20868
rect 19536 20856 19564 20896
rect 21726 20884 21732 20896
rect 21784 20884 21790 20936
rect 22646 20884 22652 20936
rect 22704 20924 22710 20936
rect 24688 20924 24716 20955
rect 22704 20896 24716 20924
rect 24765 20927 24823 20933
rect 22704 20884 22710 20896
rect 24765 20893 24777 20927
rect 24811 20924 24823 20927
rect 24854 20924 24860 20936
rect 24811 20896 24860 20924
rect 24811 20893 24823 20896
rect 24765 20887 24823 20893
rect 24854 20884 24860 20896
rect 24912 20884 24918 20936
rect 25608 20933 25636 20964
rect 31481 20961 31493 20964
rect 31527 20961 31539 20995
rect 31481 20955 31539 20961
rect 32306 20952 32312 21004
rect 32364 20992 32370 21004
rect 33873 20995 33931 21001
rect 33873 20992 33885 20995
rect 32364 20964 33885 20992
rect 32364 20952 32370 20964
rect 33873 20961 33885 20964
rect 33919 20961 33931 20995
rect 33873 20955 33931 20961
rect 35434 20952 35440 21004
rect 35492 20992 35498 21004
rect 36078 20992 36084 21004
rect 35492 20964 36084 20992
rect 35492 20952 35498 20964
rect 36078 20952 36084 20964
rect 36136 20992 36142 21004
rect 40218 20992 40224 21004
rect 36136 20964 36676 20992
rect 36136 20952 36142 20964
rect 25593 20927 25651 20933
rect 25593 20893 25605 20927
rect 25639 20893 25651 20927
rect 25593 20887 25651 20893
rect 26142 20884 26148 20936
rect 26200 20924 26206 20936
rect 28350 20924 28356 20936
rect 26200 20896 28356 20924
rect 26200 20884 26206 20896
rect 28350 20884 28356 20896
rect 28408 20884 28414 20936
rect 28534 20924 28540 20936
rect 28495 20896 28540 20924
rect 28534 20884 28540 20896
rect 28592 20884 28598 20936
rect 28810 20924 28816 20936
rect 28771 20896 28816 20924
rect 28810 20884 28816 20896
rect 28868 20884 28874 20936
rect 29733 20927 29791 20933
rect 29733 20893 29745 20927
rect 29779 20893 29791 20927
rect 30374 20924 30380 20936
rect 30335 20896 30380 20924
rect 29733 20887 29791 20893
rect 18472 20828 19564 20856
rect 19696 20859 19754 20865
rect 18472 20816 18478 20828
rect 19696 20825 19708 20859
rect 19742 20856 19754 20859
rect 20990 20856 20996 20868
rect 19742 20828 20996 20856
rect 19742 20825 19754 20828
rect 19696 20819 19754 20825
rect 20990 20816 20996 20828
rect 21048 20816 21054 20868
rect 28721 20859 28779 20865
rect 28721 20856 28733 20859
rect 22066 20828 28733 20856
rect 13780 20760 16988 20788
rect 13780 20748 13786 20760
rect 17034 20748 17040 20800
rect 17092 20788 17098 20800
rect 22066 20788 22094 20828
rect 28721 20825 28733 20828
rect 28767 20825 28779 20859
rect 29748 20856 29776 20887
rect 30374 20884 30380 20896
rect 30432 20884 30438 20936
rect 35069 20927 35127 20933
rect 35069 20893 35081 20927
rect 35115 20924 35127 20927
rect 35342 20924 35348 20936
rect 35115 20896 35348 20924
rect 35115 20893 35127 20896
rect 35069 20887 35127 20893
rect 35342 20884 35348 20896
rect 35400 20884 35406 20936
rect 36262 20884 36268 20936
rect 36320 20884 36326 20936
rect 36446 20884 36452 20936
rect 36504 20933 36510 20936
rect 36648 20933 36676 20964
rect 37384 20964 40224 20992
rect 36504 20927 36553 20933
rect 36504 20893 36507 20927
rect 36541 20893 36553 20927
rect 36504 20887 36553 20893
rect 36633 20927 36691 20933
rect 36633 20893 36645 20927
rect 36679 20893 36691 20927
rect 36633 20887 36691 20893
rect 36746 20924 36804 20930
rect 36746 20890 36758 20924
rect 36792 20890 36829 20924
rect 36504 20884 36510 20887
rect 36746 20884 36829 20890
rect 36906 20884 36912 20936
rect 36964 20924 36970 20936
rect 36964 20896 37009 20924
rect 36964 20884 36970 20896
rect 30466 20856 30472 20868
rect 29748 20828 30472 20856
rect 28721 20819 28779 20825
rect 30466 20816 30472 20828
rect 30524 20816 30530 20868
rect 33137 20859 33195 20865
rect 33137 20856 33149 20859
rect 32600 20828 33149 20856
rect 22922 20788 22928 20800
rect 17092 20760 22094 20788
rect 22883 20760 22928 20788
rect 17092 20748 17098 20760
rect 22922 20748 22928 20760
rect 22980 20748 22986 20800
rect 25133 20791 25191 20797
rect 25133 20757 25145 20791
rect 25179 20788 25191 20791
rect 25314 20788 25320 20800
rect 25179 20760 25320 20788
rect 25179 20757 25191 20760
rect 25133 20751 25191 20757
rect 25314 20748 25320 20760
rect 25372 20748 25378 20800
rect 26694 20748 26700 20800
rect 26752 20788 26758 20800
rect 27338 20788 27344 20800
rect 26752 20760 27344 20788
rect 26752 20748 26758 20760
rect 27338 20748 27344 20760
rect 27396 20748 27402 20800
rect 27706 20748 27712 20800
rect 27764 20788 27770 20800
rect 28442 20788 28448 20800
rect 27764 20760 28448 20788
rect 27764 20748 27770 20760
rect 28442 20748 28448 20760
rect 28500 20788 28506 20800
rect 32600 20788 32628 20828
rect 33137 20825 33149 20828
rect 33183 20856 33195 20859
rect 33962 20856 33968 20868
rect 33183 20828 33968 20856
rect 33183 20825 33195 20828
rect 33137 20819 33195 20825
rect 33962 20816 33968 20828
rect 34020 20816 34026 20868
rect 34885 20859 34943 20865
rect 34885 20825 34897 20859
rect 34931 20825 34943 20859
rect 35434 20856 35440 20868
rect 35395 20828 35440 20856
rect 34885 20819 34943 20825
rect 28500 20760 32628 20788
rect 28500 20748 28506 20760
rect 32674 20748 32680 20800
rect 32732 20788 32738 20800
rect 34900 20788 34928 20819
rect 35434 20816 35440 20828
rect 35492 20856 35498 20868
rect 35618 20856 35624 20868
rect 35492 20828 35624 20856
rect 35492 20816 35498 20828
rect 35618 20816 35624 20828
rect 35676 20816 35682 20868
rect 36280 20856 36308 20884
rect 36801 20856 36829 20884
rect 36998 20856 37004 20868
rect 36280 20828 36676 20856
rect 36801 20828 37004 20856
rect 36262 20788 36268 20800
rect 32732 20760 34928 20788
rect 36223 20760 36268 20788
rect 32732 20748 32738 20760
rect 36262 20748 36268 20760
rect 36320 20748 36326 20800
rect 36648 20788 36676 20828
rect 36998 20816 37004 20828
rect 37056 20816 37062 20868
rect 37384 20865 37412 20964
rect 40218 20952 40224 20964
rect 40276 20952 40282 21004
rect 41782 20992 41788 21004
rect 40880 20964 41788 20992
rect 38194 20924 38200 20936
rect 38155 20896 38200 20924
rect 38194 20884 38200 20896
rect 38252 20884 38258 20936
rect 40586 20927 40644 20933
rect 40586 20893 40598 20927
rect 40632 20924 40644 20927
rect 40880 20924 40908 20964
rect 41782 20952 41788 20964
rect 41840 20952 41846 21004
rect 43346 20992 43352 21004
rect 43307 20964 43352 20992
rect 43346 20952 43352 20964
rect 43404 20952 43410 21004
rect 43438 20952 43444 21004
rect 43496 20992 43502 21004
rect 44634 20992 44640 21004
rect 43496 20964 44640 20992
rect 43496 20952 43502 20964
rect 44634 20952 44640 20964
rect 44692 20992 44698 21004
rect 48222 20992 48228 21004
rect 44692 20964 48228 20992
rect 44692 20952 44698 20964
rect 48222 20952 48228 20964
rect 48280 20952 48286 21004
rect 56226 20992 56232 21004
rect 56187 20964 56232 20992
rect 56226 20952 56232 20964
rect 56284 20952 56290 21004
rect 56870 20992 56876 21004
rect 56831 20964 56876 20992
rect 56870 20952 56876 20964
rect 56928 20952 56934 21004
rect 40632 20896 40908 20924
rect 41061 20927 41119 20933
rect 40632 20893 40644 20896
rect 40586 20887 40644 20893
rect 41061 20893 41073 20927
rect 41107 20924 41119 20927
rect 41322 20924 41328 20936
rect 41107 20896 41328 20924
rect 41107 20893 41119 20896
rect 41061 20887 41119 20893
rect 41322 20884 41328 20896
rect 41380 20924 41386 20936
rect 42794 20924 42800 20936
rect 41380 20896 42800 20924
rect 41380 20884 41386 20896
rect 42794 20884 42800 20896
rect 42852 20884 42858 20936
rect 48130 20884 48136 20936
rect 48188 20924 48194 20936
rect 50341 20927 50399 20933
rect 50341 20924 50353 20927
rect 48188 20896 50353 20924
rect 48188 20884 48194 20896
rect 50341 20893 50353 20896
rect 50387 20924 50399 20927
rect 52362 20924 52368 20936
rect 50387 20896 52368 20924
rect 50387 20893 50399 20896
rect 50341 20887 50399 20893
rect 52362 20884 52368 20896
rect 52420 20884 52426 20936
rect 56042 20884 56048 20936
rect 56100 20924 56106 20936
rect 56326 20927 56384 20933
rect 56326 20924 56338 20927
rect 56100 20896 56338 20924
rect 56100 20884 56106 20896
rect 56326 20893 56338 20896
rect 56372 20893 56384 20927
rect 56326 20887 56384 20893
rect 37369 20859 37427 20865
rect 37369 20825 37381 20859
rect 37415 20825 37427 20859
rect 37550 20856 37556 20868
rect 37511 20828 37556 20856
rect 37369 20819 37427 20825
rect 37384 20788 37412 20819
rect 37550 20816 37556 20828
rect 37608 20816 37614 20868
rect 37642 20816 37648 20868
rect 37700 20856 37706 20868
rect 40678 20856 40684 20868
rect 37700 20828 40684 20856
rect 37700 20816 37706 20828
rect 40678 20816 40684 20828
rect 40736 20816 40742 20868
rect 41601 20859 41659 20865
rect 41601 20825 41613 20859
rect 41647 20856 41659 20859
rect 46842 20856 46848 20868
rect 41647 20828 46848 20856
rect 41647 20825 41659 20828
rect 41601 20819 41659 20825
rect 46842 20816 46848 20828
rect 46900 20816 46906 20868
rect 50430 20816 50436 20868
rect 50488 20856 50494 20868
rect 50586 20859 50644 20865
rect 50586 20856 50598 20859
rect 50488 20828 50598 20856
rect 50488 20816 50494 20828
rect 50586 20825 50598 20828
rect 50632 20825 50644 20859
rect 55953 20859 56011 20865
rect 55953 20856 55965 20859
rect 50586 20819 50644 20825
rect 51046 20828 55965 20856
rect 36648 20760 37412 20788
rect 37737 20791 37795 20797
rect 37737 20757 37749 20791
rect 37783 20788 37795 20791
rect 37918 20788 37924 20800
rect 37783 20760 37924 20788
rect 37783 20757 37795 20760
rect 37737 20751 37795 20757
rect 37918 20748 37924 20760
rect 37976 20748 37982 20800
rect 38378 20788 38384 20800
rect 38339 20760 38384 20788
rect 38378 20748 38384 20760
rect 38436 20748 38442 20800
rect 40310 20748 40316 20800
rect 40368 20788 40374 20800
rect 40405 20791 40463 20797
rect 40405 20788 40417 20791
rect 40368 20760 40417 20788
rect 40368 20748 40374 20760
rect 40405 20757 40417 20760
rect 40451 20757 40463 20791
rect 40586 20788 40592 20800
rect 40547 20760 40592 20788
rect 40405 20751 40463 20757
rect 40586 20748 40592 20760
rect 40644 20748 40650 20800
rect 45554 20748 45560 20800
rect 45612 20788 45618 20800
rect 46106 20788 46112 20800
rect 45612 20760 46112 20788
rect 45612 20748 45618 20760
rect 46106 20748 46112 20760
rect 46164 20748 46170 20800
rect 48314 20748 48320 20800
rect 48372 20788 48378 20800
rect 51046 20788 51074 20828
rect 55953 20825 55965 20828
rect 55999 20825 56011 20859
rect 56134 20856 56140 20868
rect 56095 20828 56140 20856
rect 55953 20819 56011 20825
rect 56134 20816 56140 20828
rect 56192 20816 56198 20868
rect 56229 20859 56287 20865
rect 56229 20825 56241 20859
rect 56275 20825 56287 20859
rect 56336 20856 56364 20887
rect 56962 20884 56968 20936
rect 57020 20924 57026 20936
rect 57129 20927 57187 20933
rect 57129 20924 57141 20927
rect 57020 20896 57141 20924
rect 57020 20884 57026 20896
rect 57129 20893 57141 20896
rect 57175 20893 57187 20927
rect 57129 20887 57187 20893
rect 56410 20856 56416 20868
rect 56336 20828 56416 20856
rect 56229 20819 56287 20825
rect 48372 20760 51074 20788
rect 48372 20748 48378 20760
rect 53926 20748 53932 20800
rect 53984 20788 53990 20800
rect 56152 20788 56180 20816
rect 53984 20760 56180 20788
rect 56244 20788 56272 20819
rect 56410 20816 56416 20828
rect 56468 20816 56474 20868
rect 57698 20788 57704 20800
rect 56244 20760 57704 20788
rect 53984 20748 53990 20760
rect 57698 20748 57704 20760
rect 57756 20748 57762 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 16666 20544 16672 20596
rect 16724 20584 16730 20596
rect 17405 20587 17463 20593
rect 17405 20584 17417 20587
rect 16724 20556 17417 20584
rect 16724 20544 16730 20556
rect 17405 20553 17417 20556
rect 17451 20553 17463 20587
rect 23753 20587 23811 20593
rect 17405 20547 17463 20553
rect 18340 20556 19334 20584
rect 15654 20476 15660 20528
rect 15712 20516 15718 20528
rect 18230 20516 18236 20528
rect 15712 20488 18236 20516
rect 15712 20476 15718 20488
rect 1581 20451 1639 20457
rect 1581 20417 1593 20451
rect 1627 20448 1639 20451
rect 15102 20448 15108 20460
rect 1627 20420 15108 20448
rect 1627 20417 1639 20420
rect 1581 20411 1639 20417
rect 15102 20408 15108 20420
rect 15160 20408 15166 20460
rect 15948 20457 15976 20488
rect 18230 20476 18236 20488
rect 18288 20476 18294 20528
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 17037 20451 17095 20457
rect 17037 20417 17049 20451
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 1762 20380 1768 20392
rect 1723 20352 1768 20380
rect 1762 20340 1768 20352
rect 1820 20340 1826 20392
rect 16022 20380 16028 20392
rect 15983 20352 16028 20380
rect 16022 20340 16028 20352
rect 16080 20340 16086 20392
rect 16942 20380 16948 20392
rect 16903 20352 16948 20380
rect 16942 20340 16948 20352
rect 17000 20340 17006 20392
rect 17052 20380 17080 20411
rect 17862 20408 17868 20460
rect 17920 20448 17926 20460
rect 18340 20457 18368 20556
rect 19306 20516 19334 20556
rect 23753 20553 23765 20587
rect 23799 20553 23811 20587
rect 23753 20547 23811 20553
rect 20806 20516 20812 20528
rect 19306 20488 20812 20516
rect 20806 20476 20812 20488
rect 20864 20476 20870 20528
rect 22640 20519 22698 20525
rect 22640 20485 22652 20519
rect 22686 20516 22698 20519
rect 22922 20516 22928 20528
rect 22686 20488 22928 20516
rect 22686 20485 22698 20488
rect 22640 20479 22698 20485
rect 22922 20476 22928 20488
rect 22980 20476 22986 20528
rect 23768 20516 23796 20547
rect 24854 20544 24860 20596
rect 24912 20584 24918 20596
rect 27338 20584 27344 20596
rect 24912 20556 27344 20584
rect 24912 20544 24918 20556
rect 27338 20544 27344 20556
rect 27396 20544 27402 20596
rect 27706 20544 27712 20596
rect 27764 20584 27770 20596
rect 29825 20587 29883 20593
rect 29825 20584 29837 20587
rect 27764 20556 29837 20584
rect 27764 20544 27770 20556
rect 29825 20553 29837 20556
rect 29871 20553 29883 20587
rect 37642 20584 37648 20596
rect 29825 20547 29883 20553
rect 29932 20556 37648 20584
rect 26970 20516 26976 20528
rect 23768 20488 26976 20516
rect 26970 20476 26976 20488
rect 27028 20476 27034 20528
rect 27246 20476 27252 20528
rect 27304 20516 27310 20528
rect 27430 20516 27436 20528
rect 27304 20488 27436 20516
rect 27304 20476 27310 20488
rect 27430 20476 27436 20488
rect 27488 20476 27494 20528
rect 28534 20476 28540 20528
rect 28592 20516 28598 20528
rect 29932 20516 29960 20556
rect 37642 20544 37648 20556
rect 37700 20544 37706 20596
rect 38838 20544 38844 20596
rect 38896 20584 38902 20596
rect 40405 20587 40463 20593
rect 38896 20556 40080 20584
rect 38896 20544 38902 20556
rect 28592 20488 29960 20516
rect 28592 20476 28598 20488
rect 30374 20476 30380 20528
rect 30432 20516 30438 20528
rect 30834 20516 30840 20528
rect 30432 20488 30840 20516
rect 30432 20476 30438 20488
rect 30834 20476 30840 20488
rect 30892 20476 30898 20528
rect 32490 20516 32496 20528
rect 31680 20488 32496 20516
rect 18325 20451 18383 20457
rect 18325 20448 18337 20451
rect 17920 20420 18337 20448
rect 17920 20408 17926 20420
rect 18325 20417 18337 20420
rect 18371 20417 18383 20451
rect 18325 20411 18383 20417
rect 18414 20408 18420 20460
rect 18472 20448 18478 20460
rect 19150 20448 19156 20460
rect 18472 20420 18517 20448
rect 19111 20420 19156 20448
rect 18472 20408 18478 20420
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 22370 20448 22376 20460
rect 22331 20420 22376 20448
rect 22370 20408 22376 20420
rect 22428 20408 22434 20460
rect 24305 20451 24363 20457
rect 24305 20417 24317 20451
rect 24351 20417 24363 20451
rect 27338 20448 27344 20460
rect 27299 20420 27344 20448
rect 24305 20411 24363 20417
rect 18509 20383 18567 20389
rect 17052 20352 18276 20380
rect 16040 20312 16068 20340
rect 18248 20324 18276 20352
rect 18509 20349 18521 20383
rect 18555 20349 18567 20383
rect 18509 20343 18567 20349
rect 17862 20312 17868 20324
rect 16040 20284 17868 20312
rect 17862 20272 17868 20284
rect 17920 20272 17926 20324
rect 18230 20272 18236 20324
rect 18288 20312 18294 20324
rect 18524 20312 18552 20343
rect 18598 20340 18604 20392
rect 18656 20380 18662 20392
rect 20714 20380 20720 20392
rect 18656 20352 18701 20380
rect 20675 20352 20720 20380
rect 18656 20340 18662 20352
rect 20714 20340 20720 20352
rect 20772 20340 20778 20392
rect 24320 20380 24348 20411
rect 27338 20408 27344 20420
rect 27396 20408 27402 20460
rect 27522 20408 27528 20460
rect 27580 20448 27586 20460
rect 28629 20451 28687 20457
rect 27580 20420 27625 20448
rect 27580 20408 27586 20420
rect 28629 20417 28641 20451
rect 28675 20448 28687 20451
rect 29454 20448 29460 20460
rect 28675 20420 29460 20448
rect 28675 20417 28687 20420
rect 28629 20411 28687 20417
rect 29454 20408 29460 20420
rect 29512 20408 29518 20460
rect 31389 20451 31447 20457
rect 31389 20448 31401 20451
rect 30760 20420 31401 20448
rect 28810 20380 28816 20392
rect 24320 20352 28816 20380
rect 28810 20340 28816 20352
rect 28868 20340 28874 20392
rect 30760 20380 30788 20420
rect 31389 20417 31401 20420
rect 31435 20448 31447 20451
rect 31570 20448 31576 20460
rect 31435 20420 31576 20448
rect 31435 20417 31447 20420
rect 31389 20411 31447 20417
rect 31570 20408 31576 20420
rect 31628 20408 31634 20460
rect 31680 20457 31708 20488
rect 32490 20476 32496 20488
rect 32548 20516 32554 20528
rect 32674 20516 32680 20528
rect 32548 20488 32680 20516
rect 32548 20476 32554 20488
rect 32674 20476 32680 20488
rect 32732 20476 32738 20528
rect 33318 20476 33324 20528
rect 33376 20516 33382 20528
rect 36173 20519 36231 20525
rect 36173 20516 36185 20519
rect 33376 20488 36185 20516
rect 33376 20476 33382 20488
rect 36173 20485 36185 20488
rect 36219 20485 36231 20519
rect 36173 20479 36231 20485
rect 36906 20476 36912 20528
rect 36964 20516 36970 20528
rect 37737 20519 37795 20525
rect 37737 20516 37749 20519
rect 36964 20488 37749 20516
rect 36964 20476 36970 20488
rect 37737 20485 37749 20488
rect 37783 20485 37795 20519
rect 39942 20516 39948 20528
rect 37737 20479 37795 20485
rect 38764 20488 39948 20516
rect 31665 20451 31723 20457
rect 31665 20417 31677 20451
rect 31711 20417 31723 20451
rect 31665 20411 31723 20417
rect 32309 20451 32367 20457
rect 32309 20417 32321 20451
rect 32355 20448 32367 20451
rect 35989 20451 36047 20457
rect 35989 20448 36001 20451
rect 32355 20420 36001 20448
rect 32355 20417 32367 20420
rect 32309 20411 32367 20417
rect 35989 20417 36001 20420
rect 36035 20448 36047 20451
rect 36035 20420 37412 20448
rect 36035 20417 36047 20420
rect 35989 20411 36047 20417
rect 30484 20352 30788 20380
rect 25501 20315 25559 20321
rect 25501 20312 25513 20315
rect 18288 20284 22094 20312
rect 18288 20272 18294 20284
rect 15930 20204 15936 20256
rect 15988 20244 15994 20256
rect 16301 20247 16359 20253
rect 16301 20244 16313 20247
rect 15988 20216 16313 20244
rect 15988 20204 15994 20216
rect 16301 20213 16313 20216
rect 16347 20213 16359 20247
rect 16301 20207 16359 20213
rect 18141 20247 18199 20253
rect 18141 20213 18153 20247
rect 18187 20244 18199 20247
rect 19150 20244 19156 20256
rect 18187 20216 19156 20244
rect 18187 20213 18199 20216
rect 18141 20207 18199 20213
rect 19150 20204 19156 20216
rect 19208 20204 19214 20256
rect 22066 20244 22094 20284
rect 23308 20284 25513 20312
rect 23308 20244 23336 20284
rect 25501 20281 25513 20284
rect 25547 20281 25559 20315
rect 25501 20275 25559 20281
rect 27157 20315 27215 20321
rect 27157 20281 27169 20315
rect 27203 20312 27215 20315
rect 27614 20312 27620 20324
rect 27203 20284 27620 20312
rect 27203 20281 27215 20284
rect 27157 20275 27215 20281
rect 27614 20272 27620 20284
rect 27672 20272 27678 20324
rect 27706 20272 27712 20324
rect 27764 20312 27770 20324
rect 27764 20284 27809 20312
rect 27764 20272 27770 20284
rect 28626 20272 28632 20324
rect 28684 20312 28690 20324
rect 30484 20312 30512 20352
rect 30834 20340 30840 20392
rect 30892 20380 30898 20392
rect 32324 20380 32352 20411
rect 30892 20352 32352 20380
rect 30892 20340 30898 20352
rect 33962 20340 33968 20392
rect 34020 20380 34026 20392
rect 36265 20383 36323 20389
rect 36265 20380 36277 20383
rect 34020 20352 36277 20380
rect 34020 20340 34026 20352
rect 36265 20349 36277 20352
rect 36311 20380 36323 20383
rect 36538 20380 36544 20392
rect 36311 20352 36544 20380
rect 36311 20349 36323 20352
rect 36265 20343 36323 20349
rect 36538 20340 36544 20352
rect 36596 20380 36602 20392
rect 37182 20380 37188 20392
rect 36596 20352 37188 20380
rect 36596 20340 36602 20352
rect 37182 20340 37188 20352
rect 37240 20340 37246 20392
rect 37384 20380 37412 20420
rect 37458 20408 37464 20460
rect 37516 20448 37522 20460
rect 38378 20448 38384 20460
rect 37516 20420 38384 20448
rect 37516 20408 37522 20420
rect 38378 20408 38384 20420
rect 38436 20408 38442 20460
rect 38764 20380 38792 20488
rect 39942 20476 39948 20488
rect 40000 20476 40006 20528
rect 40052 20516 40080 20556
rect 40405 20553 40417 20587
rect 40451 20584 40463 20587
rect 40494 20584 40500 20596
rect 40451 20556 40500 20584
rect 40451 20553 40463 20556
rect 40405 20547 40463 20553
rect 40494 20544 40500 20556
rect 40552 20544 40558 20596
rect 48314 20584 48320 20596
rect 40601 20556 48320 20584
rect 40601 20516 40629 20556
rect 48314 20544 48320 20556
rect 48372 20544 48378 20596
rect 50154 20544 50160 20596
rect 50212 20584 50218 20596
rect 50341 20587 50399 20593
rect 50341 20584 50353 20587
rect 50212 20556 50353 20584
rect 50212 20544 50218 20556
rect 50341 20553 50353 20556
rect 50387 20553 50399 20587
rect 50341 20547 50399 20553
rect 54294 20544 54300 20596
rect 54352 20584 54358 20596
rect 57606 20584 57612 20596
rect 54352 20556 57612 20584
rect 54352 20544 54358 20556
rect 57606 20544 57612 20556
rect 57664 20544 57670 20596
rect 48038 20516 48044 20528
rect 40052 20488 40629 20516
rect 45388 20488 48044 20516
rect 38841 20451 38899 20457
rect 38841 20417 38853 20451
rect 38887 20448 38899 20451
rect 38930 20448 38936 20460
rect 38887 20420 38936 20448
rect 38887 20417 38899 20420
rect 38841 20411 38899 20417
rect 38930 20408 38936 20420
rect 38988 20408 38994 20460
rect 40310 20448 40316 20460
rect 40271 20420 40316 20448
rect 40310 20408 40316 20420
rect 40368 20408 40374 20460
rect 40497 20451 40555 20457
rect 40497 20417 40509 20451
rect 40543 20448 40555 20451
rect 43438 20448 43444 20460
rect 40543 20420 43444 20448
rect 40543 20417 40555 20420
rect 40497 20411 40555 20417
rect 43438 20408 43444 20420
rect 43496 20408 43502 20460
rect 45388 20457 45416 20488
rect 48038 20476 48044 20488
rect 48096 20476 48102 20528
rect 48222 20476 48228 20528
rect 48280 20516 48286 20528
rect 48280 20488 55214 20516
rect 48280 20476 48286 20488
rect 45373 20451 45431 20457
rect 45373 20417 45385 20451
rect 45419 20417 45431 20451
rect 45554 20448 45560 20460
rect 45515 20420 45560 20448
rect 45373 20411 45431 20417
rect 45554 20408 45560 20420
rect 45612 20408 45618 20460
rect 45649 20451 45707 20457
rect 45649 20417 45661 20451
rect 45695 20417 45707 20451
rect 45649 20411 45707 20417
rect 37384 20352 38792 20380
rect 39025 20383 39083 20389
rect 39025 20349 39037 20383
rect 39071 20349 39083 20383
rect 45664 20380 45692 20411
rect 45738 20408 45744 20460
rect 45796 20448 45802 20460
rect 45796 20420 45841 20448
rect 45796 20408 45802 20420
rect 49694 20408 49700 20460
rect 49752 20448 49758 20460
rect 49789 20451 49847 20457
rect 49789 20448 49801 20451
rect 49752 20420 49801 20448
rect 49752 20408 49758 20420
rect 49789 20417 49801 20420
rect 49835 20417 49847 20451
rect 49970 20448 49976 20460
rect 49931 20420 49976 20448
rect 49789 20411 49847 20417
rect 49970 20408 49976 20420
rect 50028 20408 50034 20460
rect 50065 20451 50123 20457
rect 50065 20417 50077 20451
rect 50111 20417 50123 20451
rect 50065 20411 50123 20417
rect 50157 20451 50215 20457
rect 50157 20417 50169 20451
rect 50203 20448 50215 20451
rect 50706 20448 50712 20460
rect 50203 20420 50712 20448
rect 50203 20417 50215 20420
rect 50157 20411 50215 20417
rect 50080 20380 50108 20411
rect 50706 20408 50712 20420
rect 50764 20448 50770 20460
rect 50764 20420 51856 20448
rect 50764 20408 50770 20420
rect 51718 20380 51724 20392
rect 45664 20352 45876 20380
rect 50080 20352 51724 20380
rect 39025 20343 39083 20349
rect 28684 20284 30512 20312
rect 28684 20272 28690 20284
rect 30558 20272 30564 20324
rect 30616 20312 30622 20324
rect 31665 20315 31723 20321
rect 31665 20312 31677 20315
rect 30616 20284 31677 20312
rect 30616 20272 30622 20284
rect 31665 20281 31677 20284
rect 31711 20281 31723 20315
rect 31665 20275 31723 20281
rect 35713 20315 35771 20321
rect 35713 20281 35725 20315
rect 35759 20312 35771 20315
rect 38838 20312 38844 20324
rect 35759 20284 38844 20312
rect 35759 20281 35771 20284
rect 35713 20275 35771 20281
rect 38838 20272 38844 20284
rect 38896 20272 38902 20324
rect 22066 20216 23336 20244
rect 24118 20204 24124 20256
rect 24176 20244 24182 20256
rect 33505 20247 33563 20253
rect 33505 20244 33517 20247
rect 24176 20216 33517 20244
rect 24176 20204 24182 20216
rect 33505 20213 33517 20216
rect 33551 20213 33563 20247
rect 33505 20207 33563 20213
rect 35894 20204 35900 20256
rect 35952 20244 35958 20256
rect 36630 20244 36636 20256
rect 35952 20216 36636 20244
rect 35952 20204 35958 20216
rect 36630 20204 36636 20216
rect 36688 20244 36694 20256
rect 38010 20244 38016 20256
rect 36688 20216 38016 20244
rect 36688 20204 36694 20216
rect 38010 20204 38016 20216
rect 38068 20204 38074 20256
rect 38102 20204 38108 20256
rect 38160 20244 38166 20256
rect 39040 20244 39068 20343
rect 45848 20312 45876 20352
rect 51718 20340 51724 20352
rect 51776 20340 51782 20392
rect 51828 20380 51856 20420
rect 52362 20408 52368 20460
rect 52420 20448 52426 20460
rect 53190 20457 53196 20460
rect 52917 20451 52975 20457
rect 52917 20448 52929 20451
rect 52420 20420 52929 20448
rect 52420 20408 52426 20420
rect 52917 20417 52929 20420
rect 52963 20417 52975 20451
rect 52917 20411 52975 20417
rect 53184 20411 53196 20457
rect 53248 20448 53254 20460
rect 53248 20420 53284 20448
rect 53190 20408 53196 20411
rect 53248 20408 53254 20420
rect 52546 20380 52552 20392
rect 51828 20352 52552 20380
rect 52546 20340 52552 20352
rect 52604 20340 52610 20392
rect 52086 20312 52092 20324
rect 45848 20284 52092 20312
rect 52086 20272 52092 20284
rect 52144 20272 52150 20324
rect 38160 20216 39068 20244
rect 38160 20204 38166 20216
rect 45830 20204 45836 20256
rect 45888 20244 45894 20256
rect 45925 20247 45983 20253
rect 45925 20244 45937 20247
rect 45888 20216 45937 20244
rect 45888 20204 45894 20216
rect 45925 20213 45937 20216
rect 45971 20213 45983 20247
rect 45925 20207 45983 20213
rect 51810 20204 51816 20256
rect 51868 20244 51874 20256
rect 52362 20244 52368 20256
rect 51868 20216 52368 20244
rect 51868 20204 51874 20216
rect 52362 20204 52368 20216
rect 52420 20204 52426 20256
rect 54294 20244 54300 20256
rect 54255 20216 54300 20244
rect 54294 20204 54300 20216
rect 54352 20204 54358 20256
rect 55186 20244 55214 20488
rect 56778 20244 56784 20256
rect 55186 20216 56784 20244
rect 56778 20204 56784 20216
rect 56836 20204 56842 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 15194 20000 15200 20052
rect 15252 20040 15258 20052
rect 17129 20043 17187 20049
rect 17129 20040 17141 20043
rect 15252 20012 17141 20040
rect 15252 20000 15258 20012
rect 17129 20009 17141 20012
rect 17175 20009 17187 20043
rect 20990 20040 20996 20052
rect 20951 20012 20996 20040
rect 17129 20003 17187 20009
rect 20990 20000 20996 20012
rect 21048 20000 21054 20052
rect 22278 20000 22284 20052
rect 22336 20040 22342 20052
rect 24673 20043 24731 20049
rect 24673 20040 24685 20043
rect 22336 20012 24685 20040
rect 22336 20000 22342 20012
rect 24673 20009 24685 20012
rect 24719 20009 24731 20043
rect 26510 20040 26516 20052
rect 26471 20012 26516 20040
rect 24673 20003 24731 20009
rect 26510 20000 26516 20012
rect 26568 20000 26574 20052
rect 28534 20040 28540 20052
rect 28495 20012 28540 20040
rect 28534 20000 28540 20012
rect 28592 20000 28598 20052
rect 29089 20043 29147 20049
rect 29089 20009 29101 20043
rect 29135 20040 29147 20043
rect 31846 20040 31852 20052
rect 29135 20012 31852 20040
rect 29135 20009 29147 20012
rect 29089 20003 29147 20009
rect 31846 20000 31852 20012
rect 31904 20040 31910 20052
rect 32306 20040 32312 20052
rect 31904 20012 32312 20040
rect 31904 20000 31910 20012
rect 32306 20000 32312 20012
rect 32364 20000 32370 20052
rect 34146 20000 34152 20052
rect 34204 20040 34210 20052
rect 39666 20040 39672 20052
rect 34204 20012 39672 20040
rect 34204 20000 34210 20012
rect 39666 20000 39672 20012
rect 39724 20000 39730 20052
rect 40218 20040 40224 20052
rect 40179 20012 40224 20040
rect 40218 20000 40224 20012
rect 40276 20000 40282 20052
rect 41230 20000 41236 20052
rect 41288 20040 41294 20052
rect 58618 20040 58624 20052
rect 41288 20012 58624 20040
rect 41288 20000 41294 20012
rect 58618 20000 58624 20012
rect 58676 20000 58682 20052
rect 17770 19932 17776 19984
rect 17828 19972 17834 19984
rect 20254 19972 20260 19984
rect 17828 19944 20260 19972
rect 17828 19932 17834 19944
rect 20254 19932 20260 19944
rect 20312 19932 20318 19984
rect 27338 19932 27344 19984
rect 27396 19972 27402 19984
rect 27890 19972 27896 19984
rect 27396 19944 27896 19972
rect 27396 19932 27402 19944
rect 27890 19932 27896 19944
rect 27948 19972 27954 19984
rect 32677 19975 32735 19981
rect 32677 19972 32689 19975
rect 27948 19944 32689 19972
rect 27948 19932 27954 19944
rect 32677 19941 32689 19944
rect 32723 19941 32735 19975
rect 32677 19935 32735 19941
rect 39592 19944 46336 19972
rect 20438 19904 20444 19916
rect 18892 19876 20444 19904
rect 1486 19796 1492 19848
rect 1544 19836 1550 19848
rect 1581 19839 1639 19845
rect 1581 19836 1593 19839
rect 1544 19808 1593 19836
rect 1544 19796 1550 19808
rect 1581 19805 1593 19808
rect 1627 19805 1639 19839
rect 15930 19836 15936 19848
rect 15891 19808 15936 19836
rect 1581 19799 1639 19805
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 18892 19845 18920 19876
rect 20438 19864 20444 19876
rect 20496 19864 20502 19916
rect 22370 19864 22376 19916
rect 22428 19904 22434 19916
rect 22649 19907 22707 19913
rect 22649 19904 22661 19907
rect 22428 19876 22661 19904
rect 22428 19864 22434 19876
rect 22649 19873 22661 19876
rect 22695 19873 22707 19907
rect 27706 19904 27712 19916
rect 22649 19867 22707 19873
rect 24504 19876 27712 19904
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19805 18751 19839
rect 18693 19799 18751 19805
rect 18877 19839 18935 19845
rect 18877 19805 18889 19839
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 1854 19768 1860 19780
rect 1815 19740 1860 19768
rect 1854 19728 1860 19740
rect 1912 19728 1918 19780
rect 17862 19728 17868 19780
rect 17920 19768 17926 19780
rect 18414 19768 18420 19780
rect 17920 19740 18420 19768
rect 17920 19728 17926 19740
rect 18414 19728 18420 19740
rect 18472 19728 18478 19780
rect 18708 19768 18736 19799
rect 18966 19796 18972 19848
rect 19024 19836 19030 19848
rect 19797 19839 19855 19845
rect 19797 19836 19809 19839
rect 19024 19808 19809 19836
rect 19024 19796 19030 19808
rect 19797 19805 19809 19808
rect 19843 19805 19855 19839
rect 24504 19836 24532 19876
rect 27706 19864 27712 19876
rect 27764 19864 27770 19916
rect 29181 19907 29239 19913
rect 29181 19873 29193 19907
rect 29227 19904 29239 19907
rect 29454 19904 29460 19916
rect 29227 19876 29460 19904
rect 29227 19873 29239 19876
rect 29181 19867 29239 19873
rect 29454 19864 29460 19876
rect 29512 19864 29518 19916
rect 30466 19904 30472 19916
rect 30427 19876 30472 19904
rect 30466 19864 30472 19876
rect 30524 19864 30530 19916
rect 35989 19907 36047 19913
rect 35989 19904 36001 19907
rect 31496 19876 36001 19904
rect 24670 19836 24676 19848
rect 19797 19799 19855 19805
rect 22664 19808 24532 19836
rect 24631 19808 24676 19836
rect 22664 19780 22692 19808
rect 24670 19796 24676 19808
rect 24728 19796 24734 19848
rect 24762 19796 24768 19848
rect 24820 19836 24826 19848
rect 24857 19839 24915 19845
rect 24857 19836 24869 19839
rect 24820 19808 24869 19836
rect 24820 19796 24826 19808
rect 24857 19805 24869 19808
rect 24903 19805 24915 19839
rect 25314 19836 25320 19848
rect 25275 19808 25320 19836
rect 24857 19799 24915 19805
rect 25314 19796 25320 19808
rect 25372 19796 25378 19848
rect 28442 19796 28448 19848
rect 28500 19836 28506 19848
rect 28662 19839 28720 19845
rect 28662 19836 28674 19839
rect 28500 19808 28674 19836
rect 28500 19796 28506 19808
rect 28662 19805 28674 19808
rect 28708 19805 28720 19839
rect 28662 19799 28720 19805
rect 28810 19796 28816 19848
rect 28868 19836 28874 19848
rect 30377 19839 30435 19845
rect 28868 19808 29960 19836
rect 28868 19796 28874 19808
rect 21266 19768 21272 19780
rect 18708 19740 21272 19768
rect 21266 19728 21272 19740
rect 21324 19768 21330 19780
rect 21818 19768 21824 19780
rect 21324 19740 21824 19768
rect 21324 19728 21330 19740
rect 21818 19728 21824 19740
rect 21876 19728 21882 19780
rect 22646 19728 22652 19780
rect 22704 19728 22710 19780
rect 22916 19771 22974 19777
rect 22916 19737 22928 19771
rect 22962 19768 22974 19771
rect 25498 19768 25504 19780
rect 22962 19740 25504 19768
rect 22962 19737 22974 19740
rect 22916 19731 22974 19737
rect 25498 19728 25504 19740
rect 25556 19728 25562 19780
rect 29730 19768 29736 19780
rect 28552 19740 29592 19768
rect 29691 19740 29736 19768
rect 18785 19703 18843 19709
rect 18785 19669 18797 19703
rect 18831 19700 18843 19703
rect 19334 19700 19340 19712
rect 18831 19672 19340 19700
rect 18831 19669 18843 19672
rect 18785 19663 18843 19669
rect 19334 19660 19340 19672
rect 19392 19660 19398 19712
rect 24029 19703 24087 19709
rect 24029 19669 24041 19703
rect 24075 19700 24087 19703
rect 28552 19700 28580 19740
rect 28718 19700 28724 19712
rect 24075 19672 28580 19700
rect 28679 19672 28724 19700
rect 24075 19669 24087 19672
rect 24029 19663 24087 19669
rect 28718 19660 28724 19672
rect 28776 19660 28782 19712
rect 29564 19700 29592 19740
rect 29730 19728 29736 19740
rect 29788 19728 29794 19780
rect 29822 19700 29828 19712
rect 29564 19672 29828 19700
rect 29822 19660 29828 19672
rect 29880 19660 29886 19712
rect 29932 19700 29960 19808
rect 30377 19805 30389 19839
rect 30423 19805 30435 19839
rect 30742 19836 30748 19848
rect 30703 19808 30748 19836
rect 30377 19799 30435 19805
rect 30392 19768 30420 19799
rect 30742 19796 30748 19808
rect 30800 19796 30806 19848
rect 30929 19839 30987 19845
rect 30929 19805 30941 19839
rect 30975 19836 30987 19839
rect 31110 19836 31116 19848
rect 30975 19808 31116 19836
rect 30975 19805 30987 19808
rect 30929 19799 30987 19805
rect 31110 19796 31116 19808
rect 31168 19796 31174 19848
rect 31496 19845 31524 19876
rect 35989 19873 36001 19876
rect 36035 19873 36047 19907
rect 37550 19904 37556 19916
rect 35989 19867 36047 19873
rect 37200 19876 37556 19904
rect 31481 19839 31539 19845
rect 31481 19805 31493 19839
rect 31527 19805 31539 19839
rect 34882 19836 34888 19848
rect 34843 19808 34888 19836
rect 31481 19799 31539 19805
rect 34882 19796 34888 19808
rect 34940 19836 34946 19848
rect 37200 19836 37228 19876
rect 37550 19864 37556 19876
rect 37608 19904 37614 19916
rect 39025 19907 39083 19913
rect 39025 19904 39037 19907
rect 37608 19876 39037 19904
rect 37608 19864 37614 19876
rect 39025 19873 39037 19876
rect 39071 19873 39083 19907
rect 39025 19867 39083 19873
rect 34940 19808 37228 19836
rect 34940 19796 34946 19808
rect 37274 19796 37280 19848
rect 37332 19836 37338 19848
rect 37642 19836 37648 19848
rect 37332 19808 37648 19836
rect 37332 19796 37338 19808
rect 37642 19796 37648 19808
rect 37700 19796 37706 19848
rect 37734 19796 37740 19848
rect 37792 19836 37798 19848
rect 37921 19839 37979 19845
rect 37921 19836 37933 19839
rect 37792 19808 37933 19836
rect 37792 19796 37798 19808
rect 37921 19805 37933 19808
rect 37967 19805 37979 19839
rect 37921 19799 37979 19805
rect 38010 19796 38016 19848
rect 38068 19836 38074 19848
rect 39592 19836 39620 19944
rect 41322 19864 41328 19916
rect 41380 19904 41386 19916
rect 41509 19907 41567 19913
rect 41509 19904 41521 19907
rect 41380 19876 41521 19904
rect 41380 19864 41386 19876
rect 41509 19873 41521 19876
rect 41555 19904 41567 19907
rect 41874 19904 41880 19916
rect 41555 19876 41880 19904
rect 41555 19873 41567 19876
rect 41509 19867 41567 19873
rect 41874 19864 41880 19876
rect 41932 19864 41938 19916
rect 45922 19904 45928 19916
rect 45883 19876 45928 19904
rect 45922 19864 45928 19876
rect 45980 19864 45986 19916
rect 46308 19913 46336 19944
rect 46382 19932 46388 19984
rect 46440 19972 46446 19984
rect 46440 19944 55214 19972
rect 46440 19932 46446 19944
rect 46293 19907 46351 19913
rect 46293 19873 46305 19907
rect 46339 19873 46351 19907
rect 52641 19907 52699 19913
rect 46293 19867 46351 19873
rect 48286 19876 52316 19904
rect 38068 19808 39620 19836
rect 38068 19796 38074 19808
rect 39666 19796 39672 19848
rect 39724 19836 39730 19848
rect 40129 19839 40187 19845
rect 40129 19836 40141 19839
rect 39724 19808 40141 19836
rect 39724 19796 39730 19808
rect 40129 19805 40141 19808
rect 40175 19805 40187 19839
rect 40129 19799 40187 19805
rect 40586 19796 40592 19848
rect 40644 19836 40650 19848
rect 41046 19836 41052 19848
rect 40644 19808 41052 19836
rect 40644 19796 40650 19808
rect 41046 19796 41052 19808
rect 41104 19796 41110 19848
rect 41230 19836 41236 19848
rect 41191 19808 41236 19836
rect 41230 19796 41236 19808
rect 41288 19796 41294 19848
rect 45830 19836 45836 19848
rect 45791 19808 45836 19836
rect 45830 19796 45836 19808
rect 45888 19796 45894 19848
rect 46198 19836 46204 19848
rect 46159 19808 46204 19836
rect 46198 19796 46204 19808
rect 46256 19796 46262 19848
rect 48286 19836 48314 19876
rect 46308 19808 48314 19836
rect 31386 19768 31392 19780
rect 30392 19740 31392 19768
rect 31386 19728 31392 19740
rect 31444 19728 31450 19780
rect 45094 19728 45100 19780
rect 45152 19768 45158 19780
rect 45189 19771 45247 19777
rect 45189 19768 45201 19771
rect 45152 19740 45201 19768
rect 45152 19728 45158 19740
rect 45189 19737 45201 19740
rect 45235 19737 45247 19771
rect 45189 19731 45247 19737
rect 45370 19728 45376 19780
rect 45428 19768 45434 19780
rect 46308 19768 46336 19808
rect 49970 19796 49976 19848
rect 50028 19836 50034 19848
rect 52181 19839 52239 19845
rect 52181 19836 52193 19839
rect 50028 19808 52193 19836
rect 50028 19796 50034 19808
rect 52181 19805 52193 19808
rect 52227 19805 52239 19839
rect 52288 19836 52316 19876
rect 52641 19873 52653 19907
rect 52687 19904 52699 19907
rect 54294 19904 54300 19916
rect 52687 19876 54300 19904
rect 52687 19873 52699 19876
rect 52641 19867 52699 19873
rect 54294 19864 54300 19876
rect 54352 19864 54358 19916
rect 55186 19904 55214 19944
rect 57333 19907 57391 19913
rect 57333 19904 57345 19907
rect 55186 19876 57345 19904
rect 57333 19873 57345 19876
rect 57379 19873 57391 19907
rect 58158 19904 58164 19916
rect 58119 19876 58164 19904
rect 57333 19867 57391 19873
rect 58158 19864 58164 19876
rect 58216 19864 58222 19916
rect 57885 19839 57943 19845
rect 57885 19836 57897 19839
rect 52288 19808 57897 19836
rect 52181 19799 52239 19805
rect 57885 19805 57897 19808
rect 57931 19805 57943 19839
rect 57885 19799 57943 19805
rect 45428 19740 46336 19768
rect 45428 19728 45434 19740
rect 47118 19728 47124 19780
rect 47176 19768 47182 19780
rect 52273 19771 52331 19777
rect 52273 19768 52285 19771
rect 47176 19740 52285 19768
rect 47176 19728 47182 19740
rect 52273 19737 52285 19740
rect 52319 19737 52331 19771
rect 52273 19731 52331 19737
rect 52362 19728 52368 19780
rect 52420 19768 52426 19780
rect 52546 19777 52552 19780
rect 52503 19771 52552 19777
rect 52420 19740 52465 19768
rect 52420 19728 52426 19740
rect 52503 19737 52515 19771
rect 52549 19737 52552 19771
rect 52503 19731 52552 19737
rect 52546 19728 52552 19731
rect 52604 19768 52610 19780
rect 56318 19768 56324 19780
rect 52604 19740 56324 19768
rect 52604 19728 52610 19740
rect 56318 19728 56324 19740
rect 56376 19768 56382 19780
rect 56502 19768 56508 19780
rect 56376 19740 56508 19768
rect 56376 19728 56382 19740
rect 56502 19728 56508 19740
rect 56560 19728 56566 19780
rect 57054 19768 57060 19780
rect 57015 19740 57060 19768
rect 57054 19728 57060 19740
rect 57112 19728 57118 19780
rect 30650 19700 30656 19712
rect 29932 19672 30656 19700
rect 30650 19660 30656 19672
rect 30708 19660 30714 19712
rect 31110 19660 31116 19712
rect 31168 19700 31174 19712
rect 33778 19700 33784 19712
rect 31168 19672 33784 19700
rect 31168 19660 31174 19672
rect 33778 19660 33784 19672
rect 33836 19660 33842 19712
rect 34330 19660 34336 19712
rect 34388 19700 34394 19712
rect 46382 19700 46388 19712
rect 34388 19672 46388 19700
rect 34388 19660 34394 19672
rect 46382 19660 46388 19672
rect 46440 19660 46446 19712
rect 51997 19703 52055 19709
rect 51997 19669 52009 19703
rect 52043 19700 52055 19703
rect 52178 19700 52184 19712
rect 52043 19672 52184 19700
rect 52043 19669 52055 19672
rect 51997 19663 52055 19669
rect 52178 19660 52184 19672
rect 52236 19660 52242 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 15102 19496 15108 19508
rect 15063 19468 15108 19496
rect 15102 19456 15108 19468
rect 15160 19456 15166 19508
rect 18322 19456 18328 19508
rect 18380 19496 18386 19508
rect 18380 19468 18425 19496
rect 18380 19456 18386 19468
rect 19150 19456 19156 19508
rect 19208 19456 19214 19508
rect 25498 19496 25504 19508
rect 25459 19468 25504 19496
rect 25498 19456 25504 19468
rect 25556 19456 25562 19508
rect 27522 19496 27528 19508
rect 27356 19468 27528 19496
rect 17770 19428 17776 19440
rect 17420 19400 17776 19428
rect 17420 19369 17448 19400
rect 17770 19388 17776 19400
rect 17828 19388 17834 19440
rect 18049 19431 18107 19437
rect 18049 19397 18061 19431
rect 18095 19428 18107 19431
rect 18598 19428 18604 19440
rect 18095 19400 18604 19428
rect 18095 19397 18107 19400
rect 18049 19391 18107 19397
rect 18598 19388 18604 19400
rect 18656 19428 18662 19440
rect 18656 19400 19104 19428
rect 18656 19388 18662 19400
rect 17405 19363 17463 19369
rect 15028 19332 15516 19360
rect 14918 19252 14924 19304
rect 14976 19292 14982 19304
rect 15028 19292 15056 19332
rect 15488 19301 15516 19332
rect 17405 19329 17417 19363
rect 17451 19329 17463 19363
rect 17586 19360 17592 19372
rect 17547 19332 17592 19360
rect 17405 19323 17463 19329
rect 17586 19320 17592 19332
rect 17644 19320 17650 19372
rect 18230 19360 18236 19372
rect 18191 19332 18236 19360
rect 18230 19320 18236 19332
rect 18288 19320 18294 19372
rect 18414 19360 18420 19372
rect 18375 19332 18420 19360
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 14976 19264 15056 19292
rect 15289 19295 15347 19301
rect 14976 19252 14982 19264
rect 15289 19261 15301 19295
rect 15335 19261 15347 19295
rect 15289 19255 15347 19261
rect 15381 19295 15439 19301
rect 15381 19261 15393 19295
rect 15427 19261 15439 19295
rect 15381 19255 15439 19261
rect 15473 19295 15531 19301
rect 15473 19261 15485 19295
rect 15519 19261 15531 19295
rect 15473 19255 15531 19261
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 16390 19292 16396 19304
rect 15611 19264 16396 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 14734 19184 14740 19236
rect 14792 19224 14798 19236
rect 15304 19224 15332 19255
rect 14792 19196 15332 19224
rect 14792 19184 14798 19196
rect 15396 19156 15424 19255
rect 16390 19252 16396 19264
rect 16448 19252 16454 19304
rect 17497 19295 17555 19301
rect 17497 19261 17509 19295
rect 17543 19292 17555 19295
rect 18966 19292 18972 19304
rect 17543 19264 18972 19292
rect 17543 19261 17555 19264
rect 17497 19255 17555 19261
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19076 19292 19104 19400
rect 19168 19369 19196 19456
rect 23845 19431 23903 19437
rect 23845 19397 23857 19431
rect 23891 19428 23903 19431
rect 23891 19400 24624 19428
rect 23891 19397 23903 19400
rect 23845 19391 23903 19397
rect 19153 19363 19211 19369
rect 19153 19329 19165 19363
rect 19199 19329 19211 19363
rect 24118 19360 24124 19372
rect 19153 19323 19211 19329
rect 19260 19332 24124 19360
rect 19260 19292 19288 19332
rect 24118 19320 24124 19332
rect 24176 19320 24182 19372
rect 24302 19360 24308 19372
rect 24263 19332 24308 19360
rect 24302 19320 24308 19332
rect 24360 19320 24366 19372
rect 24596 19360 24624 19400
rect 27356 19372 27384 19468
rect 27522 19456 27528 19468
rect 27580 19456 27586 19508
rect 28534 19456 28540 19508
rect 28592 19496 28598 19508
rect 28592 19468 28677 19496
rect 28592 19456 28598 19468
rect 28649 19437 28677 19468
rect 34698 19456 34704 19508
rect 34756 19496 34762 19508
rect 36449 19499 36507 19505
rect 36449 19496 36461 19499
rect 34756 19468 36461 19496
rect 34756 19456 34762 19468
rect 36449 19465 36461 19468
rect 36495 19465 36507 19499
rect 36449 19459 36507 19465
rect 37461 19499 37519 19505
rect 37461 19465 37473 19499
rect 37507 19496 37519 19499
rect 37734 19496 37740 19508
rect 37507 19468 37740 19496
rect 37507 19465 37519 19468
rect 37461 19459 37519 19465
rect 37734 19456 37740 19468
rect 37792 19456 37798 19508
rect 40034 19456 40040 19508
rect 40092 19496 40098 19508
rect 45370 19496 45376 19508
rect 40092 19468 45048 19496
rect 45331 19468 45376 19496
rect 40092 19456 40098 19468
rect 28634 19431 28692 19437
rect 28634 19397 28646 19431
rect 28680 19397 28692 19431
rect 37366 19428 37372 19440
rect 28634 19391 28692 19397
rect 32324 19400 37372 19428
rect 27338 19360 27344 19372
rect 24596 19332 26234 19360
rect 27300 19332 27344 19360
rect 19076 19264 19288 19292
rect 22094 19252 22100 19304
rect 22152 19292 22158 19304
rect 22189 19295 22247 19301
rect 22189 19292 22201 19295
rect 22152 19264 22201 19292
rect 22152 19252 22158 19264
rect 22189 19261 22201 19264
rect 22235 19292 22247 19295
rect 22370 19292 22376 19304
rect 22235 19264 22376 19292
rect 22235 19261 22247 19264
rect 22189 19255 22247 19261
rect 22370 19252 22376 19264
rect 22428 19252 22434 19304
rect 22462 19252 22468 19304
rect 22520 19292 22526 19304
rect 22520 19264 22565 19292
rect 22520 19252 22526 19264
rect 21174 19224 21180 19236
rect 18432 19196 21180 19224
rect 18432 19156 18460 19196
rect 21174 19184 21180 19196
rect 21232 19184 21238 19236
rect 21266 19184 21272 19236
rect 21324 19224 21330 19236
rect 26206 19224 26234 19332
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 28258 19320 28264 19372
rect 28316 19360 28322 19372
rect 28353 19363 28411 19369
rect 28353 19360 28365 19363
rect 28316 19332 28365 19360
rect 28316 19320 28322 19332
rect 28353 19329 28365 19332
rect 28399 19329 28411 19363
rect 28534 19360 28540 19372
rect 28495 19332 28540 19360
rect 28353 19323 28411 19329
rect 28534 19320 28540 19332
rect 28592 19320 28598 19372
rect 28767 19363 28825 19369
rect 28767 19360 28779 19363
rect 28741 19329 28779 19360
rect 28813 19329 28825 19363
rect 28741 19323 28825 19329
rect 27430 19292 27436 19304
rect 27391 19264 27436 19292
rect 27430 19252 27436 19264
rect 27488 19252 27494 19304
rect 27525 19295 27583 19301
rect 27525 19261 27537 19295
rect 27571 19261 27583 19295
rect 27525 19255 27583 19261
rect 27540 19224 27568 19255
rect 27614 19252 27620 19304
rect 27672 19292 27678 19304
rect 27672 19264 27717 19292
rect 27672 19252 27678 19264
rect 27890 19224 27896 19236
rect 21324 19196 22094 19224
rect 26206 19196 27476 19224
rect 27540 19196 27896 19224
rect 21324 19184 21330 19196
rect 18598 19156 18604 19168
rect 15396 19128 18460 19156
rect 18559 19128 18604 19156
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 21358 19156 21364 19168
rect 21319 19128 21364 19156
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 22066 19156 22094 19196
rect 23382 19156 23388 19168
rect 22066 19128 23388 19156
rect 23382 19116 23388 19128
rect 23440 19116 23446 19168
rect 27154 19156 27160 19168
rect 27115 19128 27160 19156
rect 27154 19116 27160 19128
rect 27212 19116 27218 19168
rect 27448 19156 27476 19196
rect 27890 19184 27896 19196
rect 27948 19184 27954 19236
rect 28626 19184 28632 19236
rect 28684 19224 28690 19236
rect 28741 19224 28769 19323
rect 28994 19320 29000 19372
rect 29052 19360 29058 19372
rect 29454 19360 29460 19372
rect 29052 19332 29460 19360
rect 29052 19320 29058 19332
rect 29454 19320 29460 19332
rect 29512 19320 29518 19372
rect 29822 19320 29828 19372
rect 29880 19360 29886 19372
rect 32324 19369 32352 19400
rect 37366 19388 37372 19400
rect 37424 19428 37430 19440
rect 37550 19428 37556 19440
rect 37424 19400 37556 19428
rect 37424 19388 37430 19400
rect 37550 19388 37556 19400
rect 37608 19388 37614 19440
rect 37642 19388 37648 19440
rect 37700 19428 37706 19440
rect 37700 19400 41414 19428
rect 37700 19388 37706 19400
rect 32309 19363 32367 19369
rect 32309 19360 32321 19363
rect 29880 19332 32321 19360
rect 29880 19320 29886 19332
rect 32309 19329 32321 19332
rect 32355 19329 32367 19363
rect 32309 19323 32367 19329
rect 32582 19320 32588 19372
rect 32640 19360 32646 19372
rect 34698 19360 34704 19372
rect 32640 19332 34704 19360
rect 32640 19320 32646 19332
rect 34698 19320 34704 19332
rect 34756 19320 34762 19372
rect 34790 19320 34796 19372
rect 34848 19360 34854 19372
rect 35342 19369 35348 19372
rect 35069 19363 35127 19369
rect 35069 19360 35081 19363
rect 34848 19332 35081 19360
rect 34848 19320 34854 19332
rect 35069 19329 35081 19332
rect 35115 19329 35127 19363
rect 35069 19323 35127 19329
rect 35336 19323 35348 19369
rect 35400 19360 35406 19372
rect 37734 19360 37740 19372
rect 35400 19332 35436 19360
rect 37695 19332 37740 19360
rect 35342 19320 35348 19323
rect 35400 19320 35406 19332
rect 37734 19320 37740 19332
rect 37792 19320 37798 19372
rect 37829 19363 37887 19369
rect 37829 19329 37841 19363
rect 37875 19329 37887 19363
rect 37829 19323 37887 19329
rect 30650 19252 30656 19304
rect 30708 19292 30714 19304
rect 30708 19264 30753 19292
rect 30708 19252 30714 19264
rect 31294 19252 31300 19304
rect 31352 19292 31358 19304
rect 33413 19295 33471 19301
rect 33413 19292 33425 19295
rect 31352 19264 33425 19292
rect 31352 19252 31358 19264
rect 33413 19261 33425 19264
rect 33459 19261 33471 19295
rect 33413 19255 33471 19261
rect 36078 19252 36084 19304
rect 36136 19292 36142 19304
rect 37844 19292 37872 19323
rect 37918 19320 37924 19372
rect 37976 19360 37982 19372
rect 38105 19363 38163 19369
rect 37976 19332 38021 19360
rect 37976 19320 37982 19332
rect 38105 19329 38117 19363
rect 38151 19360 38163 19363
rect 38654 19360 38660 19372
rect 38151 19332 38660 19360
rect 38151 19329 38163 19332
rect 38105 19323 38163 19329
rect 38654 19320 38660 19332
rect 38712 19320 38718 19372
rect 38764 19369 38792 19400
rect 38749 19363 38807 19369
rect 38749 19329 38761 19363
rect 38795 19329 38807 19363
rect 39005 19363 39063 19369
rect 39005 19360 39017 19363
rect 38749 19323 38807 19329
rect 38856 19332 39017 19360
rect 38010 19292 38016 19304
rect 36136 19264 38016 19292
rect 36136 19252 36142 19264
rect 38010 19252 38016 19264
rect 38068 19252 38074 19304
rect 38378 19252 38384 19304
rect 38436 19292 38442 19304
rect 38856 19292 38884 19332
rect 39005 19329 39017 19332
rect 39051 19329 39063 19363
rect 41386 19360 41414 19400
rect 42610 19360 42616 19372
rect 41386 19332 42616 19360
rect 39005 19323 39063 19329
rect 42610 19320 42616 19332
rect 42668 19360 42674 19372
rect 43346 19360 43352 19372
rect 42668 19332 43352 19360
rect 42668 19320 42674 19332
rect 43346 19320 43352 19332
rect 43404 19360 43410 19372
rect 44266 19369 44272 19372
rect 43993 19363 44051 19369
rect 43993 19360 44005 19363
rect 43404 19332 44005 19360
rect 43404 19320 43410 19332
rect 43993 19329 44005 19332
rect 44039 19329 44051 19363
rect 43993 19323 44051 19329
rect 44260 19323 44272 19369
rect 44324 19360 44330 19372
rect 45020 19360 45048 19468
rect 45370 19456 45376 19468
rect 45428 19456 45434 19508
rect 46198 19456 46204 19508
rect 46256 19496 46262 19508
rect 52365 19499 52423 19505
rect 46256 19468 52316 19496
rect 46256 19456 46262 19468
rect 45094 19388 45100 19440
rect 45152 19428 45158 19440
rect 47118 19428 47124 19440
rect 45152 19400 47124 19428
rect 45152 19388 45158 19400
rect 47118 19388 47124 19400
rect 47176 19388 47182 19440
rect 49970 19360 49976 19372
rect 44324 19332 44360 19360
rect 45020 19332 49976 19360
rect 44266 19320 44272 19323
rect 44324 19320 44330 19332
rect 49970 19320 49976 19332
rect 50028 19320 50034 19372
rect 52178 19360 52184 19372
rect 52139 19332 52184 19360
rect 52178 19320 52184 19332
rect 52236 19320 52242 19372
rect 52288 19360 52316 19468
rect 52365 19465 52377 19499
rect 52411 19496 52423 19499
rect 53190 19496 53196 19508
rect 52411 19468 53196 19496
rect 52411 19465 52423 19468
rect 52365 19459 52423 19465
rect 53190 19456 53196 19468
rect 53248 19456 53254 19508
rect 56965 19499 57023 19505
rect 56965 19465 56977 19499
rect 57011 19496 57023 19499
rect 58066 19496 58072 19508
rect 57011 19468 58072 19496
rect 57011 19465 57023 19468
rect 56965 19459 57023 19465
rect 58066 19456 58072 19468
rect 58124 19456 58130 19508
rect 52454 19388 52460 19440
rect 52512 19428 52518 19440
rect 52512 19400 57100 19428
rect 52512 19388 52518 19400
rect 53190 19360 53196 19372
rect 52288 19332 53196 19360
rect 53190 19320 53196 19332
rect 53248 19320 53254 19372
rect 56778 19360 56784 19372
rect 56739 19332 56784 19360
rect 56778 19320 56784 19332
rect 56836 19320 56842 19372
rect 57072 19369 57100 19400
rect 57057 19363 57115 19369
rect 57057 19329 57069 19363
rect 57103 19329 57115 19363
rect 57057 19323 57115 19329
rect 51994 19292 52000 19304
rect 38436 19264 38884 19292
rect 51955 19264 52000 19292
rect 38436 19252 38442 19264
rect 51994 19252 52000 19264
rect 52052 19252 52058 19304
rect 28684 19196 28769 19224
rect 28905 19227 28963 19233
rect 28684 19184 28690 19196
rect 28905 19193 28917 19227
rect 28951 19224 28963 19227
rect 29086 19224 29092 19236
rect 28951 19196 29092 19224
rect 28951 19193 28963 19196
rect 28905 19187 28963 19193
rect 29086 19184 29092 19196
rect 29144 19184 29150 19236
rect 31110 19224 31116 19236
rect 30392 19196 31116 19224
rect 30392 19156 30420 19196
rect 31110 19184 31116 19196
rect 31168 19224 31174 19236
rect 34882 19224 34888 19236
rect 31168 19196 34888 19224
rect 31168 19184 31174 19196
rect 34882 19184 34888 19196
rect 34940 19184 34946 19236
rect 43438 19224 43444 19236
rect 39684 19196 43444 19224
rect 27448 19128 30420 19156
rect 30466 19116 30472 19168
rect 30524 19156 30530 19168
rect 32766 19156 32772 19168
rect 30524 19128 32772 19156
rect 30524 19116 30530 19128
rect 32766 19116 32772 19128
rect 32824 19116 32830 19168
rect 33594 19116 33600 19168
rect 33652 19156 33658 19168
rect 33778 19156 33784 19168
rect 33652 19128 33784 19156
rect 33652 19116 33658 19128
rect 33778 19116 33784 19128
rect 33836 19116 33842 19168
rect 36538 19116 36544 19168
rect 36596 19156 36602 19168
rect 39684 19156 39712 19196
rect 43438 19184 43444 19196
rect 43496 19184 43502 19236
rect 46198 19184 46204 19236
rect 46256 19224 46262 19236
rect 58986 19224 58992 19236
rect 46256 19196 58992 19224
rect 46256 19184 46262 19196
rect 58986 19184 58992 19196
rect 59044 19184 59050 19236
rect 36596 19128 39712 19156
rect 36596 19116 36602 19128
rect 39758 19116 39764 19168
rect 39816 19156 39822 19168
rect 39942 19156 39948 19168
rect 39816 19128 39948 19156
rect 39816 19116 39822 19128
rect 39942 19116 39948 19128
rect 40000 19156 40006 19168
rect 40129 19159 40187 19165
rect 40129 19156 40141 19159
rect 40000 19128 40141 19156
rect 40000 19116 40006 19128
rect 40129 19125 40141 19128
rect 40175 19125 40187 19159
rect 43456 19156 43484 19184
rect 44358 19156 44364 19168
rect 43456 19128 44364 19156
rect 40129 19119 40187 19125
rect 44358 19116 44364 19128
rect 44416 19116 44422 19168
rect 56781 19159 56839 19165
rect 56781 19125 56793 19159
rect 56827 19156 56839 19159
rect 56962 19156 56968 19168
rect 56827 19128 56968 19156
rect 56827 19125 56839 19128
rect 56781 19119 56839 19125
rect 56962 19116 56968 19128
rect 57020 19116 57026 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 10778 18952 10784 18964
rect 10739 18924 10784 18952
rect 10778 18912 10784 18924
rect 10836 18912 10842 18964
rect 16206 18912 16212 18964
rect 16264 18952 16270 18964
rect 17954 18952 17960 18964
rect 16264 18924 17960 18952
rect 16264 18912 16270 18924
rect 17954 18912 17960 18924
rect 18012 18952 18018 18964
rect 18322 18952 18328 18964
rect 18012 18924 18328 18952
rect 18012 18912 18018 18924
rect 18322 18912 18328 18924
rect 18380 18912 18386 18964
rect 25130 18952 25136 18964
rect 18524 18924 20852 18952
rect 17218 18884 17224 18896
rect 11072 18856 17224 18884
rect 11072 18825 11100 18856
rect 17218 18844 17224 18856
rect 17276 18844 17282 18896
rect 11057 18819 11115 18825
rect 11057 18785 11069 18819
rect 11103 18785 11115 18819
rect 11057 18779 11115 18785
rect 11146 18776 11152 18828
rect 11204 18816 11210 18828
rect 14918 18816 14924 18828
rect 11204 18788 14924 18816
rect 11204 18776 11210 18788
rect 14918 18776 14924 18788
rect 14976 18776 14982 18828
rect 17678 18816 17684 18828
rect 16040 18788 17684 18816
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18748 1639 18751
rect 1946 18748 1952 18760
rect 1627 18720 1952 18748
rect 1627 18717 1639 18720
rect 1581 18711 1639 18717
rect 1946 18708 1952 18720
rect 2004 18708 2010 18760
rect 10965 18751 11023 18757
rect 10965 18717 10977 18751
rect 11011 18717 11023 18751
rect 10965 18711 11023 18717
rect 1854 18680 1860 18692
rect 1815 18652 1860 18680
rect 1854 18640 1860 18652
rect 1912 18640 1918 18692
rect 10980 18612 11008 18711
rect 11238 18708 11244 18760
rect 11296 18748 11302 18760
rect 16040 18757 16068 18788
rect 17678 18776 17684 18788
rect 17736 18816 17742 18828
rect 17736 18788 18460 18816
rect 17736 18776 17742 18788
rect 16206 18757 16212 18760
rect 16025 18751 16083 18757
rect 11296 18720 11341 18748
rect 11296 18708 11302 18720
rect 16025 18717 16037 18751
rect 16071 18717 16083 18751
rect 16025 18711 16083 18717
rect 16179 18751 16212 18757
rect 16179 18717 16191 18751
rect 16179 18711 16212 18717
rect 16206 18708 16212 18711
rect 16264 18708 16270 18760
rect 16945 18751 17003 18757
rect 16945 18717 16957 18751
rect 16991 18748 17003 18751
rect 17126 18748 17132 18760
rect 16991 18720 17132 18748
rect 16991 18717 17003 18720
rect 16945 18711 17003 18717
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 17313 18751 17371 18757
rect 17313 18748 17325 18751
rect 17236 18720 17325 18748
rect 15838 18640 15844 18692
rect 15896 18680 15902 18692
rect 16393 18683 16451 18689
rect 16393 18680 16405 18683
rect 15896 18652 16405 18680
rect 15896 18640 15902 18652
rect 16393 18649 16405 18652
rect 16439 18680 16451 18683
rect 17236 18680 17264 18720
rect 17313 18717 17325 18720
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17494 18708 17500 18760
rect 17552 18748 17558 18760
rect 17552 18720 17597 18748
rect 17552 18708 17558 18720
rect 16439 18652 17264 18680
rect 18432 18680 18460 18788
rect 18524 18757 18552 18924
rect 18598 18776 18604 18828
rect 18656 18816 18662 18828
rect 18877 18819 18935 18825
rect 18656 18788 18701 18816
rect 18656 18776 18662 18788
rect 18877 18785 18889 18819
rect 18923 18785 18935 18819
rect 18877 18779 18935 18785
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18717 18567 18751
rect 18892 18748 18920 18779
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 19794 18816 19800 18828
rect 19484 18788 19800 18816
rect 19484 18776 19490 18788
rect 19794 18776 19800 18788
rect 19852 18776 19858 18828
rect 20824 18816 20852 18924
rect 22066 18924 25136 18952
rect 20898 18844 20904 18896
rect 20956 18884 20962 18896
rect 22066 18884 22094 18924
rect 25130 18912 25136 18924
rect 25188 18912 25194 18964
rect 25682 18912 25688 18964
rect 25740 18952 25746 18964
rect 28626 18952 28632 18964
rect 25740 18924 28632 18952
rect 25740 18912 25746 18924
rect 28626 18912 28632 18924
rect 28684 18912 28690 18964
rect 28810 18912 28816 18964
rect 28868 18952 28874 18964
rect 34698 18952 34704 18964
rect 28868 18924 34704 18952
rect 28868 18912 28874 18924
rect 34698 18912 34704 18924
rect 34756 18912 34762 18964
rect 35342 18912 35348 18964
rect 35400 18952 35406 18964
rect 35437 18955 35495 18961
rect 35437 18952 35449 18955
rect 35400 18924 35449 18952
rect 35400 18912 35406 18924
rect 35437 18921 35449 18924
rect 35483 18921 35495 18955
rect 35894 18952 35900 18964
rect 35437 18915 35495 18921
rect 35544 18924 35900 18952
rect 20956 18856 22094 18884
rect 20956 18844 20962 18856
rect 22554 18844 22560 18896
rect 22612 18884 22618 18896
rect 30834 18884 30840 18896
rect 22612 18856 28769 18884
rect 22612 18844 22618 18856
rect 27338 18816 27344 18828
rect 20824 18788 23428 18816
rect 21729 18751 21787 18757
rect 21729 18748 21741 18751
rect 18892 18720 21741 18748
rect 18509 18711 18567 18717
rect 21729 18717 21741 18720
rect 21775 18717 21787 18751
rect 21729 18711 21787 18717
rect 19426 18680 19432 18692
rect 18432 18652 19432 18680
rect 16439 18649 16451 18652
rect 16393 18643 16451 18649
rect 19426 18640 19432 18652
rect 19484 18640 19490 18692
rect 20064 18683 20122 18689
rect 20064 18649 20076 18683
rect 20110 18680 20122 18683
rect 20346 18680 20352 18692
rect 20110 18652 20352 18680
rect 20110 18649 20122 18652
rect 20064 18643 20122 18649
rect 20346 18640 20352 18652
rect 20404 18640 20410 18692
rect 23400 18680 23428 18788
rect 24596 18788 27344 18816
rect 23658 18708 23664 18760
rect 23716 18748 23722 18760
rect 24596 18757 24624 18788
rect 27338 18776 27344 18788
rect 27396 18776 27402 18828
rect 28074 18776 28080 18828
rect 28132 18816 28138 18828
rect 28534 18816 28540 18828
rect 28132 18788 28304 18816
rect 28132 18776 28138 18788
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 23716 18720 24593 18748
rect 23716 18708 23722 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18717 24823 18751
rect 24765 18711 24823 18717
rect 25225 18751 25283 18757
rect 25225 18717 25237 18751
rect 25271 18748 25283 18751
rect 27154 18748 27160 18760
rect 25271 18720 27160 18748
rect 25271 18717 25283 18720
rect 25225 18711 25283 18717
rect 24780 18680 24808 18711
rect 27154 18708 27160 18720
rect 27212 18708 27218 18760
rect 28276 18757 28304 18788
rect 28368 18788 28540 18816
rect 28368 18757 28396 18788
rect 28534 18776 28540 18788
rect 28592 18776 28598 18828
rect 28741 18816 28769 18856
rect 28966 18856 30840 18884
rect 28966 18816 28994 18856
rect 30834 18844 30840 18856
rect 30892 18844 30898 18896
rect 33594 18884 33600 18896
rect 32508 18856 33600 18884
rect 28741 18788 28994 18816
rect 30466 18776 30472 18828
rect 30524 18816 30530 18828
rect 30524 18788 30696 18816
rect 30524 18776 30530 18788
rect 28261 18751 28319 18757
rect 28261 18717 28273 18751
rect 28307 18717 28319 18751
rect 28261 18711 28319 18717
rect 28353 18751 28411 18757
rect 28353 18717 28365 18751
rect 28399 18717 28411 18751
rect 28353 18711 28411 18717
rect 28445 18751 28503 18757
rect 28445 18717 28457 18751
rect 28491 18748 28503 18751
rect 28629 18751 28687 18757
rect 28491 18720 28580 18748
rect 28491 18717 28503 18720
rect 28445 18711 28503 18717
rect 27522 18680 27528 18692
rect 23400 18652 27528 18680
rect 27522 18640 27528 18652
rect 27580 18640 27586 18692
rect 28552 18680 28580 18720
rect 28629 18717 28641 18751
rect 28675 18748 28687 18751
rect 30374 18748 30380 18760
rect 28675 18720 30380 18748
rect 28675 18717 28687 18720
rect 28629 18711 28687 18717
rect 30374 18708 30380 18720
rect 30432 18708 30438 18760
rect 30558 18748 30564 18760
rect 30519 18720 30564 18748
rect 30558 18708 30564 18720
rect 30616 18708 30622 18760
rect 30668 18748 30696 18788
rect 30742 18776 30748 18828
rect 30800 18816 30806 18828
rect 30800 18788 30845 18816
rect 30800 18776 30806 18788
rect 30837 18751 30895 18757
rect 30837 18748 30849 18751
rect 30668 18720 30849 18748
rect 30837 18717 30849 18720
rect 30883 18717 30895 18751
rect 30837 18711 30895 18717
rect 31018 18708 31024 18760
rect 31076 18748 31082 18760
rect 31113 18751 31171 18757
rect 31113 18748 31125 18751
rect 31076 18720 31125 18748
rect 31076 18708 31082 18720
rect 31113 18717 31125 18720
rect 31159 18717 31171 18751
rect 31570 18748 31576 18760
rect 31531 18720 31576 18748
rect 31113 18711 31171 18717
rect 31570 18708 31576 18720
rect 31628 18708 31634 18760
rect 32508 18757 32536 18856
rect 33594 18844 33600 18856
rect 33652 18844 33658 18896
rect 34882 18844 34888 18896
rect 34940 18884 34946 18896
rect 35544 18884 35572 18924
rect 35894 18912 35900 18924
rect 35952 18912 35958 18964
rect 37458 18952 37464 18964
rect 36188 18924 37464 18952
rect 36078 18884 36084 18896
rect 34940 18856 35572 18884
rect 35820 18856 36084 18884
rect 34940 18844 34946 18856
rect 32784 18788 33916 18816
rect 32784 18760 32812 18788
rect 33888 18760 33916 18788
rect 32493 18751 32551 18757
rect 32493 18717 32505 18751
rect 32539 18717 32551 18751
rect 32493 18711 32551 18717
rect 32585 18751 32643 18757
rect 32585 18717 32597 18751
rect 32631 18717 32643 18751
rect 32766 18748 32772 18760
rect 32727 18720 32772 18748
rect 32585 18711 32643 18717
rect 30006 18680 30012 18692
rect 28552 18652 30012 18680
rect 30006 18640 30012 18652
rect 30064 18640 30070 18692
rect 32214 18640 32220 18692
rect 32272 18680 32278 18692
rect 32600 18680 32628 18711
rect 32766 18708 32772 18720
rect 32824 18708 32830 18760
rect 32858 18708 32864 18760
rect 32916 18748 32922 18760
rect 33410 18748 33416 18760
rect 32916 18720 32961 18748
rect 33371 18720 33416 18748
rect 32916 18708 32922 18720
rect 33410 18708 33416 18720
rect 33468 18708 33474 18760
rect 33594 18748 33600 18760
rect 33555 18720 33600 18748
rect 33594 18708 33600 18720
rect 33652 18708 33658 18760
rect 33688 18751 33746 18757
rect 33688 18717 33700 18751
rect 33734 18717 33746 18751
rect 33870 18748 33876 18760
rect 33783 18720 33876 18748
rect 33688 18711 33746 18717
rect 32272 18652 32628 18680
rect 32272 18640 32278 18652
rect 33704 18624 33732 18711
rect 33870 18708 33876 18720
rect 33928 18708 33934 18760
rect 33965 18751 34023 18757
rect 33965 18717 33977 18751
rect 34011 18748 34023 18751
rect 35250 18748 35256 18760
rect 34011 18720 35256 18748
rect 34011 18717 34023 18720
rect 33965 18711 34023 18717
rect 35250 18708 35256 18720
rect 35308 18708 35314 18760
rect 35342 18708 35348 18760
rect 35400 18748 35406 18760
rect 35820 18757 35848 18856
rect 36078 18844 36084 18856
rect 36136 18844 36142 18896
rect 36188 18816 36216 18924
rect 37458 18912 37464 18924
rect 37516 18912 37522 18964
rect 37550 18912 37556 18964
rect 37608 18952 37614 18964
rect 37921 18955 37979 18961
rect 37921 18952 37933 18955
rect 37608 18924 37933 18952
rect 37608 18912 37614 18924
rect 37921 18921 37933 18924
rect 37967 18921 37979 18955
rect 38378 18952 38384 18964
rect 38339 18924 38384 18952
rect 37921 18915 37979 18921
rect 38378 18912 38384 18924
rect 38436 18912 38442 18964
rect 46198 18952 46204 18964
rect 38488 18924 46204 18952
rect 37734 18844 37740 18896
rect 37792 18884 37798 18896
rect 38488 18884 38516 18924
rect 46198 18912 46204 18924
rect 46256 18912 46262 18964
rect 57146 18912 57152 18964
rect 57204 18952 57210 18964
rect 57882 18952 57888 18964
rect 57204 18924 57888 18952
rect 57204 18912 57210 18924
rect 57882 18912 57888 18924
rect 57940 18952 57946 18964
rect 58253 18955 58311 18961
rect 58253 18952 58265 18955
rect 57940 18924 58265 18952
rect 57940 18912 57946 18924
rect 58253 18921 58265 18924
rect 58299 18921 58311 18955
rect 58253 18915 58311 18921
rect 37792 18856 38516 18884
rect 38580 18856 38700 18884
rect 37792 18844 37798 18856
rect 36096 18788 36216 18816
rect 36096 18760 36124 18788
rect 38010 18776 38016 18828
rect 38068 18816 38074 18828
rect 38580 18816 38608 18856
rect 38068 18788 38608 18816
rect 38672 18816 38700 18856
rect 38746 18844 38752 18896
rect 38804 18884 38810 18896
rect 43990 18884 43996 18896
rect 38804 18856 39068 18884
rect 38804 18844 38810 18856
rect 38672 18788 38792 18816
rect 38068 18776 38074 18788
rect 35713 18751 35771 18757
rect 35400 18745 35664 18748
rect 35713 18745 35725 18751
rect 35400 18720 35725 18745
rect 35400 18708 35406 18720
rect 35636 18717 35725 18720
rect 35759 18717 35771 18751
rect 35713 18711 35771 18717
rect 35805 18751 35863 18757
rect 35805 18717 35817 18751
rect 35851 18717 35863 18751
rect 35805 18711 35863 18717
rect 35897 18751 35955 18757
rect 35897 18717 35909 18751
rect 35943 18717 35955 18751
rect 35897 18711 35955 18717
rect 33778 18640 33784 18692
rect 33836 18680 33842 18692
rect 33836 18652 35756 18680
rect 33836 18640 33842 18652
rect 16850 18612 16856 18624
rect 10980 18584 16856 18612
rect 16850 18572 16856 18584
rect 16908 18572 16914 18624
rect 17034 18612 17040 18624
rect 16995 18584 17040 18612
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 17218 18572 17224 18624
rect 17276 18612 17282 18624
rect 21082 18612 21088 18624
rect 17276 18584 21088 18612
rect 17276 18572 17282 18584
rect 21082 18572 21088 18584
rect 21140 18572 21146 18624
rect 21177 18615 21235 18621
rect 21177 18581 21189 18615
rect 21223 18612 21235 18615
rect 22554 18612 22560 18624
rect 21223 18584 22560 18612
rect 21223 18581 21235 18584
rect 21177 18575 21235 18581
rect 22554 18572 22560 18584
rect 22612 18572 22618 18624
rect 22922 18612 22928 18624
rect 22883 18584 22928 18612
rect 22922 18572 22928 18584
rect 22980 18572 22986 18624
rect 24765 18615 24823 18621
rect 24765 18581 24777 18615
rect 24811 18612 24823 18615
rect 25314 18612 25320 18624
rect 24811 18584 25320 18612
rect 24811 18581 24823 18584
rect 24765 18575 24823 18581
rect 25314 18572 25320 18584
rect 25372 18572 25378 18624
rect 25406 18572 25412 18624
rect 25464 18612 25470 18624
rect 26421 18615 26479 18621
rect 26421 18612 26433 18615
rect 25464 18584 26433 18612
rect 25464 18572 25470 18584
rect 26421 18581 26433 18584
rect 26467 18581 26479 18615
rect 26421 18575 26479 18581
rect 27985 18615 28043 18621
rect 27985 18581 27997 18615
rect 28031 18612 28043 18615
rect 28074 18612 28080 18624
rect 28031 18584 28080 18612
rect 28031 18581 28043 18584
rect 27985 18575 28043 18581
rect 28074 18572 28080 18584
rect 28132 18572 28138 18624
rect 28258 18572 28264 18624
rect 28316 18612 28322 18624
rect 31294 18612 31300 18624
rect 28316 18584 31300 18612
rect 28316 18572 28322 18584
rect 31294 18572 31300 18584
rect 31352 18572 31358 18624
rect 31570 18572 31576 18624
rect 31628 18612 31634 18624
rect 32309 18615 32367 18621
rect 32309 18612 32321 18615
rect 31628 18584 32321 18612
rect 31628 18572 31634 18584
rect 32309 18581 32321 18584
rect 32355 18581 32367 18615
rect 32309 18575 32367 18581
rect 33686 18572 33692 18624
rect 33744 18572 33750 18624
rect 35728 18612 35756 18652
rect 35912 18612 35940 18711
rect 36078 18708 36084 18760
rect 36136 18748 36142 18760
rect 36538 18748 36544 18760
rect 36136 18720 36181 18748
rect 36451 18720 36544 18748
rect 36136 18708 36142 18720
rect 36538 18708 36544 18720
rect 36596 18748 36602 18760
rect 37642 18748 37648 18760
rect 36596 18720 37648 18748
rect 36596 18708 36602 18720
rect 37642 18708 37648 18720
rect 37700 18708 37706 18760
rect 38562 18708 38568 18760
rect 38620 18748 38626 18760
rect 38764 18757 38792 18788
rect 39040 18760 39068 18856
rect 41386 18856 43996 18884
rect 41046 18776 41052 18828
rect 41104 18816 41110 18828
rect 41386 18816 41414 18856
rect 43990 18844 43996 18856
rect 44048 18844 44054 18896
rect 44358 18884 44364 18896
rect 44319 18856 44364 18884
rect 44358 18844 44364 18856
rect 44416 18844 44422 18896
rect 41104 18788 41414 18816
rect 43073 18819 43131 18825
rect 41104 18776 41110 18788
rect 43073 18785 43085 18819
rect 43119 18816 43131 18819
rect 44266 18816 44272 18828
rect 43119 18788 44272 18816
rect 43119 18785 43131 18788
rect 43073 18779 43131 18785
rect 44266 18776 44272 18788
rect 44324 18776 44330 18828
rect 45370 18816 45376 18828
rect 44376 18788 45376 18816
rect 38657 18751 38715 18757
rect 38657 18748 38669 18751
rect 38620 18720 38669 18748
rect 38620 18708 38626 18720
rect 38657 18717 38669 18720
rect 38703 18717 38715 18751
rect 38657 18711 38715 18717
rect 38746 18751 38804 18757
rect 38746 18717 38758 18751
rect 38792 18717 38804 18751
rect 38746 18711 38804 18717
rect 38862 18745 38920 18751
rect 38862 18711 38874 18745
rect 38908 18742 38920 18745
rect 38908 18714 38976 18742
rect 38908 18711 38920 18714
rect 38862 18705 38920 18711
rect 36262 18640 36268 18692
rect 36320 18680 36326 18692
rect 36786 18683 36844 18689
rect 36786 18680 36798 18683
rect 36320 18652 36798 18680
rect 36320 18640 36326 18652
rect 36786 18649 36798 18652
rect 36832 18649 36844 18683
rect 38948 18680 38976 18714
rect 39022 18708 39028 18760
rect 39080 18748 39086 18760
rect 42981 18751 43039 18757
rect 39080 18720 39173 18748
rect 39080 18708 39086 18720
rect 42981 18717 42993 18751
rect 43027 18717 43039 18751
rect 43162 18748 43168 18760
rect 43123 18720 43168 18748
rect 42981 18711 43039 18717
rect 39206 18680 39212 18692
rect 38948 18652 39212 18680
rect 36786 18643 36844 18649
rect 39206 18640 39212 18652
rect 39264 18640 39270 18692
rect 42996 18680 43024 18711
rect 43162 18708 43168 18720
rect 43220 18708 43226 18760
rect 43990 18751 44048 18757
rect 43990 18717 44002 18751
rect 44036 18748 44048 18751
rect 44376 18748 44404 18788
rect 45370 18776 45376 18788
rect 45428 18776 45434 18828
rect 44036 18720 44404 18748
rect 44036 18717 44048 18720
rect 43990 18711 44048 18717
rect 44450 18708 44456 18760
rect 44508 18748 44514 18760
rect 56870 18748 56876 18760
rect 44508 18720 44553 18748
rect 56831 18720 56876 18748
rect 44508 18708 44514 18720
rect 56870 18708 56876 18720
rect 56928 18708 56934 18760
rect 56962 18708 56968 18760
rect 57020 18748 57026 18760
rect 57129 18751 57187 18757
rect 57129 18748 57141 18751
rect 57020 18720 57141 18748
rect 57020 18708 57026 18720
rect 57129 18717 57141 18720
rect 57175 18717 57187 18751
rect 57129 18711 57187 18717
rect 42996 18652 43852 18680
rect 35728 18584 35940 18612
rect 38378 18572 38384 18624
rect 38436 18612 38442 18624
rect 41874 18612 41880 18624
rect 38436 18584 41880 18612
rect 38436 18572 38442 18584
rect 41874 18572 41880 18584
rect 41932 18612 41938 18624
rect 42426 18612 42432 18624
rect 41932 18584 42432 18612
rect 41932 18572 41938 18584
rect 42426 18572 42432 18584
rect 42484 18572 42490 18624
rect 43438 18612 43444 18624
rect 43399 18584 43444 18612
rect 43438 18572 43444 18584
rect 43496 18572 43502 18624
rect 43824 18621 43852 18652
rect 43898 18640 43904 18692
rect 43956 18680 43962 18692
rect 43956 18652 51074 18680
rect 43956 18640 43962 18652
rect 43809 18615 43867 18621
rect 43809 18581 43821 18615
rect 43855 18581 43867 18615
rect 43990 18612 43996 18624
rect 43951 18584 43996 18612
rect 43809 18575 43867 18581
rect 43990 18572 43996 18584
rect 44048 18572 44054 18624
rect 51046 18612 51074 18652
rect 59170 18612 59176 18624
rect 51046 18584 59176 18612
rect 59170 18572 59176 18584
rect 59228 18572 59234 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 10505 18411 10563 18417
rect 10505 18377 10517 18411
rect 10551 18408 10563 18411
rect 11238 18408 11244 18420
rect 10551 18380 11244 18408
rect 10551 18377 10563 18380
rect 10505 18371 10563 18377
rect 11238 18368 11244 18380
rect 11296 18368 11302 18420
rect 13078 18368 13084 18420
rect 13136 18408 13142 18420
rect 16209 18411 16267 18417
rect 16209 18408 16221 18411
rect 13136 18380 16221 18408
rect 13136 18368 13142 18380
rect 16209 18377 16221 18380
rect 16255 18377 16267 18411
rect 16209 18371 16267 18377
rect 16850 18368 16856 18420
rect 16908 18408 16914 18420
rect 18690 18408 18696 18420
rect 16908 18380 18696 18408
rect 16908 18368 16914 18380
rect 18690 18368 18696 18380
rect 18748 18408 18754 18420
rect 19242 18408 19248 18420
rect 18748 18380 19248 18408
rect 18748 18368 18754 18380
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 19978 18368 19984 18420
rect 20036 18408 20042 18420
rect 20346 18408 20352 18420
rect 20036 18380 20208 18408
rect 20307 18380 20352 18408
rect 20036 18368 20042 18380
rect 10045 18343 10103 18349
rect 10045 18309 10057 18343
rect 10091 18340 10103 18343
rect 11146 18340 11152 18352
rect 10091 18312 11152 18340
rect 10091 18309 10103 18312
rect 10045 18303 10103 18309
rect 11146 18300 11152 18312
rect 11204 18300 11210 18352
rect 16114 18300 16120 18352
rect 16172 18340 16178 18352
rect 16172 18312 17448 18340
rect 16172 18300 16178 18312
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18272 1639 18275
rect 1627 18244 12434 18272
rect 1627 18241 1639 18244
rect 1581 18235 1639 18241
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 12406 18204 12434 18244
rect 14918 18232 14924 18284
rect 14976 18272 14982 18284
rect 15197 18275 15255 18281
rect 15197 18272 15209 18275
rect 14976 18244 15209 18272
rect 14976 18232 14982 18244
rect 15197 18241 15209 18244
rect 15243 18241 15255 18275
rect 15838 18272 15844 18284
rect 15799 18244 15844 18272
rect 15197 18235 15255 18241
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 17126 18272 17132 18284
rect 17087 18244 17132 18272
rect 17126 18232 17132 18244
rect 17184 18232 17190 18284
rect 17221 18275 17279 18281
rect 17221 18241 17233 18275
rect 17267 18272 17279 18275
rect 17310 18272 17316 18284
rect 17267 18244 17316 18272
rect 17267 18241 17279 18244
rect 17221 18235 17279 18241
rect 17310 18232 17316 18244
rect 17368 18232 17374 18284
rect 17420 18281 17448 18312
rect 17494 18300 17500 18352
rect 17552 18340 17558 18352
rect 20070 18340 20076 18352
rect 17552 18312 20076 18340
rect 17552 18300 17558 18312
rect 17405 18275 17463 18281
rect 17405 18241 17417 18275
rect 17451 18241 17463 18275
rect 18046 18272 18052 18284
rect 17405 18235 17463 18241
rect 17512 18244 18052 18272
rect 14829 18207 14887 18213
rect 14829 18204 14841 18207
rect 12406 18176 14841 18204
rect 14829 18173 14841 18176
rect 14875 18173 14887 18207
rect 14829 18167 14887 18173
rect 15013 18207 15071 18213
rect 15013 18173 15025 18207
rect 15059 18173 15071 18207
rect 15013 18167 15071 18173
rect 15105 18207 15163 18213
rect 15105 18173 15117 18207
rect 15151 18173 15163 18207
rect 15105 18167 15163 18173
rect 7558 18096 7564 18148
rect 7616 18136 7622 18148
rect 10321 18139 10379 18145
rect 10321 18136 10333 18139
rect 7616 18108 10333 18136
rect 7616 18096 7622 18108
rect 10321 18105 10333 18108
rect 10367 18105 10379 18139
rect 10321 18099 10379 18105
rect 14734 18096 14740 18148
rect 14792 18136 14798 18148
rect 15028 18136 15056 18167
rect 14792 18108 15056 18136
rect 15120 18136 15148 18167
rect 15286 18164 15292 18216
rect 15344 18204 15350 18216
rect 15344 18176 15389 18204
rect 15344 18164 15350 18176
rect 15562 18164 15568 18216
rect 15620 18204 15626 18216
rect 15933 18207 15991 18213
rect 15933 18204 15945 18207
rect 15620 18176 15945 18204
rect 15620 18164 15626 18176
rect 15933 18173 15945 18176
rect 15979 18173 15991 18207
rect 15933 18167 15991 18173
rect 16942 18164 16948 18216
rect 17000 18204 17006 18216
rect 17512 18204 17540 18244
rect 18046 18232 18052 18244
rect 18104 18272 18110 18284
rect 18616 18281 18644 18312
rect 20070 18300 20076 18312
rect 20128 18300 20134 18352
rect 20180 18340 20208 18380
rect 20346 18368 20352 18380
rect 20404 18368 20410 18420
rect 22462 18368 22468 18420
rect 22520 18408 22526 18420
rect 25501 18411 25559 18417
rect 25501 18408 25513 18411
rect 22520 18380 25513 18408
rect 22520 18368 22526 18380
rect 25501 18377 25513 18380
rect 25547 18377 25559 18411
rect 25501 18371 25559 18377
rect 27430 18368 27436 18420
rect 27488 18408 27494 18420
rect 29730 18408 29736 18420
rect 27488 18380 29736 18408
rect 27488 18368 27494 18380
rect 29730 18368 29736 18380
rect 29788 18408 29794 18420
rect 32769 18411 32827 18417
rect 29788 18380 30880 18408
rect 29788 18368 29794 18380
rect 22094 18340 22100 18352
rect 20180 18312 22100 18340
rect 22094 18300 22100 18312
rect 22152 18340 22158 18352
rect 22640 18343 22698 18349
rect 22152 18312 22416 18340
rect 22152 18300 22158 18312
rect 18325 18275 18383 18281
rect 18325 18272 18337 18275
rect 18104 18244 18337 18272
rect 18104 18232 18110 18244
rect 18325 18241 18337 18244
rect 18371 18241 18383 18275
rect 18325 18235 18383 18241
rect 18601 18275 18659 18281
rect 18601 18241 18613 18275
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 19153 18275 19211 18281
rect 19153 18241 19165 18275
rect 19199 18272 19211 18275
rect 20990 18272 20996 18284
rect 19199 18244 20996 18272
rect 19199 18241 19211 18244
rect 19153 18235 19211 18241
rect 20990 18232 20996 18244
rect 21048 18232 21054 18284
rect 22388 18281 22416 18312
rect 22640 18309 22652 18343
rect 22686 18340 22698 18343
rect 22922 18340 22928 18352
rect 22686 18312 22928 18340
rect 22686 18309 22698 18312
rect 22640 18303 22698 18309
rect 22922 18300 22928 18312
rect 22980 18300 22986 18352
rect 25130 18300 25136 18352
rect 25188 18340 25194 18352
rect 27706 18340 27712 18352
rect 25188 18312 27712 18340
rect 25188 18300 25194 18312
rect 27706 18300 27712 18312
rect 27764 18300 27770 18352
rect 28902 18340 28908 18352
rect 27816 18312 28908 18340
rect 22373 18275 22431 18281
rect 22373 18241 22385 18275
rect 22419 18272 22431 18275
rect 22462 18272 22468 18284
rect 22419 18244 22468 18272
rect 22419 18241 22431 18244
rect 22373 18235 22431 18241
rect 22462 18232 22468 18244
rect 22520 18232 22526 18284
rect 24305 18275 24363 18281
rect 24305 18241 24317 18275
rect 24351 18272 24363 18275
rect 25774 18272 25780 18284
rect 24351 18244 25780 18272
rect 24351 18241 24363 18244
rect 24305 18235 24363 18241
rect 25774 18232 25780 18244
rect 25832 18232 25838 18284
rect 26326 18232 26332 18284
rect 26384 18272 26390 18284
rect 26970 18272 26976 18284
rect 26384 18244 26976 18272
rect 26384 18232 26390 18244
rect 26970 18232 26976 18244
rect 27028 18232 27034 18284
rect 27154 18272 27160 18284
rect 27115 18244 27160 18272
rect 27154 18232 27160 18244
rect 27212 18232 27218 18284
rect 27816 18281 27844 18312
rect 28902 18300 28908 18312
rect 28960 18300 28966 18352
rect 28074 18281 28080 18284
rect 27341 18275 27399 18281
rect 27341 18241 27353 18275
rect 27387 18241 27399 18275
rect 27341 18235 27399 18241
rect 27801 18275 27859 18281
rect 27801 18241 27813 18275
rect 27847 18241 27859 18275
rect 28068 18272 28080 18281
rect 28035 18244 28080 18272
rect 27801 18235 27859 18241
rect 28068 18235 28080 18244
rect 17000 18176 17540 18204
rect 17865 18207 17923 18213
rect 17000 18164 17006 18176
rect 17865 18173 17877 18207
rect 17911 18204 17923 18207
rect 20438 18204 20444 18216
rect 17911 18176 20444 18204
rect 17911 18173 17923 18176
rect 17865 18167 17923 18173
rect 20438 18164 20444 18176
rect 20496 18164 20502 18216
rect 20622 18164 20628 18216
rect 20680 18164 20686 18216
rect 25038 18164 25044 18216
rect 25096 18204 25102 18216
rect 27356 18204 27384 18235
rect 28074 18232 28080 18235
rect 28132 18232 28138 18284
rect 28810 18232 28816 18284
rect 28868 18272 28874 18284
rect 30374 18272 30380 18284
rect 28868 18244 30380 18272
rect 28868 18232 28874 18244
rect 30374 18232 30380 18244
rect 30432 18232 30438 18284
rect 30852 18281 30880 18380
rect 32769 18377 32781 18411
rect 32815 18408 32827 18411
rect 33778 18408 33784 18420
rect 32815 18380 33784 18408
rect 32815 18377 32827 18380
rect 32769 18371 32827 18377
rect 33778 18368 33784 18380
rect 33836 18368 33842 18420
rect 35342 18368 35348 18420
rect 35400 18408 35406 18420
rect 35802 18408 35808 18420
rect 35400 18380 35808 18408
rect 35400 18368 35406 18380
rect 35802 18368 35808 18380
rect 35860 18408 35866 18420
rect 37734 18408 37740 18420
rect 35860 18380 37740 18408
rect 35860 18368 35866 18380
rect 37734 18368 37740 18380
rect 37792 18368 37798 18420
rect 37921 18411 37979 18417
rect 37921 18377 37933 18411
rect 37967 18408 37979 18411
rect 52454 18408 52460 18420
rect 37967 18380 52460 18408
rect 37967 18377 37979 18380
rect 37921 18371 37979 18377
rect 52454 18368 52460 18380
rect 52512 18368 52518 18420
rect 56778 18368 56784 18420
rect 56836 18408 56842 18420
rect 56965 18411 57023 18417
rect 56965 18408 56977 18411
rect 56836 18380 56977 18408
rect 56836 18368 56842 18380
rect 56965 18377 56977 18380
rect 57011 18377 57023 18411
rect 56965 18371 57023 18377
rect 58066 18368 58072 18420
rect 58124 18408 58130 18420
rect 58161 18411 58219 18417
rect 58161 18408 58173 18411
rect 58124 18380 58173 18408
rect 58124 18368 58130 18380
rect 58161 18377 58173 18380
rect 58207 18377 58219 18411
rect 58161 18371 58219 18377
rect 31018 18300 31024 18352
rect 31076 18340 31082 18352
rect 31662 18340 31668 18352
rect 31076 18312 31668 18340
rect 31076 18300 31082 18312
rect 30837 18275 30895 18281
rect 30837 18241 30849 18275
rect 30883 18241 30895 18275
rect 31110 18272 31116 18284
rect 31071 18244 31116 18272
rect 30837 18235 30895 18241
rect 31110 18232 31116 18244
rect 31168 18232 31174 18284
rect 31496 18281 31524 18312
rect 31662 18300 31668 18312
rect 31720 18300 31726 18352
rect 31754 18300 31760 18352
rect 31812 18340 31818 18352
rect 32306 18340 32312 18352
rect 31812 18312 32312 18340
rect 31812 18300 31818 18312
rect 32306 18300 32312 18312
rect 32364 18340 32370 18352
rect 32401 18343 32459 18349
rect 32401 18340 32413 18343
rect 32364 18312 32413 18340
rect 32364 18300 32370 18312
rect 32401 18309 32413 18312
rect 32447 18309 32459 18343
rect 32582 18340 32588 18352
rect 32543 18312 32588 18340
rect 32401 18303 32459 18309
rect 32582 18300 32588 18312
rect 32640 18300 32646 18352
rect 34238 18340 34244 18352
rect 33612 18312 34244 18340
rect 31481 18275 31539 18281
rect 31481 18241 31493 18275
rect 31527 18241 31539 18275
rect 33134 18272 33140 18284
rect 31481 18235 31539 18241
rect 31726 18244 33140 18272
rect 25096 18176 27384 18204
rect 25096 18164 25102 18176
rect 28994 18164 29000 18216
rect 29052 18204 29058 18216
rect 30650 18204 30656 18216
rect 29052 18176 30656 18204
rect 29052 18164 29058 18176
rect 30650 18164 30656 18176
rect 30708 18164 30714 18216
rect 30742 18164 30748 18216
rect 30800 18204 30806 18216
rect 30800 18176 30845 18204
rect 30800 18164 30806 18176
rect 20640 18136 20668 18164
rect 15120 18108 20668 18136
rect 14792 18096 14798 18108
rect 23382 18096 23388 18148
rect 23440 18136 23446 18148
rect 31726 18136 31754 18244
rect 33134 18232 33140 18244
rect 33192 18232 33198 18284
rect 33502 18272 33508 18284
rect 33463 18244 33508 18272
rect 33502 18232 33508 18244
rect 33560 18232 33566 18284
rect 33612 18281 33640 18312
rect 34238 18300 34244 18312
rect 34296 18300 34302 18352
rect 34514 18300 34520 18352
rect 34572 18340 34578 18352
rect 34609 18343 34667 18349
rect 34609 18340 34621 18343
rect 34572 18312 34621 18340
rect 34572 18300 34578 18312
rect 34609 18309 34621 18312
rect 34655 18340 34667 18343
rect 35618 18340 35624 18352
rect 34655 18312 35624 18340
rect 34655 18309 34667 18312
rect 34609 18303 34667 18309
rect 35618 18300 35624 18312
rect 35676 18300 35682 18352
rect 39206 18340 39212 18352
rect 39167 18312 39212 18340
rect 39206 18300 39212 18312
rect 39264 18300 39270 18352
rect 41230 18340 41236 18352
rect 39776 18312 41236 18340
rect 33597 18275 33655 18281
rect 33597 18241 33609 18275
rect 33643 18241 33655 18275
rect 33781 18275 33839 18281
rect 33781 18272 33793 18275
rect 33597 18235 33655 18241
rect 33704 18244 33793 18272
rect 33704 18204 33732 18244
rect 33781 18241 33793 18244
rect 33827 18241 33839 18275
rect 33781 18235 33839 18241
rect 33870 18232 33876 18284
rect 33928 18272 33934 18284
rect 34333 18275 34391 18281
rect 34333 18272 34345 18275
rect 33928 18244 33973 18272
rect 34256 18244 34345 18272
rect 33928 18232 33934 18244
rect 33962 18204 33968 18216
rect 33704 18176 33968 18204
rect 33962 18164 33968 18176
rect 34020 18204 34026 18216
rect 34256 18204 34284 18244
rect 34333 18241 34345 18244
rect 34379 18241 34391 18275
rect 34333 18235 34391 18241
rect 34422 18232 34428 18284
rect 34480 18272 34486 18284
rect 34480 18244 34525 18272
rect 34480 18232 34486 18244
rect 34698 18232 34704 18284
rect 34756 18272 34762 18284
rect 34882 18281 34888 18284
rect 34839 18275 34888 18281
rect 34756 18244 34801 18272
rect 34756 18232 34762 18244
rect 34839 18241 34851 18275
rect 34885 18241 34888 18275
rect 34839 18235 34888 18241
rect 34882 18232 34888 18235
rect 34940 18232 34946 18284
rect 35342 18232 35348 18284
rect 35400 18272 35406 18284
rect 37737 18275 37795 18281
rect 37737 18272 37749 18275
rect 35400 18244 37749 18272
rect 35400 18232 35406 18244
rect 37737 18241 37749 18244
rect 37783 18241 37795 18275
rect 38102 18272 38108 18284
rect 38063 18244 38108 18272
rect 37737 18235 37795 18241
rect 38102 18232 38108 18244
rect 38160 18232 38166 18284
rect 38378 18272 38384 18284
rect 38339 18244 38384 18272
rect 38378 18232 38384 18244
rect 38436 18232 38442 18284
rect 38838 18272 38844 18284
rect 38799 18244 38844 18272
rect 38838 18232 38844 18244
rect 38896 18232 38902 18284
rect 39025 18275 39083 18281
rect 39025 18241 39037 18275
rect 39071 18272 39083 18275
rect 39666 18272 39672 18284
rect 39071 18244 39672 18272
rect 39071 18241 39083 18244
rect 39025 18235 39083 18241
rect 39666 18232 39672 18244
rect 39724 18232 39730 18284
rect 39776 18281 39804 18312
rect 41230 18300 41236 18312
rect 41288 18300 41294 18352
rect 41877 18343 41935 18349
rect 41877 18309 41889 18343
rect 41923 18340 41935 18343
rect 42858 18343 42916 18349
rect 42858 18340 42870 18343
rect 41923 18312 42870 18340
rect 41923 18309 41935 18312
rect 41877 18303 41935 18309
rect 42858 18309 42870 18312
rect 42904 18309 42916 18343
rect 42858 18303 42916 18309
rect 56502 18300 56508 18352
rect 56560 18340 56566 18352
rect 56560 18312 57008 18340
rect 56560 18300 56566 18312
rect 39761 18275 39819 18281
rect 39761 18241 39773 18275
rect 39807 18241 39819 18275
rect 39761 18235 39819 18241
rect 40221 18275 40279 18281
rect 40221 18241 40233 18275
rect 40267 18272 40279 18275
rect 41046 18272 41052 18284
rect 40267 18244 41052 18272
rect 40267 18241 40279 18244
rect 40221 18235 40279 18241
rect 36078 18204 36084 18216
rect 34020 18176 34284 18204
rect 35176 18176 36084 18204
rect 34020 18164 34026 18176
rect 23440 18108 27384 18136
rect 23440 18096 23446 18108
rect 16025 18071 16083 18077
rect 16025 18037 16037 18071
rect 16071 18068 16083 18071
rect 18414 18068 18420 18080
rect 16071 18040 18420 18068
rect 16071 18037 16083 18040
rect 16025 18031 16083 18037
rect 18414 18028 18420 18040
rect 18472 18028 18478 18080
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 20622 18068 20628 18080
rect 18656 18040 20628 18068
rect 18656 18028 18662 18040
rect 20622 18028 20628 18040
rect 20680 18068 20686 18080
rect 23658 18068 23664 18080
rect 20680 18040 23664 18068
rect 20680 18028 20686 18040
rect 23658 18028 23664 18040
rect 23716 18028 23722 18080
rect 23753 18071 23811 18077
rect 23753 18037 23765 18071
rect 23799 18068 23811 18071
rect 26326 18068 26332 18080
rect 23799 18040 26332 18068
rect 23799 18037 23811 18040
rect 23753 18031 23811 18037
rect 26326 18028 26332 18040
rect 26384 18028 26390 18080
rect 26418 18028 26424 18080
rect 26476 18068 26482 18080
rect 27249 18071 27307 18077
rect 27249 18068 27261 18071
rect 26476 18040 27261 18068
rect 26476 18028 26482 18040
rect 27249 18037 27261 18040
rect 27295 18037 27307 18071
rect 27356 18068 27384 18108
rect 28966 18108 31754 18136
rect 28966 18068 28994 18108
rect 32674 18096 32680 18148
rect 32732 18136 32738 18148
rect 35176 18136 35204 18176
rect 36078 18164 36084 18176
rect 36136 18164 36142 18216
rect 38562 18164 38568 18216
rect 38620 18204 38626 18216
rect 39776 18204 39804 18235
rect 41046 18232 41052 18244
rect 41104 18232 41110 18284
rect 41782 18272 41788 18284
rect 41743 18244 41788 18272
rect 41782 18232 41788 18244
rect 41840 18232 41846 18284
rect 41969 18275 42027 18281
rect 41969 18241 41981 18275
rect 42015 18241 42027 18275
rect 42610 18272 42616 18284
rect 42571 18244 42616 18272
rect 41969 18235 42027 18241
rect 38620 18176 39804 18204
rect 38620 18164 38626 18176
rect 40034 18164 40040 18216
rect 40092 18204 40098 18216
rect 40313 18207 40371 18213
rect 40313 18204 40325 18207
rect 40092 18176 40325 18204
rect 40092 18164 40098 18176
rect 40313 18173 40325 18176
rect 40359 18173 40371 18207
rect 41984 18204 42012 18235
rect 42610 18232 42616 18244
rect 42668 18232 42674 18284
rect 43162 18272 43168 18284
rect 42720 18244 43168 18272
rect 42720 18204 42748 18244
rect 43162 18232 43168 18244
rect 43220 18232 43226 18284
rect 56686 18232 56692 18284
rect 56744 18272 56750 18284
rect 56873 18275 56931 18281
rect 56873 18272 56885 18275
rect 56744 18244 56885 18272
rect 56744 18232 56750 18244
rect 56873 18241 56885 18244
rect 56919 18241 56931 18275
rect 56980 18272 57008 18312
rect 57882 18300 57888 18352
rect 57940 18340 57946 18352
rect 57940 18312 58296 18340
rect 57940 18300 57946 18312
rect 57974 18272 57980 18284
rect 56980 18244 57980 18272
rect 56873 18235 56931 18241
rect 57974 18232 57980 18244
rect 58032 18272 58038 18284
rect 58268 18281 58296 18312
rect 58069 18275 58127 18281
rect 58069 18272 58081 18275
rect 58032 18244 58081 18272
rect 58032 18232 58038 18244
rect 58069 18241 58081 18244
rect 58115 18241 58127 18275
rect 58069 18235 58127 18241
rect 58253 18275 58311 18281
rect 58253 18241 58265 18275
rect 58299 18241 58311 18275
rect 58253 18235 58311 18241
rect 41984 18176 42748 18204
rect 40313 18167 40371 18173
rect 32732 18108 35204 18136
rect 32732 18096 32738 18108
rect 35250 18096 35256 18148
rect 35308 18136 35314 18148
rect 44266 18136 44272 18148
rect 35308 18108 41414 18136
rect 35308 18096 35314 18108
rect 29178 18068 29184 18080
rect 27356 18040 28994 18068
rect 29139 18040 29184 18068
rect 27249 18031 27307 18037
rect 29178 18028 29184 18040
rect 29236 18028 29242 18080
rect 30742 18028 30748 18080
rect 30800 18068 30806 18080
rect 32766 18068 32772 18080
rect 30800 18040 32772 18068
rect 30800 18028 30806 18040
rect 32766 18028 32772 18040
rect 32824 18028 32830 18080
rect 33318 18068 33324 18080
rect 33279 18040 33324 18068
rect 33318 18028 33324 18040
rect 33376 18028 33382 18080
rect 34698 18028 34704 18080
rect 34756 18068 34762 18080
rect 34977 18071 35035 18077
rect 34977 18068 34989 18071
rect 34756 18040 34989 18068
rect 34756 18028 34762 18040
rect 34977 18037 34989 18040
rect 35023 18037 35035 18071
rect 34977 18031 35035 18037
rect 36354 18028 36360 18080
rect 36412 18068 36418 18080
rect 38105 18071 38163 18077
rect 38105 18068 38117 18071
rect 36412 18040 38117 18068
rect 36412 18028 36418 18040
rect 38105 18037 38117 18040
rect 38151 18037 38163 18071
rect 38105 18031 38163 18037
rect 38838 18028 38844 18080
rect 38896 18068 38902 18080
rect 40218 18068 40224 18080
rect 38896 18040 40224 18068
rect 38896 18028 38902 18040
rect 40218 18028 40224 18040
rect 40276 18028 40282 18080
rect 41386 18068 41414 18108
rect 43548 18108 44272 18136
rect 43548 18068 43576 18108
rect 44266 18096 44272 18108
rect 44324 18096 44330 18148
rect 43990 18068 43996 18080
rect 41386 18040 43576 18068
rect 43951 18040 43996 18068
rect 43990 18028 43996 18040
rect 44048 18028 44054 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 14826 17824 14832 17876
rect 14884 17864 14890 17876
rect 14884 17836 20024 17864
rect 14884 17824 14890 17836
rect 15749 17799 15807 17805
rect 15749 17765 15761 17799
rect 15795 17796 15807 17799
rect 17586 17796 17592 17808
rect 15795 17768 17592 17796
rect 15795 17765 15807 17768
rect 15749 17759 15807 17765
rect 17586 17756 17592 17768
rect 17644 17756 17650 17808
rect 17678 17756 17684 17808
rect 17736 17796 17742 17808
rect 19886 17796 19892 17808
rect 17736 17768 19892 17796
rect 17736 17756 17742 17768
rect 19886 17756 19892 17768
rect 19944 17756 19950 17808
rect 19996 17796 20024 17836
rect 20254 17824 20260 17876
rect 20312 17864 20318 17876
rect 20993 17867 21051 17873
rect 20993 17864 21005 17867
rect 20312 17836 21005 17864
rect 20312 17824 20318 17836
rect 20993 17833 21005 17836
rect 21039 17833 21051 17867
rect 33042 17864 33048 17876
rect 20993 17827 21051 17833
rect 22066 17836 33048 17864
rect 22066 17796 22094 17836
rect 33042 17824 33048 17836
rect 33100 17824 33106 17876
rect 41782 17864 41788 17876
rect 35636 17836 41414 17864
rect 41743 17836 41788 17864
rect 25774 17796 25780 17808
rect 19996 17768 22094 17796
rect 25735 17768 25780 17796
rect 25774 17756 25780 17768
rect 25832 17756 25838 17808
rect 26142 17756 26148 17808
rect 26200 17796 26206 17808
rect 30098 17796 30104 17808
rect 26200 17768 30104 17796
rect 26200 17756 26206 17768
rect 30098 17756 30104 17768
rect 30156 17756 30162 17808
rect 30282 17796 30288 17808
rect 30243 17768 30288 17796
rect 30282 17756 30288 17768
rect 30340 17756 30346 17808
rect 32766 17756 32772 17808
rect 32824 17796 32830 17808
rect 32861 17799 32919 17805
rect 32861 17796 32873 17799
rect 32824 17768 32873 17796
rect 32824 17756 32830 17768
rect 32861 17765 32873 17768
rect 32907 17796 32919 17799
rect 35342 17796 35348 17808
rect 32907 17768 35348 17796
rect 32907 17765 32919 17768
rect 32861 17759 32919 17765
rect 35342 17756 35348 17768
rect 35400 17756 35406 17808
rect 17957 17731 18015 17737
rect 17957 17728 17969 17731
rect 16501 17700 17969 17728
rect 1581 17663 1639 17669
rect 1581 17629 1593 17663
rect 1627 17660 1639 17663
rect 2038 17660 2044 17672
rect 1627 17632 2044 17660
rect 1627 17629 1639 17632
rect 1581 17623 1639 17629
rect 2038 17620 2044 17632
rect 2096 17620 2102 17672
rect 15654 17660 15660 17672
rect 15615 17632 15660 17660
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 16501 17669 16529 17700
rect 17957 17697 17969 17700
rect 18003 17728 18015 17731
rect 18003 17700 22416 17728
rect 18003 17697 18015 17700
rect 17957 17691 18015 17697
rect 16485 17663 16543 17669
rect 16485 17629 16497 17663
rect 16531 17629 16543 17663
rect 17402 17660 17408 17672
rect 17363 17632 17408 17660
rect 16485 17623 16543 17629
rect 17402 17620 17408 17632
rect 17460 17620 17466 17672
rect 18138 17620 18144 17672
rect 18196 17660 18202 17672
rect 18509 17663 18567 17669
rect 18509 17660 18521 17663
rect 18196 17632 18521 17660
rect 18196 17620 18202 17632
rect 18509 17629 18521 17632
rect 18555 17629 18567 17663
rect 18509 17623 18567 17629
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17660 18751 17663
rect 19058 17660 19064 17672
rect 18739 17632 19064 17660
rect 18739 17629 18751 17632
rect 18693 17623 18751 17629
rect 1854 17592 1860 17604
rect 1815 17564 1860 17592
rect 1854 17552 1860 17564
rect 1912 17552 1918 17604
rect 16301 17595 16359 17601
rect 16301 17561 16313 17595
rect 16347 17592 16359 17595
rect 17126 17592 17132 17604
rect 16347 17564 17132 17592
rect 16347 17561 16359 17564
rect 16301 17555 16359 17561
rect 17126 17552 17132 17564
rect 17184 17592 17190 17604
rect 17310 17592 17316 17604
rect 17184 17564 17316 17592
rect 17184 17552 17190 17564
rect 17310 17552 17316 17564
rect 17368 17552 17374 17604
rect 17954 17552 17960 17604
rect 18012 17592 18018 17604
rect 18708 17592 18736 17623
rect 19058 17620 19064 17632
rect 19116 17620 19122 17672
rect 19334 17620 19340 17672
rect 19392 17660 19398 17672
rect 19797 17663 19855 17669
rect 19797 17660 19809 17663
rect 19392 17632 19809 17660
rect 19392 17620 19398 17632
rect 19797 17629 19809 17632
rect 19843 17629 19855 17663
rect 22388 17660 22416 17700
rect 22462 17688 22468 17740
rect 22520 17728 22526 17740
rect 22557 17731 22615 17737
rect 22557 17728 22569 17731
rect 22520 17700 22569 17728
rect 22520 17688 22526 17700
rect 22557 17697 22569 17700
rect 22603 17697 22615 17731
rect 25314 17728 25320 17740
rect 25275 17700 25320 17728
rect 22557 17691 22615 17697
rect 25314 17688 25320 17700
rect 25372 17688 25378 17740
rect 27982 17688 27988 17740
rect 28040 17728 28046 17740
rect 30742 17728 30748 17740
rect 28040 17700 30748 17728
rect 28040 17688 28046 17700
rect 30742 17688 30748 17700
rect 30800 17688 30806 17740
rect 33502 17728 33508 17740
rect 33060 17700 33508 17728
rect 23382 17660 23388 17672
rect 22388 17632 23388 17660
rect 19797 17623 19855 17629
rect 23382 17620 23388 17632
rect 23440 17620 23446 17672
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 24854 17660 24860 17672
rect 24627 17632 24860 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 24854 17620 24860 17632
rect 24912 17620 24918 17672
rect 25409 17663 25467 17669
rect 25409 17629 25421 17663
rect 25455 17629 25467 17663
rect 25409 17623 25467 17629
rect 20346 17592 20352 17604
rect 18012 17564 18736 17592
rect 18800 17564 20352 17592
rect 18012 17552 18018 17564
rect 13078 17484 13084 17536
rect 13136 17524 13142 17536
rect 16577 17527 16635 17533
rect 16577 17524 16589 17527
rect 13136 17496 16589 17524
rect 13136 17484 13142 17496
rect 16577 17493 16589 17496
rect 16623 17524 16635 17527
rect 17678 17524 17684 17536
rect 16623 17496 17684 17524
rect 16623 17493 16635 17496
rect 16577 17487 16635 17493
rect 17678 17484 17684 17496
rect 17736 17484 17742 17536
rect 18322 17484 18328 17536
rect 18380 17524 18386 17536
rect 18800 17524 18828 17564
rect 20346 17552 20352 17564
rect 20404 17552 20410 17604
rect 22824 17595 22882 17601
rect 22824 17561 22836 17595
rect 22870 17592 22882 17595
rect 22922 17592 22928 17604
rect 22870 17564 22928 17592
rect 22870 17561 22882 17564
rect 22824 17555 22882 17561
rect 22922 17552 22928 17564
rect 22980 17552 22986 17604
rect 25424 17592 25452 17623
rect 25498 17620 25504 17672
rect 25556 17660 25562 17672
rect 26237 17663 26295 17669
rect 26237 17660 26249 17663
rect 25556 17632 26249 17660
rect 25556 17620 25562 17632
rect 26237 17629 26249 17632
rect 26283 17660 26295 17663
rect 29178 17660 29184 17672
rect 26283 17632 29184 17660
rect 26283 17629 26295 17632
rect 26237 17623 26295 17629
rect 29178 17620 29184 17632
rect 29236 17620 29242 17672
rect 29753 17663 29811 17669
rect 29753 17660 29765 17663
rect 29288 17632 29765 17660
rect 27890 17592 27896 17604
rect 25424 17564 27896 17592
rect 27890 17552 27896 17564
rect 27948 17552 27954 17604
rect 29086 17552 29092 17604
rect 29144 17592 29150 17604
rect 29288 17592 29316 17632
rect 29753 17629 29765 17632
rect 29799 17629 29811 17663
rect 29753 17623 29811 17629
rect 30106 17663 30164 17669
rect 30106 17629 30118 17663
rect 30152 17660 30164 17663
rect 30558 17660 30564 17672
rect 30152 17632 30564 17660
rect 30152 17629 30164 17632
rect 30106 17623 30164 17629
rect 30558 17620 30564 17632
rect 30616 17620 30622 17672
rect 30834 17620 30840 17672
rect 30892 17660 30898 17672
rect 31110 17660 31116 17672
rect 30892 17632 30937 17660
rect 31071 17632 31116 17660
rect 30892 17620 30898 17632
rect 31110 17620 31116 17632
rect 31168 17620 31174 17672
rect 31570 17620 31576 17672
rect 31628 17660 31634 17672
rect 31757 17663 31815 17669
rect 31757 17660 31769 17663
rect 31628 17632 31769 17660
rect 31628 17620 31634 17632
rect 31757 17629 31769 17632
rect 31803 17629 31815 17663
rect 32030 17660 32036 17672
rect 31991 17632 32036 17660
rect 31757 17623 31815 17629
rect 32030 17620 32036 17632
rect 32088 17620 32094 17672
rect 32125 17663 32183 17669
rect 32125 17629 32137 17663
rect 32171 17660 32183 17663
rect 32858 17660 32864 17672
rect 32171 17632 32864 17660
rect 32171 17629 32183 17632
rect 32125 17623 32183 17629
rect 32858 17620 32864 17632
rect 32916 17620 32922 17672
rect 33060 17669 33088 17700
rect 33502 17688 33508 17700
rect 33560 17688 33566 17740
rect 33045 17663 33103 17669
rect 33045 17629 33057 17663
rect 33091 17629 33103 17663
rect 33045 17623 33103 17629
rect 33134 17620 33140 17672
rect 33192 17660 33198 17672
rect 33321 17663 33379 17669
rect 33192 17632 33237 17660
rect 33192 17620 33198 17632
rect 33321 17629 33333 17663
rect 33367 17629 33379 17663
rect 33321 17623 33379 17629
rect 33413 17663 33471 17669
rect 33413 17629 33425 17663
rect 33459 17660 33471 17663
rect 35636 17660 35664 17836
rect 37645 17799 37703 17805
rect 37645 17796 37657 17799
rect 36832 17768 37657 17796
rect 33459 17632 35664 17660
rect 35713 17663 35771 17669
rect 33459 17629 33471 17632
rect 33413 17623 33471 17629
rect 35713 17629 35725 17663
rect 35759 17660 35771 17663
rect 36538 17660 36544 17672
rect 35759 17632 36544 17660
rect 35759 17629 35771 17632
rect 35713 17623 35771 17629
rect 29144 17564 29316 17592
rect 29144 17552 29150 17564
rect 29454 17552 29460 17604
rect 29512 17592 29518 17604
rect 29917 17595 29975 17601
rect 29917 17592 29929 17595
rect 29512 17564 29929 17592
rect 29512 17552 29518 17564
rect 29917 17561 29929 17564
rect 29963 17561 29975 17595
rect 29917 17555 29975 17561
rect 30009 17595 30067 17601
rect 30009 17561 30021 17595
rect 30055 17592 30067 17595
rect 30055 17564 30144 17592
rect 30055 17561 30067 17564
rect 30009 17555 30067 17561
rect 30116 17536 30144 17564
rect 30190 17552 30196 17604
rect 30248 17592 30254 17604
rect 31938 17592 31944 17604
rect 30248 17564 31754 17592
rect 31851 17564 31944 17592
rect 30248 17552 30254 17564
rect 31726 17536 31754 17564
rect 31938 17552 31944 17564
rect 31996 17592 32002 17604
rect 32582 17592 32588 17604
rect 31996 17564 32588 17592
rect 31996 17552 32002 17564
rect 32582 17552 32588 17564
rect 32640 17552 32646 17604
rect 32876 17592 32904 17620
rect 33226 17592 33232 17604
rect 32876 17564 33232 17592
rect 33226 17552 33232 17564
rect 33284 17552 33290 17604
rect 33336 17592 33364 17623
rect 36538 17620 36544 17632
rect 36596 17620 36602 17672
rect 33962 17592 33968 17604
rect 33336 17564 33968 17592
rect 33962 17552 33968 17564
rect 34020 17552 34026 17604
rect 35980 17595 36038 17601
rect 35980 17561 35992 17595
rect 36026 17592 36038 17595
rect 36832 17592 36860 17768
rect 37645 17765 37657 17768
rect 37691 17765 37703 17799
rect 41386 17796 41414 17836
rect 41782 17824 41788 17836
rect 41840 17824 41846 17876
rect 42242 17796 42248 17808
rect 41386 17768 42248 17796
rect 37645 17759 37703 17765
rect 42242 17756 42248 17768
rect 42300 17756 42306 17808
rect 37918 17688 37924 17740
rect 37976 17728 37982 17740
rect 38197 17731 38255 17737
rect 38197 17728 38209 17731
rect 37976 17700 38209 17728
rect 37976 17688 37982 17700
rect 38197 17697 38209 17700
rect 38243 17697 38255 17731
rect 58158 17728 58164 17740
rect 38197 17691 38255 17697
rect 42260 17700 44036 17728
rect 58119 17700 58164 17728
rect 37826 17620 37832 17672
rect 37884 17660 37890 17672
rect 38013 17663 38071 17669
rect 38013 17660 38025 17663
rect 37884 17632 38025 17660
rect 37884 17620 37890 17632
rect 38013 17629 38025 17632
rect 38059 17629 38071 17663
rect 38013 17623 38071 17629
rect 38102 17620 38108 17672
rect 38160 17660 38166 17672
rect 41230 17660 41236 17672
rect 38160 17632 41236 17660
rect 38160 17620 38166 17632
rect 41230 17620 41236 17632
rect 41288 17620 41294 17672
rect 41966 17663 42024 17669
rect 41966 17629 41978 17663
rect 42012 17660 42024 17663
rect 42260 17660 42288 17700
rect 44008 17672 44036 17700
rect 58158 17688 58164 17700
rect 58216 17688 58222 17740
rect 42012 17632 42288 17660
rect 42337 17663 42395 17669
rect 42012 17629 42024 17632
rect 41966 17623 42024 17629
rect 42337 17629 42349 17663
rect 42383 17629 42395 17663
rect 42337 17623 42395 17629
rect 36026 17564 36860 17592
rect 36026 17561 36038 17564
rect 35980 17555 36038 17561
rect 37734 17552 37740 17604
rect 37792 17592 37798 17604
rect 42352 17592 42380 17623
rect 42426 17620 42432 17672
rect 42484 17660 42490 17672
rect 42484 17632 42529 17660
rect 42484 17620 42490 17632
rect 43990 17620 43996 17672
rect 44048 17660 44054 17672
rect 57885 17663 57943 17669
rect 57885 17660 57897 17663
rect 44048 17632 57897 17660
rect 44048 17620 44054 17632
rect 57885 17629 57897 17632
rect 57931 17629 57943 17663
rect 57885 17623 57943 17629
rect 57054 17592 57060 17604
rect 37792 17564 42380 17592
rect 57015 17564 57060 17592
rect 37792 17552 37798 17564
rect 57054 17552 57060 17564
rect 57112 17552 57118 17604
rect 18380 17496 18828 17524
rect 18877 17527 18935 17533
rect 18380 17484 18386 17496
rect 18877 17493 18889 17527
rect 18923 17524 18935 17527
rect 18966 17524 18972 17536
rect 18923 17496 18972 17524
rect 18923 17493 18935 17496
rect 18877 17487 18935 17493
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 20438 17484 20444 17536
rect 20496 17524 20502 17536
rect 21910 17524 21916 17536
rect 20496 17496 21916 17524
rect 20496 17484 20502 17496
rect 21910 17484 21916 17496
rect 21968 17484 21974 17536
rect 23934 17484 23940 17536
rect 23992 17524 23998 17536
rect 24673 17527 24731 17533
rect 23992 17496 24037 17524
rect 23992 17484 23998 17496
rect 24673 17493 24685 17527
rect 24719 17524 24731 17527
rect 25038 17524 25044 17536
rect 24719 17496 25044 17524
rect 24719 17493 24731 17496
rect 24673 17487 24731 17493
rect 25038 17484 25044 17496
rect 25096 17484 25102 17536
rect 25314 17484 25320 17536
rect 25372 17524 25378 17536
rect 27433 17527 27491 17533
rect 27433 17524 27445 17527
rect 25372 17496 27445 17524
rect 25372 17484 25378 17496
rect 27433 17493 27445 17496
rect 27479 17493 27491 17527
rect 27433 17487 27491 17493
rect 30098 17484 30104 17536
rect 30156 17484 30162 17536
rect 30374 17484 30380 17536
rect 30432 17524 30438 17536
rect 30929 17527 30987 17533
rect 30929 17524 30941 17527
rect 30432 17496 30941 17524
rect 30432 17484 30438 17496
rect 30929 17493 30941 17496
rect 30975 17493 30987 17527
rect 31726 17496 31760 17536
rect 30929 17487 30987 17493
rect 31754 17484 31760 17496
rect 31812 17484 31818 17536
rect 32309 17527 32367 17533
rect 32309 17493 32321 17527
rect 32355 17524 32367 17527
rect 32766 17524 32772 17536
rect 32355 17496 32772 17524
rect 32355 17493 32367 17496
rect 32309 17487 32367 17493
rect 32766 17484 32772 17496
rect 32824 17484 32830 17536
rect 33042 17484 33048 17536
rect 33100 17524 33106 17536
rect 37093 17527 37151 17533
rect 37093 17524 37105 17527
rect 33100 17496 37105 17524
rect 33100 17484 33106 17496
rect 37093 17493 37105 17496
rect 37139 17524 37151 17527
rect 38105 17527 38163 17533
rect 38105 17524 38117 17527
rect 37139 17496 38117 17524
rect 37139 17493 37151 17496
rect 37093 17487 37151 17493
rect 38105 17493 38117 17496
rect 38151 17493 38163 17527
rect 38105 17487 38163 17493
rect 41046 17484 41052 17536
rect 41104 17524 41110 17536
rect 41969 17527 42027 17533
rect 41969 17524 41981 17527
rect 41104 17496 41981 17524
rect 41104 17484 41110 17496
rect 41969 17493 41981 17496
rect 42015 17493 42027 17527
rect 41969 17487 42027 17493
rect 46198 17484 46204 17536
rect 46256 17524 46262 17536
rect 57149 17527 57207 17533
rect 57149 17524 57161 17527
rect 46256 17496 57161 17524
rect 46256 17484 46262 17496
rect 57149 17493 57161 17496
rect 57195 17493 57207 17527
rect 57149 17487 57207 17493
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 15654 17280 15660 17332
rect 15712 17320 15718 17332
rect 16942 17320 16948 17332
rect 15712 17292 16948 17320
rect 15712 17280 15718 17292
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 18414 17320 18420 17332
rect 17604 17292 18420 17320
rect 2130 17212 2136 17264
rect 2188 17252 2194 17264
rect 11606 17252 11612 17264
rect 2188 17224 11612 17252
rect 2188 17212 2194 17224
rect 11606 17212 11612 17224
rect 11664 17212 11670 17264
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17184 1639 17187
rect 12342 17184 12348 17196
rect 1627 17156 12348 17184
rect 1627 17153 1639 17156
rect 1581 17147 1639 17153
rect 12342 17144 12348 17156
rect 12400 17144 12406 17196
rect 15657 17187 15715 17193
rect 15657 17153 15669 17187
rect 15703 17184 15715 17187
rect 17034 17184 17040 17196
rect 15703 17156 17040 17184
rect 15703 17153 15715 17156
rect 15657 17147 15715 17153
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 17402 17184 17408 17196
rect 17363 17156 17408 17184
rect 17402 17144 17408 17156
rect 17460 17144 17466 17196
rect 17604 17184 17632 17292
rect 18414 17280 18420 17292
rect 18472 17320 18478 17332
rect 19150 17320 19156 17332
rect 18472 17292 19156 17320
rect 18472 17280 18478 17292
rect 19150 17280 19156 17292
rect 19208 17280 19214 17332
rect 19981 17323 20039 17329
rect 19981 17289 19993 17323
rect 20027 17289 20039 17323
rect 19981 17283 20039 17289
rect 21453 17323 21511 17329
rect 21453 17289 21465 17323
rect 21499 17320 21511 17323
rect 24302 17320 24308 17332
rect 21499 17292 24308 17320
rect 21499 17289 21511 17292
rect 21453 17283 21511 17289
rect 17678 17212 17684 17264
rect 17736 17252 17742 17264
rect 18874 17252 18880 17264
rect 17736 17224 18880 17252
rect 17736 17212 17742 17224
rect 18874 17212 18880 17224
rect 18932 17212 18938 17264
rect 19058 17252 19064 17264
rect 18971 17224 19064 17252
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 17604 17156 17785 17184
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 17773 17147 17831 17153
rect 17862 17144 17868 17196
rect 17920 17184 17926 17196
rect 18984 17193 19012 17224
rect 19058 17212 19064 17224
rect 19116 17252 19122 17264
rect 19996 17252 20024 17283
rect 24302 17280 24308 17292
rect 24360 17280 24366 17332
rect 24394 17280 24400 17332
rect 24452 17320 24458 17332
rect 30190 17320 30196 17332
rect 24452 17292 30196 17320
rect 24452 17280 24458 17292
rect 30190 17280 30196 17292
rect 30248 17280 30254 17332
rect 30374 17280 30380 17332
rect 30432 17280 30438 17332
rect 30558 17280 30564 17332
rect 30616 17320 30622 17332
rect 31846 17320 31852 17332
rect 30616 17292 31852 17320
rect 30616 17280 30622 17292
rect 31846 17280 31852 17292
rect 31904 17280 31910 17332
rect 33502 17280 33508 17332
rect 33560 17320 33566 17332
rect 34885 17323 34943 17329
rect 34885 17320 34897 17323
rect 33560 17292 34897 17320
rect 33560 17280 33566 17292
rect 34885 17289 34897 17292
rect 34931 17289 34943 17323
rect 34885 17283 34943 17289
rect 39390 17280 39396 17332
rect 39448 17320 39454 17332
rect 40954 17320 40960 17332
rect 39448 17292 40960 17320
rect 39448 17280 39454 17292
rect 40954 17280 40960 17292
rect 41012 17280 41018 17332
rect 41046 17280 41052 17332
rect 41104 17280 41110 17332
rect 41230 17280 41236 17332
rect 41288 17320 41294 17332
rect 45554 17320 45560 17332
rect 41288 17292 45560 17320
rect 41288 17280 41294 17292
rect 45554 17280 45560 17292
rect 45612 17280 45618 17332
rect 19116 17224 20024 17252
rect 20993 17255 21051 17261
rect 19116 17212 19122 17224
rect 20993 17221 21005 17255
rect 21039 17252 21051 17255
rect 21082 17252 21088 17264
rect 21039 17224 21088 17252
rect 21039 17221 21051 17224
rect 20993 17215 21051 17221
rect 21082 17212 21088 17224
rect 21140 17212 21146 17264
rect 21174 17212 21180 17264
rect 21232 17252 21238 17264
rect 21232 17224 22784 17252
rect 21232 17212 21238 17224
rect 18693 17187 18751 17193
rect 18693 17184 18705 17187
rect 17920 17156 18705 17184
rect 17920 17144 17926 17156
rect 18693 17153 18705 17156
rect 18739 17153 18751 17187
rect 18693 17147 18751 17153
rect 18969 17187 19027 17193
rect 18969 17153 18981 17187
rect 19015 17153 19027 17187
rect 19886 17184 19892 17196
rect 18969 17147 19027 17153
rect 19076 17156 19892 17184
rect 1762 17116 1768 17128
rect 1723 17088 1768 17116
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 14734 17076 14740 17128
rect 14792 17116 14798 17128
rect 19076 17116 19104 17156
rect 19886 17144 19892 17156
rect 19944 17144 19950 17196
rect 19981 17187 20039 17193
rect 19981 17153 19993 17187
rect 20027 17184 20039 17187
rect 20070 17184 20076 17196
rect 20027 17156 20076 17184
rect 20027 17153 20039 17156
rect 19981 17147 20039 17153
rect 20070 17144 20076 17156
rect 20128 17144 20134 17196
rect 20165 17187 20223 17193
rect 20165 17153 20177 17187
rect 20211 17153 20223 17187
rect 20346 17184 20352 17196
rect 20307 17156 20352 17184
rect 20165 17147 20223 17153
rect 19242 17116 19248 17128
rect 14792 17088 19104 17116
rect 19203 17088 19248 17116
rect 14792 17076 14798 17088
rect 19242 17076 19248 17088
rect 19300 17076 19306 17128
rect 19426 17076 19432 17128
rect 19484 17116 19490 17128
rect 20180 17116 20208 17147
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 21910 17144 21916 17196
rect 21968 17184 21974 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21968 17156 22017 17184
rect 21968 17144 21974 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22189 17187 22247 17193
rect 22189 17153 22201 17187
rect 22235 17184 22247 17187
rect 22646 17184 22652 17196
rect 22235 17156 22652 17184
rect 22235 17153 22247 17156
rect 22189 17147 22247 17153
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 22756 17187 22784 17224
rect 23934 17212 23940 17264
rect 23992 17252 23998 17264
rect 25498 17252 25504 17264
rect 23992 17224 25504 17252
rect 23992 17212 23998 17224
rect 25498 17212 25504 17224
rect 25556 17212 25562 17264
rect 25682 17212 25688 17264
rect 25740 17252 25746 17264
rect 26142 17252 26148 17264
rect 25740 17224 26148 17252
rect 25740 17212 25746 17224
rect 26142 17212 26148 17224
rect 26200 17212 26206 17264
rect 27062 17252 27068 17264
rect 26344 17224 27068 17252
rect 22833 17187 22891 17193
rect 22756 17159 22845 17187
rect 22833 17153 22845 17159
rect 22879 17153 22891 17187
rect 26234 17184 26240 17196
rect 26195 17156 26240 17184
rect 22833 17147 22891 17153
rect 26234 17144 26240 17156
rect 26292 17144 26298 17196
rect 26344 17193 26372 17224
rect 27062 17212 27068 17224
rect 27120 17212 27126 17264
rect 28902 17252 28908 17264
rect 28863 17224 28908 17252
rect 28902 17212 28908 17224
rect 28960 17212 28966 17264
rect 29454 17212 29460 17264
rect 29512 17252 29518 17264
rect 30392 17252 30420 17280
rect 31662 17252 31668 17264
rect 29512 17224 29960 17252
rect 29512 17212 29518 17224
rect 26329 17187 26387 17193
rect 26329 17153 26341 17187
rect 26375 17153 26387 17187
rect 26329 17147 26387 17153
rect 26418 17144 26424 17196
rect 26476 17184 26482 17196
rect 26605 17187 26663 17193
rect 26476 17156 26521 17184
rect 26476 17144 26482 17156
rect 26605 17153 26617 17187
rect 26651 17153 26663 17187
rect 26605 17147 26663 17153
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17184 27215 17187
rect 29822 17184 29828 17196
rect 27203 17156 29828 17184
rect 27203 17153 27215 17156
rect 27157 17147 27215 17153
rect 25406 17116 25412 17128
rect 19484 17088 20208 17116
rect 21376 17088 25412 17116
rect 19484 17076 19490 17088
rect 17126 17008 17132 17060
rect 17184 17048 17190 17060
rect 17221 17051 17279 17057
rect 17221 17048 17233 17051
rect 17184 17020 17233 17048
rect 17184 17008 17190 17020
rect 17221 17017 17233 17020
rect 17267 17017 17279 17051
rect 17221 17011 17279 17017
rect 17494 17008 17500 17060
rect 17552 17048 17558 17060
rect 18785 17051 18843 17057
rect 18785 17048 18797 17051
rect 17552 17020 18797 17048
rect 17552 17008 17558 17020
rect 18785 17017 18797 17020
rect 18831 17017 18843 17051
rect 18785 17011 18843 17017
rect 18874 17008 18880 17060
rect 18932 17048 18938 17060
rect 21376 17057 21404 17088
rect 25406 17076 25412 17088
rect 25464 17076 25470 17128
rect 26620 17116 26648 17147
rect 29822 17144 29828 17156
rect 29880 17144 29886 17196
rect 29932 17184 29960 17224
rect 30208 17224 30420 17252
rect 30484 17224 31668 17252
rect 30208 17193 30236 17224
rect 30484 17196 30512 17224
rect 31662 17212 31668 17224
rect 31720 17212 31726 17264
rect 32493 17255 32551 17261
rect 32493 17252 32505 17255
rect 32140 17224 32505 17252
rect 29989 17187 30047 17193
rect 29989 17184 30001 17187
rect 29932 17156 30001 17184
rect 29989 17153 30001 17156
rect 30035 17153 30047 17187
rect 29989 17147 30047 17153
rect 30082 17187 30140 17193
rect 30082 17153 30094 17187
rect 30128 17184 30140 17187
rect 30193 17187 30251 17193
rect 30128 17153 30141 17184
rect 30082 17147 30141 17153
rect 30193 17153 30205 17187
rect 30239 17153 30251 17187
rect 30193 17147 30251 17153
rect 30377 17187 30435 17193
rect 30377 17153 30389 17187
rect 30423 17184 30435 17187
rect 30466 17184 30472 17196
rect 30423 17156 30472 17184
rect 30423 17153 30435 17156
rect 30377 17147 30435 17153
rect 26878 17116 26884 17128
rect 26620 17088 26884 17116
rect 26878 17076 26884 17088
rect 26936 17116 26942 17128
rect 29730 17116 29736 17128
rect 26936 17088 29736 17116
rect 26936 17076 26942 17088
rect 29730 17076 29736 17088
rect 29788 17076 29794 17128
rect 30113 17116 30141 17147
rect 30466 17144 30472 17156
rect 30524 17144 30530 17196
rect 30837 17187 30895 17193
rect 30837 17153 30849 17187
rect 30883 17184 30895 17187
rect 31478 17184 31484 17196
rect 30883 17156 31484 17184
rect 30883 17153 30895 17156
rect 30837 17147 30895 17153
rect 31478 17144 31484 17156
rect 31536 17144 31542 17196
rect 31938 17144 31944 17196
rect 31996 17184 32002 17196
rect 32140 17184 32168 17224
rect 32493 17221 32505 17224
rect 32539 17221 32551 17255
rect 32493 17215 32551 17221
rect 33226 17212 33232 17264
rect 33284 17252 33290 17264
rect 33597 17255 33655 17261
rect 33597 17252 33609 17255
rect 33284 17224 33609 17252
rect 33284 17212 33290 17224
rect 33597 17221 33609 17224
rect 33643 17252 33655 17255
rect 35894 17252 35900 17264
rect 33643 17224 35900 17252
rect 33643 17221 33655 17224
rect 33597 17215 33655 17221
rect 35894 17212 35900 17224
rect 35952 17252 35958 17264
rect 38102 17252 38108 17264
rect 35952 17224 38108 17252
rect 35952 17212 35958 17224
rect 38102 17212 38108 17224
rect 38160 17212 38166 17264
rect 40034 17252 40040 17264
rect 39224 17224 40040 17252
rect 32306 17184 32312 17196
rect 31996 17156 32168 17184
rect 32267 17156 32312 17184
rect 31996 17144 32002 17156
rect 32306 17144 32312 17156
rect 32364 17144 32370 17196
rect 32766 17144 32772 17196
rect 32824 17184 32830 17196
rect 33321 17187 33379 17193
rect 33321 17184 33333 17187
rect 32824 17156 33333 17184
rect 32824 17144 32830 17156
rect 33321 17153 33333 17156
rect 33367 17153 33379 17187
rect 33321 17147 33379 17153
rect 33469 17187 33527 17193
rect 33469 17153 33481 17187
rect 33515 17153 33527 17187
rect 33686 17187 33744 17193
rect 33686 17184 33698 17187
rect 33469 17147 33527 17153
rect 33612 17156 33698 17184
rect 30926 17116 30932 17128
rect 30113 17088 30932 17116
rect 30926 17076 30932 17088
rect 30984 17116 30990 17128
rect 31021 17119 31079 17125
rect 31021 17116 31033 17119
rect 30984 17088 31033 17116
rect 30984 17076 30990 17088
rect 31021 17085 31033 17088
rect 31067 17085 31079 17119
rect 31021 17079 31079 17085
rect 32122 17076 32128 17128
rect 32180 17116 32186 17128
rect 32677 17119 32735 17125
rect 32677 17116 32689 17119
rect 32180 17088 32689 17116
rect 32180 17076 32186 17088
rect 32677 17085 32689 17088
rect 32723 17085 32735 17119
rect 32677 17079 32735 17085
rect 21361 17051 21419 17057
rect 18932 17020 21312 17048
rect 18932 17008 18938 17020
rect 15194 16940 15200 16992
rect 15252 16980 15258 16992
rect 15749 16983 15807 16989
rect 15749 16980 15761 16983
rect 15252 16952 15761 16980
rect 15252 16940 15258 16952
rect 15749 16949 15761 16952
rect 15795 16949 15807 16983
rect 15749 16943 15807 16949
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 21174 16980 21180 16992
rect 16724 16952 21180 16980
rect 16724 16940 16730 16952
rect 21174 16940 21180 16952
rect 21232 16940 21238 16992
rect 21284 16980 21312 17020
rect 21361 17017 21373 17051
rect 21407 17017 21419 17051
rect 24029 17051 24087 17057
rect 24029 17048 24041 17051
rect 21361 17011 21419 17017
rect 21468 17020 24041 17048
rect 21468 16980 21496 17020
rect 24029 17017 24041 17020
rect 24075 17017 24087 17051
rect 24029 17011 24087 17017
rect 25498 17008 25504 17060
rect 25556 17048 25562 17060
rect 25556 17020 30149 17048
rect 25556 17008 25562 17020
rect 21284 16952 21496 16980
rect 22373 16983 22431 16989
rect 22373 16949 22385 16983
rect 22419 16980 22431 16983
rect 25682 16980 25688 16992
rect 22419 16952 25688 16980
rect 22419 16949 22431 16952
rect 22373 16943 22431 16949
rect 25682 16940 25688 16952
rect 25740 16940 25746 16992
rect 25961 16983 26019 16989
rect 25961 16949 25973 16983
rect 26007 16980 26019 16983
rect 29546 16980 29552 16992
rect 26007 16952 29552 16980
rect 26007 16949 26019 16952
rect 25961 16943 26019 16949
rect 29546 16940 29552 16952
rect 29604 16940 29610 16992
rect 29730 16980 29736 16992
rect 29691 16952 29736 16980
rect 29730 16940 29736 16952
rect 29788 16940 29794 16992
rect 30121 16980 30149 17020
rect 30190 17008 30196 17060
rect 30248 17048 30254 17060
rect 31110 17048 31116 17060
rect 30248 17020 31116 17048
rect 30248 17008 30254 17020
rect 31110 17008 31116 17020
rect 31168 17008 31174 17060
rect 31018 16980 31024 16992
rect 30121 16952 31024 16980
rect 31018 16940 31024 16952
rect 31076 16940 31082 16992
rect 31846 16940 31852 16992
rect 31904 16980 31910 16992
rect 32306 16980 32312 16992
rect 31904 16952 32312 16980
rect 31904 16940 31910 16952
rect 32306 16940 32312 16952
rect 32364 16940 32370 16992
rect 33484 16980 33512 17147
rect 33612 17060 33640 17156
rect 33686 17153 33698 17156
rect 33732 17153 33744 17187
rect 33686 17147 33744 17153
rect 33778 17144 33784 17196
rect 33836 17193 33842 17196
rect 33836 17184 33844 17193
rect 33836 17156 33881 17184
rect 33836 17147 33844 17156
rect 33836 17144 33842 17147
rect 33962 17144 33968 17196
rect 34020 17184 34026 17196
rect 34425 17187 34483 17193
rect 34425 17184 34437 17187
rect 34020 17156 34437 17184
rect 34020 17144 34026 17156
rect 34425 17153 34437 17156
rect 34471 17153 34483 17187
rect 34698 17184 34704 17196
rect 34659 17156 34704 17184
rect 34425 17147 34483 17153
rect 34698 17144 34704 17156
rect 34756 17144 34762 17196
rect 39022 17184 39028 17196
rect 38983 17156 39028 17184
rect 39022 17144 39028 17156
rect 39080 17144 39086 17196
rect 39224 17193 39252 17224
rect 40034 17212 40040 17224
rect 40092 17212 40098 17264
rect 40129 17255 40187 17261
rect 40129 17221 40141 17255
rect 40175 17252 40187 17255
rect 40586 17252 40592 17264
rect 40175 17224 40592 17252
rect 40175 17221 40187 17224
rect 40129 17215 40187 17221
rect 40586 17212 40592 17224
rect 40644 17252 40650 17264
rect 41064 17252 41092 17280
rect 40644 17224 41092 17252
rect 40644 17212 40650 17224
rect 39209 17187 39267 17193
rect 39209 17153 39221 17187
rect 39255 17153 39267 17187
rect 39209 17147 39267 17153
rect 39853 17187 39911 17193
rect 39853 17153 39865 17187
rect 39899 17184 39911 17187
rect 40402 17184 40408 17196
rect 39899 17156 40408 17184
rect 39899 17153 39911 17156
rect 39853 17147 39911 17153
rect 40402 17144 40408 17156
rect 40460 17184 40466 17196
rect 41414 17184 41420 17196
rect 40460 17156 41420 17184
rect 40460 17144 40466 17156
rect 41414 17144 41420 17156
rect 41472 17144 41478 17196
rect 57054 17184 57060 17196
rect 57015 17156 57060 17184
rect 57054 17144 57060 17156
rect 57112 17144 57118 17196
rect 34517 17119 34575 17125
rect 34517 17085 34529 17119
rect 34563 17116 34575 17119
rect 36814 17116 36820 17128
rect 34563 17088 36820 17116
rect 34563 17085 34575 17088
rect 34517 17079 34575 17085
rect 36814 17076 36820 17088
rect 36872 17076 36878 17128
rect 36998 17076 37004 17128
rect 37056 17116 37062 17128
rect 46198 17116 46204 17128
rect 37056 17088 46204 17116
rect 37056 17076 37062 17088
rect 46198 17076 46204 17088
rect 46256 17076 46262 17128
rect 57330 17116 57336 17128
rect 57291 17088 57336 17116
rect 57330 17076 57336 17088
rect 57388 17076 57394 17128
rect 33594 17008 33600 17060
rect 33652 17008 33658 17060
rect 33962 17008 33968 17060
rect 34020 17048 34026 17060
rect 40678 17048 40684 17060
rect 34020 17020 34065 17048
rect 39316 17020 40684 17048
rect 34020 17008 34026 17020
rect 39316 16980 39344 17020
rect 40678 17008 40684 17020
rect 40736 17008 40742 17060
rect 33484 16952 39344 16980
rect 39393 16983 39451 16989
rect 39393 16949 39405 16983
rect 39439 16980 39451 16983
rect 39758 16980 39764 16992
rect 39439 16952 39764 16980
rect 39439 16949 39451 16952
rect 39393 16943 39451 16949
rect 39758 16940 39764 16952
rect 39816 16940 39822 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 14826 16736 14832 16788
rect 14884 16736 14890 16788
rect 16666 16776 16672 16788
rect 16627 16748 16672 16776
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 22554 16776 22560 16788
rect 16960 16748 22560 16776
rect 9646 16680 11744 16708
rect 2222 16600 2228 16652
rect 2280 16640 2286 16652
rect 9646 16640 9674 16680
rect 11330 16640 11336 16652
rect 2280 16612 9674 16640
rect 11291 16612 11336 16640
rect 2280 16600 2286 16612
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 11716 16649 11744 16680
rect 11701 16643 11759 16649
rect 11701 16609 11713 16643
rect 11747 16609 11759 16643
rect 14734 16640 14740 16652
rect 14695 16612 14740 16640
rect 11701 16603 11759 16609
rect 14734 16600 14740 16612
rect 14792 16600 14798 16652
rect 14844 16649 14872 16736
rect 14829 16643 14887 16649
rect 14829 16609 14841 16643
rect 14875 16609 14887 16643
rect 14829 16603 14887 16609
rect 15013 16643 15071 16649
rect 15013 16609 15025 16643
rect 15059 16609 15071 16643
rect 15013 16603 15071 16609
rect 11238 16572 11244 16584
rect 11199 16544 11244 16572
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 11606 16572 11612 16584
rect 11567 16544 11612 16572
rect 11606 16532 11612 16544
rect 11664 16532 11670 16584
rect 14918 16572 14924 16584
rect 14879 16544 14924 16572
rect 14918 16532 14924 16544
rect 14976 16532 14982 16584
rect 10502 16464 10508 16516
rect 10560 16504 10566 16516
rect 10597 16507 10655 16513
rect 10597 16504 10609 16507
rect 10560 16476 10609 16504
rect 10560 16464 10566 16476
rect 10597 16473 10609 16476
rect 10643 16473 10655 16507
rect 10597 16467 10655 16473
rect 12342 16396 12348 16448
rect 12400 16436 12406 16448
rect 14553 16439 14611 16445
rect 14553 16436 14565 16439
rect 12400 16408 14565 16436
rect 12400 16396 12406 16408
rect 14553 16405 14565 16408
rect 14599 16405 14611 16439
rect 14553 16399 14611 16405
rect 14918 16396 14924 16448
rect 14976 16436 14982 16448
rect 15028 16436 15056 16603
rect 16025 16575 16083 16581
rect 16025 16541 16037 16575
rect 16071 16541 16083 16575
rect 16206 16572 16212 16584
rect 16167 16544 16212 16572
rect 16025 16535 16083 16541
rect 16040 16504 16068 16535
rect 16206 16532 16212 16544
rect 16264 16532 16270 16584
rect 16666 16572 16672 16584
rect 16627 16544 16672 16572
rect 16666 16532 16672 16544
rect 16724 16532 16730 16584
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16572 16911 16575
rect 16960 16572 16988 16748
rect 22554 16736 22560 16748
rect 22612 16736 22618 16788
rect 22922 16776 22928 16788
rect 22883 16748 22928 16776
rect 22922 16736 22928 16748
rect 22980 16736 22986 16788
rect 24578 16776 24584 16788
rect 24539 16748 24584 16776
rect 24578 16736 24584 16748
rect 24636 16736 24642 16788
rect 24854 16736 24860 16788
rect 24912 16776 24918 16788
rect 26142 16776 26148 16788
rect 24912 16748 26148 16776
rect 24912 16736 24918 16748
rect 26142 16736 26148 16748
rect 26200 16736 26206 16788
rect 26804 16748 27016 16776
rect 17865 16711 17923 16717
rect 17865 16677 17877 16711
rect 17911 16708 17923 16711
rect 19567 16711 19625 16717
rect 19567 16708 19579 16711
rect 17911 16680 19579 16708
rect 17911 16677 17923 16680
rect 17865 16671 17923 16677
rect 19567 16677 19579 16680
rect 19613 16677 19625 16711
rect 19567 16671 19625 16677
rect 20993 16711 21051 16717
rect 20993 16677 21005 16711
rect 21039 16708 21051 16711
rect 21358 16708 21364 16720
rect 21039 16680 21364 16708
rect 21039 16677 21051 16680
rect 20993 16671 21051 16677
rect 21358 16668 21364 16680
rect 21416 16668 21422 16720
rect 25682 16708 25688 16720
rect 24964 16680 25688 16708
rect 18966 16600 18972 16652
rect 19024 16640 19030 16652
rect 19797 16643 19855 16649
rect 19797 16640 19809 16643
rect 19024 16612 19809 16640
rect 19024 16600 19030 16612
rect 19797 16609 19809 16612
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 19886 16600 19892 16652
rect 19944 16640 19950 16652
rect 24394 16640 24400 16652
rect 19944 16612 24400 16640
rect 19944 16600 19950 16612
rect 24394 16600 24400 16612
rect 24452 16600 24458 16652
rect 24486 16600 24492 16652
rect 24544 16640 24550 16652
rect 24964 16640 24992 16680
rect 25682 16668 25688 16680
rect 25740 16668 25746 16720
rect 26804 16708 26832 16748
rect 26068 16680 26832 16708
rect 24544 16612 24808 16640
rect 24544 16600 24550 16612
rect 16899 16544 16988 16572
rect 17313 16575 17371 16581
rect 16899 16541 16911 16544
rect 16853 16535 16911 16541
rect 17313 16541 17325 16575
rect 17359 16541 17371 16575
rect 17586 16572 17592 16584
rect 17547 16544 17592 16572
rect 17313 16535 17371 16541
rect 16574 16504 16580 16516
rect 16040 16476 16580 16504
rect 16574 16464 16580 16476
rect 16632 16464 16638 16516
rect 16758 16464 16764 16516
rect 16816 16504 16822 16516
rect 17328 16504 17356 16535
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 17681 16575 17739 16581
rect 17681 16541 17693 16575
rect 17727 16572 17739 16575
rect 17770 16572 17776 16584
rect 17727 16544 17776 16572
rect 17727 16541 17739 16544
rect 17681 16535 17739 16541
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 18506 16572 18512 16584
rect 17880 16544 18512 16572
rect 16816 16476 17356 16504
rect 16816 16464 16822 16476
rect 14976 16408 15056 16436
rect 14976 16396 14982 16408
rect 16022 16396 16028 16448
rect 16080 16436 16086 16448
rect 16117 16439 16175 16445
rect 16117 16436 16129 16439
rect 16080 16408 16129 16436
rect 16080 16396 16086 16408
rect 16117 16405 16129 16408
rect 16163 16405 16175 16439
rect 17328 16436 17356 16476
rect 17497 16507 17555 16513
rect 17497 16473 17509 16507
rect 17543 16504 17555 16507
rect 17880 16504 17908 16544
rect 18506 16532 18512 16544
rect 18564 16532 18570 16584
rect 18601 16575 18659 16581
rect 18601 16541 18613 16575
rect 18647 16541 18659 16575
rect 18782 16572 18788 16584
rect 18743 16544 18788 16572
rect 18601 16535 18659 16541
rect 18616 16504 18644 16535
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16572 18935 16575
rect 19058 16572 19064 16584
rect 18923 16544 19064 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19058 16532 19064 16544
rect 19116 16532 19122 16584
rect 19242 16532 19248 16584
rect 19300 16572 19306 16584
rect 19659 16575 19717 16581
rect 19659 16572 19671 16575
rect 19300 16544 19671 16572
rect 19300 16532 19306 16544
rect 19659 16541 19671 16544
rect 19705 16541 19717 16575
rect 20622 16572 20628 16584
rect 20583 16544 20628 16572
rect 19659 16535 19717 16541
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 21726 16572 21732 16584
rect 21687 16544 21732 16572
rect 21726 16532 21732 16544
rect 21784 16532 21790 16584
rect 24780 16581 24808 16612
rect 24872 16612 24992 16640
rect 25041 16643 25099 16649
rect 24872 16581 24900 16612
rect 25041 16609 25053 16643
rect 25087 16640 25099 16643
rect 26068 16640 26096 16680
rect 26878 16668 26884 16720
rect 26936 16668 26942 16720
rect 26326 16640 26332 16652
rect 25087 16612 26096 16640
rect 26160 16612 26332 16640
rect 25087 16609 25099 16612
rect 25041 16603 25099 16609
rect 24765 16575 24823 16581
rect 24765 16541 24777 16575
rect 24811 16541 24823 16575
rect 24765 16535 24823 16541
rect 24857 16575 24915 16581
rect 24857 16541 24869 16575
rect 24903 16541 24915 16575
rect 25130 16572 25136 16584
rect 25091 16544 25136 16572
rect 24857 16535 24915 16541
rect 25130 16532 25136 16544
rect 25188 16532 25194 16584
rect 25406 16532 25412 16584
rect 25464 16572 25470 16584
rect 26160 16581 26188 16612
rect 26326 16600 26332 16612
rect 26384 16600 26390 16652
rect 26896 16640 26924 16668
rect 26436 16612 26924 16640
rect 26988 16640 27016 16748
rect 30466 16736 30472 16788
rect 30524 16776 30530 16788
rect 31665 16779 31723 16785
rect 30524 16748 31616 16776
rect 30524 16736 30530 16748
rect 28534 16668 28540 16720
rect 28592 16708 28598 16720
rect 29362 16708 29368 16720
rect 28592 16680 29368 16708
rect 28592 16668 28598 16680
rect 29362 16668 29368 16680
rect 29420 16668 29426 16720
rect 31588 16708 31616 16748
rect 31665 16745 31677 16779
rect 31711 16776 31723 16779
rect 37734 16776 37740 16788
rect 31711 16748 37740 16776
rect 31711 16745 31723 16748
rect 31665 16739 31723 16745
rect 37734 16736 37740 16748
rect 37792 16736 37798 16788
rect 40034 16776 40040 16788
rect 39995 16748 40040 16776
rect 40034 16736 40040 16748
rect 40092 16736 40098 16788
rect 33045 16711 33103 16717
rect 33045 16708 33057 16711
rect 31588 16680 33057 16708
rect 33045 16677 33057 16680
rect 33091 16677 33103 16711
rect 33045 16671 33103 16677
rect 34422 16668 34428 16720
rect 34480 16708 34486 16720
rect 34480 16680 40264 16708
rect 34480 16668 34486 16680
rect 29822 16640 29828 16652
rect 26988 16612 29684 16640
rect 29783 16612 29828 16640
rect 26053 16575 26111 16581
rect 26053 16572 26065 16575
rect 25464 16544 26065 16572
rect 25464 16532 25470 16544
rect 26053 16541 26065 16544
rect 26099 16541 26111 16575
rect 26053 16535 26111 16541
rect 26145 16575 26203 16581
rect 26145 16541 26157 16575
rect 26191 16541 26203 16575
rect 26145 16535 26203 16541
rect 26234 16532 26240 16584
rect 26292 16572 26298 16584
rect 26436 16581 26464 16612
rect 26421 16575 26479 16581
rect 26292 16544 26337 16572
rect 26292 16532 26298 16544
rect 26421 16541 26433 16575
rect 26467 16541 26479 16575
rect 26878 16572 26884 16584
rect 26839 16544 26884 16572
rect 26421 16535 26479 16541
rect 26878 16532 26884 16544
rect 26936 16572 26942 16584
rect 26936 16544 28994 16572
rect 26936 16532 26942 16544
rect 17543 16476 17908 16504
rect 18248 16476 18644 16504
rect 17543 16473 17555 16476
rect 17497 16467 17555 16473
rect 18248 16436 18276 16476
rect 18966 16464 18972 16516
rect 19024 16504 19030 16516
rect 19429 16507 19487 16513
rect 19429 16504 19441 16507
rect 19024 16476 19441 16504
rect 19024 16464 19030 16476
rect 19429 16473 19441 16476
rect 19475 16473 19487 16507
rect 19429 16467 19487 16473
rect 20165 16507 20223 16513
rect 20165 16473 20177 16507
rect 20211 16504 20223 16507
rect 20438 16504 20444 16516
rect 20211 16476 20444 16504
rect 20211 16473 20223 16476
rect 20165 16467 20223 16473
rect 20438 16464 20444 16476
rect 20496 16464 20502 16516
rect 21174 16464 21180 16516
rect 21232 16504 21238 16516
rect 21232 16476 28120 16504
rect 21232 16464 21238 16476
rect 17328 16408 18276 16436
rect 18325 16439 18383 16445
rect 16117 16399 16175 16405
rect 18325 16405 18337 16439
rect 18371 16436 18383 16439
rect 18782 16436 18788 16448
rect 18371 16408 18788 16436
rect 18371 16405 18383 16408
rect 18325 16399 18383 16405
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 20990 16396 20996 16448
rect 21048 16436 21054 16448
rect 21085 16439 21143 16445
rect 21085 16436 21097 16439
rect 21048 16408 21097 16436
rect 21048 16396 21054 16408
rect 21085 16405 21097 16408
rect 21131 16405 21143 16439
rect 25406 16436 25412 16448
rect 25367 16408 25412 16436
rect 21085 16399 21143 16405
rect 25406 16396 25412 16408
rect 25464 16396 25470 16448
rect 25777 16439 25835 16445
rect 25777 16405 25789 16439
rect 25823 16436 25835 16439
rect 27430 16436 27436 16448
rect 25823 16408 27436 16436
rect 25823 16405 25835 16408
rect 25777 16399 25835 16405
rect 27430 16396 27436 16408
rect 27488 16396 27494 16448
rect 28092 16445 28120 16476
rect 28077 16439 28135 16445
rect 28077 16405 28089 16439
rect 28123 16405 28135 16439
rect 28966 16436 28994 16544
rect 29656 16504 29684 16612
rect 29822 16600 29828 16612
rect 29880 16600 29886 16652
rect 31754 16600 31760 16652
rect 31812 16640 31818 16652
rect 32125 16643 32183 16649
rect 31812 16612 31984 16640
rect 31812 16600 31818 16612
rect 29730 16532 29736 16584
rect 29788 16572 29794 16584
rect 30081 16575 30139 16581
rect 30081 16572 30093 16575
rect 29788 16544 30093 16572
rect 29788 16532 29794 16544
rect 30081 16541 30093 16544
rect 30127 16541 30139 16575
rect 30081 16535 30139 16541
rect 31570 16532 31576 16584
rect 31628 16572 31634 16584
rect 31956 16581 31984 16612
rect 32125 16609 32137 16643
rect 32171 16640 32183 16643
rect 32306 16640 32312 16652
rect 32171 16612 32312 16640
rect 32171 16609 32183 16612
rect 32125 16603 32183 16609
rect 32306 16600 32312 16612
rect 32364 16600 32370 16652
rect 36722 16600 36728 16652
rect 36780 16640 36786 16652
rect 36817 16643 36875 16649
rect 36817 16640 36829 16643
rect 36780 16612 36829 16640
rect 36780 16600 36786 16612
rect 36817 16609 36829 16612
rect 36863 16640 36875 16643
rect 37918 16640 37924 16652
rect 36863 16612 37924 16640
rect 36863 16609 36875 16612
rect 36817 16603 36875 16609
rect 37918 16600 37924 16612
rect 37976 16600 37982 16652
rect 39114 16600 39120 16652
rect 39172 16640 39178 16652
rect 40236 16649 40264 16680
rect 39209 16643 39267 16649
rect 39209 16640 39221 16643
rect 39172 16612 39221 16640
rect 39172 16600 39178 16612
rect 39209 16609 39221 16612
rect 39255 16609 39267 16643
rect 39209 16603 39267 16609
rect 40221 16643 40279 16649
rect 40221 16609 40233 16643
rect 40267 16609 40279 16643
rect 40586 16640 40592 16652
rect 40547 16612 40592 16640
rect 40221 16603 40279 16609
rect 40586 16600 40592 16612
rect 40644 16600 40650 16652
rect 51994 16600 52000 16652
rect 52052 16640 52058 16652
rect 56045 16643 56103 16649
rect 56045 16640 56057 16643
rect 52052 16612 56057 16640
rect 52052 16600 52058 16612
rect 56045 16609 56057 16612
rect 56091 16609 56103 16643
rect 56045 16603 56103 16609
rect 56413 16643 56471 16649
rect 56413 16609 56425 16643
rect 56459 16640 56471 16643
rect 56870 16640 56876 16652
rect 56459 16612 56732 16640
rect 56831 16612 56876 16640
rect 56459 16609 56471 16612
rect 56413 16603 56471 16609
rect 31849 16575 31907 16581
rect 31849 16572 31861 16575
rect 31628 16544 31861 16572
rect 31628 16532 31634 16544
rect 31849 16541 31861 16544
rect 31895 16541 31907 16575
rect 31849 16535 31907 16541
rect 31941 16575 31999 16581
rect 31941 16541 31953 16575
rect 31987 16541 31999 16575
rect 31941 16535 31999 16541
rect 32030 16532 32036 16584
rect 32088 16572 32094 16584
rect 32217 16575 32275 16581
rect 32217 16572 32229 16575
rect 32088 16544 32229 16572
rect 32088 16532 32094 16544
rect 32217 16541 32229 16544
rect 32263 16541 32275 16575
rect 32217 16535 32275 16541
rect 36170 16532 36176 16584
rect 36228 16572 36234 16584
rect 36633 16575 36691 16581
rect 36633 16572 36645 16575
rect 36228 16544 36645 16572
rect 36228 16532 36234 16544
rect 36633 16541 36645 16544
rect 36679 16541 36691 16575
rect 36633 16535 36691 16541
rect 39025 16575 39083 16581
rect 39025 16541 39037 16575
rect 39071 16572 39083 16575
rect 39666 16572 39672 16584
rect 39071 16544 39672 16572
rect 39071 16541 39083 16544
rect 39025 16535 39083 16541
rect 39666 16532 39672 16544
rect 39724 16532 39730 16584
rect 40313 16575 40371 16581
rect 40313 16541 40325 16575
rect 40359 16572 40371 16575
rect 42426 16572 42432 16584
rect 40359 16544 42432 16572
rect 40359 16541 40371 16544
rect 40313 16535 40371 16541
rect 42426 16532 42432 16544
rect 42484 16532 42490 16584
rect 56229 16575 56287 16581
rect 56229 16541 56241 16575
rect 56275 16572 56287 16575
rect 56594 16572 56600 16584
rect 56275 16544 56600 16572
rect 56275 16541 56287 16544
rect 56229 16535 56287 16541
rect 56594 16532 56600 16544
rect 56652 16532 56658 16584
rect 56704 16572 56732 16612
rect 56870 16600 56876 16612
rect 56928 16600 56934 16652
rect 57129 16575 57187 16581
rect 57129 16572 57141 16575
rect 56704 16544 57141 16572
rect 57129 16541 57141 16544
rect 57175 16541 57187 16575
rect 57129 16535 57187 16541
rect 30558 16504 30564 16516
rect 29656 16476 30564 16504
rect 30558 16464 30564 16476
rect 30616 16464 30622 16516
rect 32398 16464 32404 16516
rect 32456 16504 32462 16516
rect 32677 16507 32735 16513
rect 32677 16504 32689 16507
rect 32456 16476 32689 16504
rect 32456 16464 32462 16476
rect 32677 16473 32689 16476
rect 32723 16473 32735 16507
rect 32677 16467 32735 16473
rect 32861 16507 32919 16513
rect 32861 16473 32873 16507
rect 32907 16473 32919 16507
rect 32861 16467 32919 16473
rect 40681 16507 40739 16513
rect 40681 16473 40693 16507
rect 40727 16504 40739 16507
rect 40862 16504 40868 16516
rect 40727 16476 40868 16504
rect 40727 16473 40739 16476
rect 40681 16467 40739 16473
rect 30742 16436 30748 16448
rect 28966 16408 30748 16436
rect 28077 16399 28135 16405
rect 30742 16396 30748 16408
rect 30800 16436 30806 16448
rect 31205 16439 31263 16445
rect 31205 16436 31217 16439
rect 30800 16408 31217 16436
rect 30800 16396 30806 16408
rect 31205 16405 31217 16408
rect 31251 16436 31263 16439
rect 32876 16436 32904 16467
rect 40862 16464 40868 16476
rect 40920 16504 40926 16516
rect 56042 16504 56048 16516
rect 40920 16476 56048 16504
rect 40920 16464 40926 16476
rect 56042 16464 56048 16476
rect 56100 16464 56106 16516
rect 36262 16436 36268 16448
rect 31251 16408 32904 16436
rect 36223 16408 36268 16436
rect 31251 16405 31263 16408
rect 31205 16399 31263 16405
rect 36262 16396 36268 16408
rect 36320 16396 36326 16448
rect 36725 16439 36783 16445
rect 36725 16405 36737 16439
rect 36771 16436 36783 16439
rect 36814 16436 36820 16448
rect 36771 16408 36820 16436
rect 36771 16405 36783 16408
rect 36725 16399 36783 16405
rect 36814 16396 36820 16408
rect 36872 16396 36878 16448
rect 56962 16396 56968 16448
rect 57020 16436 57026 16448
rect 58253 16439 58311 16445
rect 58253 16436 58265 16439
rect 57020 16408 58265 16436
rect 57020 16396 57026 16408
rect 58253 16405 58265 16408
rect 58299 16405 58311 16439
rect 58253 16399 58311 16405
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 16758 16232 16764 16244
rect 12584 16204 16764 16232
rect 12584 16192 12590 16204
rect 16758 16192 16764 16204
rect 16816 16192 16822 16244
rect 16945 16235 17003 16241
rect 16945 16201 16957 16235
rect 16991 16232 17003 16235
rect 17402 16232 17408 16244
rect 16991 16204 17408 16232
rect 16991 16201 17003 16204
rect 16945 16195 17003 16201
rect 17402 16192 17408 16204
rect 17460 16192 17466 16244
rect 17865 16235 17923 16241
rect 17865 16201 17877 16235
rect 17911 16232 17923 16235
rect 18966 16232 18972 16244
rect 17911 16204 18972 16232
rect 17911 16201 17923 16204
rect 17865 16195 17923 16201
rect 18966 16192 18972 16204
rect 19024 16192 19030 16244
rect 19058 16192 19064 16244
rect 19116 16192 19122 16244
rect 22646 16232 22652 16244
rect 19168 16204 22652 16232
rect 15933 16167 15991 16173
rect 15933 16133 15945 16167
rect 15979 16164 15991 16167
rect 16574 16164 16580 16176
rect 15979 16136 16580 16164
rect 15979 16133 15991 16136
rect 15933 16127 15991 16133
rect 16574 16124 16580 16136
rect 16632 16164 16638 16176
rect 17494 16164 17500 16176
rect 16632 16136 16804 16164
rect 16632 16124 16638 16136
rect 1581 16099 1639 16105
rect 1581 16065 1593 16099
rect 1627 16096 1639 16099
rect 2682 16096 2688 16108
rect 1627 16068 2688 16096
rect 1627 16065 1639 16068
rect 1581 16059 1639 16065
rect 2682 16056 2688 16068
rect 2740 16056 2746 16108
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16206 16096 16212 16108
rect 16163 16068 16212 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 1762 16028 1768 16040
rect 1723 16000 1768 16028
rect 1762 15988 1768 16000
rect 1820 15988 1826 16040
rect 16132 15960 16160 16059
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 16776 16028 16804 16136
rect 17144 16136 17500 16164
rect 16850 16056 16856 16108
rect 16908 16096 16914 16108
rect 17144 16105 17172 16136
rect 17494 16124 17500 16136
rect 17552 16124 17558 16176
rect 19076 16164 19104 16192
rect 18064 16136 19104 16164
rect 17129 16099 17187 16105
rect 17129 16096 17141 16099
rect 16908 16068 17141 16096
rect 16908 16056 16914 16068
rect 17129 16065 17141 16068
rect 17175 16065 17187 16099
rect 17310 16096 17316 16108
rect 17271 16068 17316 16096
rect 17129 16059 17187 16065
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16096 17463 16099
rect 17954 16096 17960 16108
rect 17451 16068 17960 16096
rect 17451 16065 17463 16068
rect 17405 16059 17463 16065
rect 17954 16056 17960 16068
rect 18012 16056 18018 16108
rect 18064 16105 18092 16136
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16065 18107 16099
rect 18230 16096 18236 16108
rect 18191 16068 18236 16096
rect 18049 16059 18107 16065
rect 18230 16056 18236 16068
rect 18288 16056 18294 16108
rect 18782 16096 18788 16108
rect 18743 16068 18788 16096
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 18874 16056 18880 16108
rect 18932 16096 18938 16108
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 18932 16068 19073 16096
rect 18932 16056 18938 16068
rect 19061 16065 19073 16068
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 17218 16028 17224 16040
rect 16776 16000 17224 16028
rect 17218 15988 17224 16000
rect 17276 15988 17282 16040
rect 17586 15988 17592 16040
rect 17644 16028 17650 16040
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 17644 16000 18337 16028
rect 17644 15988 17650 16000
rect 18325 15997 18337 16000
rect 18371 15997 18383 16031
rect 19168 16028 19196 16204
rect 22646 16192 22652 16204
rect 22704 16192 22710 16244
rect 23845 16235 23903 16241
rect 23845 16201 23857 16235
rect 23891 16232 23903 16235
rect 26878 16232 26884 16244
rect 23891 16204 26884 16232
rect 23891 16201 23903 16204
rect 23845 16195 23903 16201
rect 26878 16192 26884 16204
rect 26936 16192 26942 16244
rect 31297 16235 31355 16241
rect 31297 16232 31309 16235
rect 27172 16204 31309 16232
rect 21361 16167 21419 16173
rect 21361 16164 21373 16167
rect 20364 16136 21373 16164
rect 19978 16056 19984 16108
rect 20036 16096 20042 16108
rect 20364 16105 20392 16136
rect 21361 16133 21373 16136
rect 21407 16164 21419 16167
rect 22732 16167 22790 16173
rect 21407 16136 22692 16164
rect 21407 16133 21419 16136
rect 21361 16127 21419 16133
rect 20349 16099 20407 16105
rect 20349 16096 20361 16099
rect 20036 16068 20361 16096
rect 20036 16056 20042 16068
rect 20349 16065 20361 16068
rect 20395 16065 20407 16099
rect 21174 16096 21180 16108
rect 21135 16068 21180 16096
rect 20349 16059 20407 16065
rect 21174 16056 21180 16068
rect 21232 16056 21238 16108
rect 21450 16096 21456 16108
rect 21411 16068 21456 16096
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 22664 16096 22692 16136
rect 22732 16133 22744 16167
rect 22778 16164 22790 16167
rect 24854 16164 24860 16176
rect 22778 16136 24860 16164
rect 22778 16133 22790 16136
rect 22732 16127 22790 16133
rect 24854 16124 24860 16136
rect 24912 16124 24918 16176
rect 24305 16099 24363 16105
rect 22664 16068 23888 16096
rect 19334 16028 19340 16040
rect 18325 15991 18383 15997
rect 18432 16000 19196 16028
rect 19295 16000 19340 16028
rect 18432 15960 18460 16000
rect 19334 15988 19340 16000
rect 19392 15988 19398 16040
rect 20441 16031 20499 16037
rect 20441 16028 20453 16031
rect 19444 16000 20453 16028
rect 18874 15960 18880 15972
rect 16132 15932 18460 15960
rect 18835 15932 18880 15960
rect 18874 15920 18880 15932
rect 18932 15960 18938 15972
rect 19242 15960 19248 15972
rect 18932 15932 19248 15960
rect 18932 15920 18938 15932
rect 19242 15920 19248 15932
rect 19300 15920 19306 15972
rect 15746 15852 15752 15904
rect 15804 15892 15810 15904
rect 16301 15895 16359 15901
rect 16301 15892 16313 15895
rect 15804 15864 16313 15892
rect 15804 15852 15810 15864
rect 16301 15861 16313 15864
rect 16347 15861 16359 15895
rect 16301 15855 16359 15861
rect 18506 15852 18512 15904
rect 18564 15892 18570 15904
rect 19444 15892 19472 16000
rect 20441 15997 20453 16000
rect 20487 16028 20499 16031
rect 21468 16028 21496 16056
rect 22462 16028 22468 16040
rect 20487 16000 21496 16028
rect 22423 16000 22468 16028
rect 20487 15997 20499 16000
rect 20441 15991 20499 15997
rect 22462 15988 22468 16000
rect 22520 15988 22526 16040
rect 23860 16028 23888 16068
rect 24305 16065 24317 16099
rect 24351 16096 24363 16099
rect 24578 16096 24584 16108
rect 24351 16068 24584 16096
rect 24351 16065 24363 16068
rect 24305 16059 24363 16065
rect 24578 16056 24584 16068
rect 24636 16056 24642 16108
rect 24946 16056 24952 16108
rect 25004 16096 25010 16108
rect 27172 16105 27200 16204
rect 31297 16201 31309 16204
rect 31343 16201 31355 16235
rect 31297 16195 31355 16201
rect 32582 16192 32588 16244
rect 32640 16232 32646 16244
rect 33962 16232 33968 16244
rect 32640 16204 33968 16232
rect 32640 16192 32646 16204
rect 33962 16192 33968 16204
rect 34020 16192 34026 16244
rect 34054 16192 34060 16244
rect 34112 16232 34118 16244
rect 34149 16235 34207 16241
rect 34149 16232 34161 16235
rect 34112 16204 34161 16232
rect 34112 16192 34118 16204
rect 34149 16201 34161 16204
rect 34195 16201 34207 16235
rect 34149 16195 34207 16201
rect 34514 16192 34520 16244
rect 34572 16232 34578 16244
rect 34572 16204 55214 16232
rect 34572 16192 34578 16204
rect 29546 16124 29552 16176
rect 29604 16164 29610 16176
rect 30162 16167 30220 16173
rect 30162 16164 30174 16167
rect 29604 16136 30174 16164
rect 29604 16124 29610 16136
rect 30162 16133 30174 16136
rect 30208 16133 30220 16167
rect 40494 16164 40500 16176
rect 30162 16127 30220 16133
rect 35452 16136 40500 16164
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 25004 16068 27169 16096
rect 25004 16056 25010 16068
rect 27157 16065 27169 16068
rect 27203 16065 27215 16099
rect 27157 16059 27215 16065
rect 28902 16056 28908 16108
rect 28960 16096 28966 16108
rect 29917 16099 29975 16105
rect 29917 16096 29929 16099
rect 28960 16068 29929 16096
rect 28960 16056 28966 16068
rect 29917 16065 29929 16068
rect 29963 16065 29975 16099
rect 29917 16059 29975 16065
rect 32493 16099 32551 16105
rect 32493 16065 32505 16099
rect 32539 16096 32551 16099
rect 32766 16096 32772 16108
rect 32539 16068 32772 16096
rect 32539 16065 32551 16068
rect 32493 16059 32551 16065
rect 32766 16056 32772 16068
rect 32824 16056 32830 16108
rect 35452 16105 35480 16136
rect 35437 16099 35495 16105
rect 35437 16065 35449 16099
rect 35483 16065 35495 16099
rect 35437 16059 35495 16065
rect 35704 16099 35762 16105
rect 35704 16065 35716 16099
rect 35750 16096 35762 16099
rect 36262 16096 36268 16108
rect 35750 16068 36268 16096
rect 35750 16065 35762 16068
rect 35704 16059 35762 16065
rect 36262 16056 36268 16068
rect 36320 16056 36326 16108
rect 39500 16105 39528 16136
rect 40494 16124 40500 16136
rect 40552 16164 40558 16176
rect 48130 16164 48136 16176
rect 40552 16136 48136 16164
rect 40552 16124 40558 16136
rect 48130 16124 48136 16136
rect 48188 16124 48194 16176
rect 39758 16105 39764 16108
rect 39485 16099 39543 16105
rect 39485 16065 39497 16099
rect 39531 16065 39543 16099
rect 39752 16096 39764 16105
rect 39719 16068 39764 16096
rect 39485 16059 39543 16065
rect 39752 16059 39764 16068
rect 39758 16056 39764 16059
rect 39816 16056 39822 16108
rect 55186 16096 55214 16204
rect 56594 16192 56600 16244
rect 56652 16232 56658 16244
rect 57241 16235 57299 16241
rect 57241 16232 57253 16235
rect 56652 16204 57253 16232
rect 56652 16192 56658 16204
rect 57241 16201 57253 16204
rect 57287 16201 57299 16235
rect 57241 16195 57299 16201
rect 56134 16124 56140 16176
rect 56192 16164 56198 16176
rect 56962 16164 56968 16176
rect 56192 16136 56824 16164
rect 56923 16136 56968 16164
rect 56192 16124 56198 16136
rect 56689 16099 56747 16105
rect 56689 16096 56701 16099
rect 55186 16068 56701 16096
rect 56689 16065 56701 16068
rect 56735 16065 56747 16099
rect 56796 16096 56824 16136
rect 56962 16124 56968 16136
rect 57020 16124 57026 16176
rect 56873 16099 56931 16105
rect 56873 16096 56885 16099
rect 56796 16068 56885 16096
rect 56689 16059 56747 16065
rect 56873 16065 56885 16068
rect 56919 16065 56931 16099
rect 56873 16059 56931 16065
rect 57057 16099 57115 16105
rect 57057 16065 57069 16099
rect 57103 16096 57115 16099
rect 58066 16096 58072 16108
rect 57103 16068 58072 16096
rect 57103 16065 57115 16068
rect 57057 16059 57115 16065
rect 58066 16056 58072 16068
rect 58124 16056 58130 16108
rect 27062 16028 27068 16040
rect 23860 16000 27068 16028
rect 27062 15988 27068 16000
rect 27120 15988 27126 16040
rect 28460 16000 28994 16028
rect 26142 15920 26148 15972
rect 26200 15960 26206 15972
rect 28353 15963 28411 15969
rect 28353 15960 28365 15963
rect 26200 15932 28365 15960
rect 26200 15920 26206 15932
rect 28353 15929 28365 15932
rect 28399 15929 28411 15963
rect 28353 15923 28411 15929
rect 20714 15892 20720 15904
rect 18564 15864 19472 15892
rect 20675 15864 20720 15892
rect 18564 15852 18570 15864
rect 20714 15852 20720 15864
rect 20772 15852 20778 15904
rect 21177 15895 21235 15901
rect 21177 15861 21189 15895
rect 21223 15892 21235 15895
rect 23474 15892 23480 15904
rect 21223 15864 23480 15892
rect 21223 15861 21235 15864
rect 21177 15855 21235 15861
rect 23474 15852 23480 15864
rect 23532 15852 23538 15904
rect 24118 15852 24124 15904
rect 24176 15892 24182 15904
rect 25501 15895 25559 15901
rect 25501 15892 25513 15895
rect 24176 15864 25513 15892
rect 24176 15852 24182 15864
rect 25501 15861 25513 15864
rect 25547 15861 25559 15895
rect 25501 15855 25559 15861
rect 25958 15852 25964 15904
rect 26016 15892 26022 15904
rect 28460 15892 28488 16000
rect 26016 15864 28488 15892
rect 28966 15892 28994 16000
rect 31018 15988 31024 16040
rect 31076 16028 31082 16040
rect 32677 16031 32735 16037
rect 32677 16028 32689 16031
rect 31076 16000 32689 16028
rect 31076 15988 31082 16000
rect 32677 15997 32689 16000
rect 32723 15997 32735 16031
rect 34238 16028 34244 16040
rect 34199 16000 34244 16028
rect 32677 15991 32735 15997
rect 34238 15988 34244 16000
rect 34296 15988 34302 16040
rect 34333 16031 34391 16037
rect 34333 15997 34345 16031
rect 34379 15997 34391 16031
rect 34333 15991 34391 15997
rect 34348 15960 34376 15991
rect 34698 15960 34704 15972
rect 33060 15932 34704 15960
rect 33060 15892 33088 15932
rect 34698 15920 34704 15932
rect 34756 15920 34762 15972
rect 40862 15960 40868 15972
rect 40823 15932 40868 15960
rect 40862 15920 40868 15932
rect 40920 15920 40926 15972
rect 28966 15864 33088 15892
rect 26016 15852 26022 15864
rect 33134 15852 33140 15904
rect 33192 15892 33198 15904
rect 33781 15895 33839 15901
rect 33781 15892 33793 15895
rect 33192 15864 33793 15892
rect 33192 15852 33198 15864
rect 33781 15861 33793 15864
rect 33827 15861 33839 15895
rect 36814 15892 36820 15904
rect 36775 15864 36820 15892
rect 33781 15855 33839 15861
rect 36814 15852 36820 15864
rect 36872 15852 36878 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 18693 15691 18751 15697
rect 18693 15657 18705 15691
rect 18739 15688 18751 15691
rect 19797 15691 19855 15697
rect 19797 15688 19809 15691
rect 18739 15660 19809 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 19797 15657 19809 15660
rect 19843 15688 19855 15691
rect 23290 15688 23296 15700
rect 19843 15660 23296 15688
rect 19843 15657 19855 15660
rect 19797 15651 19855 15657
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 25314 15688 25320 15700
rect 23400 15660 25320 15688
rect 17865 15623 17923 15629
rect 17865 15589 17877 15623
rect 17911 15620 17923 15623
rect 21726 15620 21732 15632
rect 17911 15592 21732 15620
rect 17911 15589 17923 15592
rect 17865 15583 17923 15589
rect 21726 15580 21732 15592
rect 21784 15580 21790 15632
rect 22554 15580 22560 15632
rect 22612 15620 22618 15632
rect 23017 15623 23075 15629
rect 23017 15620 23029 15623
rect 22612 15592 23029 15620
rect 22612 15580 22618 15592
rect 23017 15589 23029 15592
rect 23063 15620 23075 15623
rect 23400 15620 23428 15660
rect 25314 15648 25320 15660
rect 25372 15648 25378 15700
rect 29454 15648 29460 15700
rect 29512 15688 29518 15700
rect 48130 15688 48136 15700
rect 29512 15660 41414 15688
rect 48091 15660 48136 15688
rect 29512 15648 29518 15660
rect 23063 15592 23428 15620
rect 23063 15589 23075 15592
rect 23017 15583 23075 15589
rect 34698 15580 34704 15632
rect 34756 15620 34762 15632
rect 36722 15620 36728 15632
rect 34756 15592 36728 15620
rect 34756 15580 34762 15592
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 19334 15552 19340 15564
rect 11296 15524 19340 15552
rect 11296 15512 11302 15524
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15552 19487 15555
rect 21174 15552 21180 15564
rect 19475 15524 21180 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 21174 15512 21180 15524
rect 21232 15512 21238 15564
rect 22462 15512 22468 15564
rect 22520 15552 22526 15564
rect 24581 15555 24639 15561
rect 24581 15552 24593 15555
rect 22520 15524 24593 15552
rect 22520 15512 22526 15524
rect 24581 15521 24593 15524
rect 24627 15521 24639 15555
rect 24581 15515 24639 15521
rect 26418 15512 26424 15564
rect 26476 15552 26482 15564
rect 30837 15555 30895 15561
rect 30837 15552 30849 15555
rect 26476 15524 30849 15552
rect 26476 15512 26482 15524
rect 30837 15521 30849 15524
rect 30883 15521 30895 15555
rect 30837 15515 30895 15521
rect 34241 15555 34299 15561
rect 34241 15521 34253 15555
rect 34287 15552 34299 15555
rect 34790 15552 34796 15564
rect 34287 15524 34796 15552
rect 34287 15521 34299 15524
rect 34241 15515 34299 15521
rect 34790 15512 34796 15524
rect 34848 15512 34854 15564
rect 35452 15561 35480 15592
rect 36722 15580 36728 15592
rect 36780 15580 36786 15632
rect 35437 15555 35495 15561
rect 35437 15521 35449 15555
rect 35483 15521 35495 15555
rect 41386 15552 41414 15660
rect 48130 15648 48136 15660
rect 48188 15648 48194 15700
rect 58253 15555 58311 15561
rect 58253 15552 58265 15555
rect 41386 15524 58265 15552
rect 35437 15515 35495 15521
rect 58253 15521 58265 15524
rect 58299 15521 58311 15555
rect 58253 15515 58311 15521
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15484 1639 15487
rect 13998 15484 14004 15496
rect 1627 15456 14004 15484
rect 1627 15453 1639 15456
rect 1581 15447 1639 15453
rect 13998 15444 14004 15456
rect 14056 15444 14062 15496
rect 15105 15487 15163 15493
rect 15105 15453 15117 15487
rect 15151 15484 15163 15487
rect 15470 15484 15476 15496
rect 15151 15456 15476 15484
rect 15151 15453 15163 15456
rect 15105 15447 15163 15453
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 17678 15444 17684 15496
rect 17736 15484 17742 15496
rect 17865 15487 17923 15493
rect 17865 15484 17877 15487
rect 17736 15456 17877 15484
rect 17736 15444 17742 15456
rect 17865 15453 17877 15456
rect 17911 15453 17923 15487
rect 17865 15447 17923 15453
rect 18049 15487 18107 15493
rect 18049 15453 18061 15487
rect 18095 15484 18107 15487
rect 19518 15484 19524 15496
rect 18095 15456 19524 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 19518 15444 19524 15456
rect 19576 15444 19582 15496
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15484 19671 15487
rect 19978 15484 19984 15496
rect 19659 15456 19984 15484
rect 19659 15453 19671 15456
rect 19613 15447 19671 15453
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 20257 15487 20315 15493
rect 20257 15453 20269 15487
rect 20303 15484 20315 15487
rect 20714 15484 20720 15496
rect 20303 15456 20720 15484
rect 20303 15453 20315 15456
rect 20257 15447 20315 15453
rect 20714 15444 20720 15456
rect 20772 15444 20778 15496
rect 23566 15484 23572 15496
rect 23527 15456 23572 15484
rect 23566 15444 23572 15456
rect 23624 15444 23630 15496
rect 26878 15484 26884 15496
rect 26839 15456 26884 15484
rect 26878 15444 26884 15456
rect 26936 15444 26942 15496
rect 29730 15484 29736 15496
rect 29691 15456 29736 15484
rect 29730 15444 29736 15456
rect 29788 15444 29794 15496
rect 29914 15444 29920 15496
rect 29972 15484 29978 15496
rect 32493 15487 32551 15493
rect 32493 15484 32505 15487
rect 29972 15456 32505 15484
rect 29972 15444 29978 15456
rect 32493 15453 32505 15456
rect 32539 15484 32551 15487
rect 39942 15484 39948 15496
rect 32539 15456 39948 15484
rect 32539 15453 32551 15456
rect 32493 15447 32551 15453
rect 39942 15444 39948 15456
rect 40000 15484 40006 15496
rect 40000 15456 41414 15484
rect 40000 15444 40006 15456
rect 1854 15416 1860 15428
rect 1815 15388 1860 15416
rect 1854 15376 1860 15388
rect 1912 15376 1918 15428
rect 18506 15416 18512 15428
rect 18467 15388 18512 15416
rect 18506 15376 18512 15388
rect 18564 15376 18570 15428
rect 18725 15419 18783 15425
rect 18725 15385 18737 15419
rect 18771 15416 18783 15419
rect 23385 15419 23443 15425
rect 23385 15416 23397 15419
rect 18771 15388 23397 15416
rect 18771 15385 18783 15388
rect 18725 15379 18783 15385
rect 23385 15385 23397 15388
rect 23431 15416 23443 15419
rect 23842 15416 23848 15428
rect 23431 15388 23848 15416
rect 23431 15385 23443 15388
rect 23385 15379 23443 15385
rect 23842 15376 23848 15388
rect 23900 15376 23906 15428
rect 24848 15419 24906 15425
rect 24848 15385 24860 15419
rect 24894 15416 24906 15419
rect 25682 15416 25688 15428
rect 24894 15388 25688 15416
rect 24894 15385 24906 15388
rect 24848 15379 24906 15385
rect 25682 15376 25688 15388
rect 25740 15376 25746 15428
rect 29270 15376 29276 15428
rect 29328 15416 29334 15428
rect 30098 15416 30104 15428
rect 29328 15388 30104 15416
rect 29328 15376 29334 15388
rect 30098 15376 30104 15388
rect 30156 15376 30162 15428
rect 35253 15419 35311 15425
rect 35253 15385 35265 15419
rect 35299 15416 35311 15419
rect 35802 15416 35808 15428
rect 35299 15388 35808 15416
rect 35299 15385 35311 15388
rect 35253 15379 35311 15385
rect 35802 15376 35808 15388
rect 35860 15376 35866 15428
rect 41386 15416 41414 15456
rect 56042 15444 56048 15496
rect 56100 15484 56106 15496
rect 56965 15487 57023 15493
rect 56965 15484 56977 15487
rect 56100 15456 56977 15484
rect 56100 15444 56106 15456
rect 56965 15453 56977 15456
rect 57011 15453 57023 15487
rect 57974 15484 57980 15496
rect 57935 15456 57980 15484
rect 56965 15447 57023 15453
rect 57974 15444 57980 15456
rect 58032 15444 58038 15496
rect 46842 15416 46848 15428
rect 41386 15388 46848 15416
rect 46842 15376 46848 15388
rect 46900 15376 46906 15428
rect 57238 15416 57244 15428
rect 57199 15388 57244 15416
rect 57238 15376 57244 15388
rect 57296 15376 57302 15428
rect 15102 15308 15108 15360
rect 15160 15348 15166 15360
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 15160 15320 16313 15348
rect 15160 15308 15166 15320
rect 16301 15317 16313 15320
rect 16347 15317 16359 15351
rect 16301 15311 16359 15317
rect 16666 15308 16672 15360
rect 16724 15348 16730 15360
rect 18877 15351 18935 15357
rect 18877 15348 18889 15351
rect 16724 15320 18889 15348
rect 16724 15308 16730 15320
rect 18877 15317 18889 15320
rect 18923 15348 18935 15351
rect 20806 15348 20812 15360
rect 18923 15320 20812 15348
rect 18923 15317 18935 15320
rect 18877 15311 18935 15317
rect 20806 15308 20812 15320
rect 20864 15308 20870 15360
rect 21450 15348 21456 15360
rect 21411 15320 21456 15348
rect 21450 15308 21456 15320
rect 21508 15308 21514 15360
rect 23198 15348 23204 15360
rect 23159 15320 23204 15348
rect 23198 15308 23204 15320
rect 23256 15308 23262 15360
rect 23290 15308 23296 15360
rect 23348 15348 23354 15360
rect 25961 15351 26019 15357
rect 23348 15320 23393 15348
rect 23348 15308 23354 15320
rect 25961 15317 25973 15351
rect 26007 15348 26019 15351
rect 26878 15348 26884 15360
rect 26007 15320 26884 15348
rect 26007 15317 26019 15320
rect 25961 15311 26019 15317
rect 26878 15308 26884 15320
rect 26936 15308 26942 15360
rect 29086 15348 29092 15360
rect 29047 15320 29092 15348
rect 29086 15308 29092 15320
rect 29144 15308 29150 15360
rect 34885 15351 34943 15357
rect 34885 15317 34897 15351
rect 34931 15348 34943 15351
rect 34974 15348 34980 15360
rect 34931 15320 34980 15348
rect 34931 15317 34943 15320
rect 34885 15311 34943 15317
rect 34974 15308 34980 15320
rect 35032 15308 35038 15360
rect 35342 15308 35348 15360
rect 35400 15348 35406 15360
rect 35400 15320 35445 15348
rect 35400 15308 35406 15320
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 14185 15147 14243 15153
rect 14185 15113 14197 15147
rect 14231 15144 14243 15147
rect 14918 15144 14924 15156
rect 14231 15116 14924 15144
rect 14231 15113 14243 15116
rect 14185 15107 14243 15113
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 19334 15104 19340 15156
rect 19392 15144 19398 15156
rect 32398 15144 32404 15156
rect 19392 15116 32404 15144
rect 19392 15104 19398 15116
rect 32398 15104 32404 15116
rect 32456 15104 32462 15156
rect 18049 15079 18107 15085
rect 18049 15045 18061 15079
rect 18095 15076 18107 15079
rect 18506 15076 18512 15088
rect 18095 15048 18512 15076
rect 18095 15045 18107 15048
rect 18049 15039 18107 15045
rect 18506 15036 18512 15048
rect 18564 15036 18570 15088
rect 19978 15076 19984 15088
rect 19076 15048 19984 15076
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 15008 1639 15011
rect 16758 15008 16764 15020
rect 1627 14980 16764 15008
rect 1627 14977 1639 14980
rect 1581 14971 1639 14977
rect 16758 14968 16764 14980
rect 16816 14968 16822 15020
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 13725 14943 13783 14949
rect 13725 14909 13737 14943
rect 13771 14940 13783 14943
rect 13814 14940 13820 14952
rect 13771 14912 13820 14940
rect 13771 14909 13783 14912
rect 13725 14903 13783 14909
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 14642 14940 14648 14952
rect 14603 14912 14648 14940
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 14918 14940 14924 14952
rect 14879 14912 14924 14940
rect 14918 14900 14924 14912
rect 14976 14900 14982 14952
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 17218 14940 17224 14952
rect 17175 14912 17224 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 17218 14900 17224 14912
rect 17276 14900 17282 14952
rect 19076 14949 19104 15048
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 20248 15079 20306 15085
rect 20248 15045 20260 15079
rect 20294 15076 20306 15079
rect 21450 15076 21456 15088
rect 20294 15048 21456 15076
rect 20294 15045 20306 15048
rect 20248 15039 20306 15045
rect 21450 15036 21456 15048
rect 21508 15036 21514 15088
rect 22732 15079 22790 15085
rect 22732 15045 22744 15079
rect 22778 15076 22790 15079
rect 24118 15076 24124 15088
rect 22778 15048 24124 15076
rect 22778 15045 22790 15048
rect 22732 15039 22790 15045
rect 24118 15036 24124 15048
rect 24176 15036 24182 15088
rect 26970 15076 26976 15088
rect 24228 15048 26976 15076
rect 19153 15011 19211 15017
rect 19153 14977 19165 15011
rect 19199 15008 19211 15011
rect 19334 15008 19340 15020
rect 19199 14980 19340 15008
rect 19199 14977 19211 14980
rect 19153 14971 19211 14977
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 19061 14943 19119 14949
rect 19061 14909 19073 14943
rect 19107 14909 19119 14943
rect 19061 14903 19119 14909
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 19981 14943 20039 14949
rect 19981 14940 19993 14943
rect 19484 14912 19993 14940
rect 19484 14900 19490 14912
rect 19981 14909 19993 14912
rect 20027 14909 20039 14943
rect 19981 14903 20039 14909
rect 22002 14900 22008 14952
rect 22060 14940 22066 14952
rect 22462 14940 22468 14952
rect 22060 14912 22468 14940
rect 22060 14900 22066 14912
rect 22462 14900 22468 14912
rect 22520 14900 22526 14952
rect 24228 14940 24256 15048
rect 26970 15036 26976 15048
rect 27028 15076 27034 15088
rect 30190 15076 30196 15088
rect 27028 15048 30196 15076
rect 27028 15036 27034 15048
rect 30190 15036 30196 15048
rect 30248 15036 30254 15088
rect 30300 15048 34744 15076
rect 30300 15020 30328 15048
rect 24305 15011 24363 15017
rect 24305 14977 24317 15011
rect 24351 15008 24363 15011
rect 26326 15008 26332 15020
rect 24351 14980 26332 15008
rect 24351 14977 24363 14980
rect 24305 14971 24363 14977
rect 26326 14968 26332 14980
rect 26384 14968 26390 15020
rect 27154 15008 27160 15020
rect 27115 14980 27160 15008
rect 27154 14968 27160 14980
rect 27212 14968 27218 15020
rect 29822 14968 29828 15020
rect 29880 15008 29886 15020
rect 30282 15008 30288 15020
rect 29880 14980 30288 15008
rect 29880 14968 29886 14980
rect 30282 14968 30288 14980
rect 30340 14968 30346 15020
rect 30552 15011 30610 15017
rect 30552 14977 30564 15011
rect 30598 15008 30610 15011
rect 31110 15008 31116 15020
rect 30598 14980 31116 15008
rect 30598 14977 30610 14980
rect 30552 14971 30610 14977
rect 31110 14968 31116 14980
rect 31168 14968 31174 15020
rect 32876 15017 32904 15048
rect 33134 15017 33140 15020
rect 32861 15011 32919 15017
rect 32861 14977 32873 15011
rect 32907 14977 32919 15011
rect 33128 15008 33140 15017
rect 33095 14980 33140 15008
rect 32861 14971 32919 14977
rect 33128 14971 33140 14980
rect 33134 14968 33140 14971
rect 33192 14968 33198 15020
rect 34716 15017 34744 15048
rect 34701 15011 34759 15017
rect 34701 14977 34713 15011
rect 34747 15008 34759 15011
rect 34790 15008 34796 15020
rect 34747 14980 34796 15008
rect 34747 14977 34759 14980
rect 34701 14971 34759 14977
rect 34790 14968 34796 14980
rect 34848 14968 34854 15020
rect 34974 15017 34980 15020
rect 34968 15008 34980 15017
rect 34935 14980 34980 15008
rect 34968 14971 34980 14980
rect 34974 14968 34980 14971
rect 35032 14968 35038 15020
rect 23768 14912 24256 14940
rect 13170 14832 13176 14884
rect 13228 14872 13234 14884
rect 14001 14875 14059 14881
rect 14001 14872 14013 14875
rect 13228 14844 14013 14872
rect 13228 14832 13234 14844
rect 14001 14841 14013 14844
rect 14047 14841 14059 14875
rect 14001 14835 14059 14841
rect 17497 14875 17555 14881
rect 17497 14841 17509 14875
rect 17543 14872 17555 14875
rect 18138 14872 18144 14884
rect 17543 14844 18144 14872
rect 17543 14841 17555 14844
rect 17497 14835 17555 14841
rect 18138 14832 18144 14844
rect 18196 14832 18202 14884
rect 18414 14872 18420 14884
rect 18375 14844 18420 14872
rect 18414 14832 18420 14844
rect 18472 14832 18478 14884
rect 18509 14875 18567 14881
rect 18509 14841 18521 14875
rect 18555 14872 18567 14875
rect 18555 14844 20024 14872
rect 18555 14841 18567 14844
rect 18509 14835 18567 14841
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 14826 14804 14832 14816
rect 13872 14776 14832 14804
rect 13872 14764 13878 14776
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 16206 14804 16212 14816
rect 16167 14776 16212 14804
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 16574 14764 16580 14816
rect 16632 14804 16638 14816
rect 17589 14807 17647 14813
rect 17589 14804 17601 14807
rect 16632 14776 17601 14804
rect 16632 14764 16638 14776
rect 17589 14773 17601 14776
rect 17635 14773 17647 14807
rect 17589 14767 17647 14773
rect 19150 14764 19156 14816
rect 19208 14804 19214 14816
rect 19429 14807 19487 14813
rect 19429 14804 19441 14807
rect 19208 14776 19441 14804
rect 19208 14764 19214 14776
rect 19429 14773 19441 14776
rect 19475 14773 19487 14807
rect 19996 14804 20024 14844
rect 21082 14804 21088 14816
rect 19996 14776 21088 14804
rect 19429 14767 19487 14773
rect 21082 14764 21088 14776
rect 21140 14764 21146 14816
rect 21358 14804 21364 14816
rect 21319 14776 21364 14804
rect 21358 14764 21364 14776
rect 21416 14764 21422 14816
rect 21450 14764 21456 14816
rect 21508 14804 21514 14816
rect 23768 14804 23796 14912
rect 24762 14900 24768 14952
rect 24820 14940 24826 14952
rect 28261 14943 28319 14949
rect 28261 14940 28273 14943
rect 24820 14912 28273 14940
rect 24820 14900 24826 14912
rect 28261 14909 28273 14912
rect 28307 14909 28319 14943
rect 28261 14903 28319 14909
rect 23845 14875 23903 14881
rect 23845 14841 23857 14875
rect 23891 14872 23903 14875
rect 24946 14872 24952 14884
rect 23891 14844 24952 14872
rect 23891 14841 23903 14844
rect 23845 14835 23903 14841
rect 24946 14832 24952 14844
rect 25004 14832 25010 14884
rect 21508 14776 23796 14804
rect 21508 14764 21514 14776
rect 24670 14764 24676 14816
rect 24728 14804 24734 14816
rect 25501 14807 25559 14813
rect 25501 14804 25513 14807
rect 24728 14776 25513 14804
rect 24728 14764 24734 14776
rect 25501 14773 25513 14776
rect 25547 14773 25559 14807
rect 25501 14767 25559 14773
rect 29730 14764 29736 14816
rect 29788 14804 29794 14816
rect 31665 14807 31723 14813
rect 31665 14804 31677 14807
rect 29788 14776 31677 14804
rect 29788 14764 29794 14776
rect 31665 14773 31677 14776
rect 31711 14804 31723 14807
rect 32490 14804 32496 14816
rect 31711 14776 32496 14804
rect 31711 14773 31723 14776
rect 31665 14767 31723 14773
rect 32490 14764 32496 14776
rect 32548 14764 32554 14816
rect 33778 14764 33784 14816
rect 33836 14804 33842 14816
rect 34238 14804 34244 14816
rect 33836 14776 34244 14804
rect 33836 14764 33842 14776
rect 34238 14764 34244 14776
rect 34296 14764 34302 14816
rect 35342 14764 35348 14816
rect 35400 14804 35406 14816
rect 36081 14807 36139 14813
rect 36081 14804 36093 14807
rect 35400 14776 36093 14804
rect 35400 14764 35406 14776
rect 36081 14773 36093 14776
rect 36127 14773 36139 14807
rect 36081 14767 36139 14773
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 15470 14600 15476 14612
rect 15431 14572 15476 14600
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 18414 14560 18420 14612
rect 18472 14600 18478 14612
rect 22925 14603 22983 14609
rect 22925 14600 22937 14603
rect 18472 14572 22937 14600
rect 18472 14560 18478 14572
rect 22925 14569 22937 14572
rect 22971 14569 22983 14603
rect 22925 14563 22983 14569
rect 23014 14560 23020 14612
rect 23072 14600 23078 14612
rect 30650 14600 30656 14612
rect 23072 14572 30656 14600
rect 23072 14560 23078 14572
rect 30650 14560 30656 14572
rect 30708 14560 30714 14612
rect 31110 14560 31116 14612
rect 31168 14600 31174 14612
rect 31205 14603 31263 14609
rect 31205 14600 31217 14603
rect 31168 14572 31217 14600
rect 31168 14560 31174 14572
rect 31205 14569 31217 14572
rect 31251 14569 31263 14603
rect 31205 14563 31263 14569
rect 31478 14560 31484 14612
rect 31536 14600 31542 14612
rect 36722 14600 36728 14612
rect 31536 14572 36728 14600
rect 31536 14560 31542 14572
rect 36722 14560 36728 14572
rect 36780 14560 36786 14612
rect 58066 14600 58072 14612
rect 58027 14572 58072 14600
rect 58066 14560 58072 14572
rect 58124 14560 58130 14612
rect 21818 14492 21824 14544
rect 21876 14532 21882 14544
rect 30285 14535 30343 14541
rect 21876 14504 30144 14532
rect 21876 14492 21882 14504
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14464 15347 14467
rect 15378 14464 15384 14476
rect 15335 14436 15384 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 15378 14424 15384 14436
rect 15436 14464 15442 14476
rect 17129 14467 17187 14473
rect 17129 14464 17141 14467
rect 15436 14436 17141 14464
rect 15436 14424 15442 14436
rect 17129 14433 17141 14436
rect 17175 14433 17187 14467
rect 17129 14427 17187 14433
rect 24673 14467 24731 14473
rect 24673 14433 24685 14467
rect 24719 14433 24731 14467
rect 29270 14464 29276 14476
rect 24673 14427 24731 14433
rect 24964 14436 29276 14464
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14396 1639 14399
rect 13906 14396 13912 14408
rect 1627 14368 13912 14396
rect 1627 14365 1639 14368
rect 1581 14359 1639 14365
rect 13906 14356 13912 14368
rect 13964 14356 13970 14408
rect 15197 14399 15255 14405
rect 15197 14365 15209 14399
rect 15243 14396 15255 14399
rect 15838 14396 15844 14408
rect 15243 14368 15844 14396
rect 15243 14365 15255 14368
rect 15197 14359 15255 14365
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 16022 14396 16028 14408
rect 15983 14368 16028 14396
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 19426 14356 19432 14408
rect 19484 14396 19490 14408
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 19484 14368 19625 14396
rect 19484 14356 19490 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14396 19947 14399
rect 20346 14396 20352 14408
rect 19935 14368 20352 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 20346 14356 20352 14368
rect 20404 14356 20410 14408
rect 21726 14396 21732 14408
rect 21687 14368 21732 14396
rect 21726 14356 21732 14368
rect 21784 14356 21790 14408
rect 23934 14356 23940 14408
rect 23992 14396 23998 14408
rect 24688 14396 24716 14427
rect 23992 14368 24716 14396
rect 23992 14356 23998 14368
rect 24762 14356 24768 14408
rect 24820 14396 24826 14408
rect 24820 14368 24865 14396
rect 24820 14356 24826 14368
rect 1854 14328 1860 14340
rect 1815 14300 1860 14328
rect 1854 14288 1860 14300
rect 1912 14288 1918 14340
rect 21177 14263 21235 14269
rect 21177 14229 21189 14263
rect 21223 14260 21235 14263
rect 24964 14260 24992 14436
rect 29270 14424 29276 14436
rect 29328 14424 29334 14476
rect 26145 14399 26203 14405
rect 26145 14365 26157 14399
rect 26191 14396 26203 14399
rect 26418 14396 26424 14408
rect 26191 14368 26424 14396
rect 26191 14365 26203 14368
rect 26145 14359 26203 14365
rect 26418 14356 26424 14368
rect 26476 14356 26482 14408
rect 27062 14356 27068 14408
rect 27120 14396 27126 14408
rect 28445 14399 28503 14405
rect 28445 14396 28457 14399
rect 27120 14368 28457 14396
rect 27120 14356 27126 14368
rect 28445 14365 28457 14368
rect 28491 14365 28503 14399
rect 29086 14396 29092 14408
rect 29047 14368 29092 14396
rect 28445 14359 28503 14365
rect 29086 14356 29092 14368
rect 29144 14356 29150 14408
rect 29178 14356 29184 14408
rect 29236 14396 29242 14408
rect 29917 14399 29975 14405
rect 29917 14396 29929 14399
rect 29236 14368 29929 14396
rect 29236 14356 29242 14368
rect 29917 14365 29929 14368
rect 29963 14396 29975 14399
rect 30006 14396 30012 14408
rect 29963 14368 30012 14396
rect 29963 14365 29975 14368
rect 29917 14359 29975 14365
rect 30006 14356 30012 14368
rect 30064 14356 30070 14408
rect 30116 14405 30144 14504
rect 30285 14501 30297 14535
rect 30331 14532 30343 14535
rect 34422 14532 34428 14544
rect 30331 14504 34428 14532
rect 30331 14501 30343 14504
rect 30285 14495 30343 14501
rect 34422 14492 34428 14504
rect 34480 14492 34486 14544
rect 30190 14424 30196 14476
rect 30248 14464 30254 14476
rect 30926 14464 30932 14476
rect 30248 14436 30932 14464
rect 30248 14424 30254 14436
rect 30926 14424 30932 14436
rect 30984 14424 30990 14476
rect 31294 14424 31300 14476
rect 31352 14464 31358 14476
rect 32677 14467 32735 14473
rect 32677 14464 32689 14467
rect 31352 14436 31616 14464
rect 31352 14424 31358 14436
rect 30101 14399 30159 14405
rect 30101 14365 30113 14399
rect 30147 14365 30159 14399
rect 30101 14359 30159 14365
rect 30377 14399 30435 14405
rect 30377 14365 30389 14399
rect 30423 14365 30435 14399
rect 30377 14359 30435 14365
rect 30745 14399 30803 14405
rect 30745 14365 30757 14399
rect 30791 14396 30803 14399
rect 31018 14396 31024 14408
rect 30791 14368 31024 14396
rect 30791 14365 30803 14368
rect 30745 14359 30803 14365
rect 25406 14288 25412 14340
rect 25464 14328 25470 14340
rect 29730 14328 29736 14340
rect 25464 14300 29736 14328
rect 25464 14288 25470 14300
rect 29730 14288 29736 14300
rect 29788 14328 29794 14340
rect 30392 14328 30420 14359
rect 31018 14356 31024 14368
rect 31076 14356 31082 14408
rect 31478 14396 31484 14408
rect 31439 14368 31484 14396
rect 31478 14356 31484 14368
rect 31536 14356 31542 14408
rect 31588 14405 31616 14436
rect 31680 14436 32689 14464
rect 31680 14405 31708 14436
rect 32677 14433 32689 14436
rect 32723 14433 32735 14467
rect 32677 14427 32735 14433
rect 31573 14399 31631 14405
rect 31573 14365 31585 14399
rect 31619 14365 31631 14399
rect 31573 14359 31631 14365
rect 31665 14399 31723 14405
rect 31665 14365 31677 14399
rect 31711 14365 31723 14399
rect 31665 14359 31723 14365
rect 31849 14399 31907 14405
rect 31849 14365 31861 14399
rect 31895 14365 31907 14399
rect 32490 14396 32496 14408
rect 32451 14368 32496 14396
rect 31849 14359 31907 14365
rect 31754 14328 31760 14340
rect 29788 14300 30420 14328
rect 30484 14300 31760 14328
rect 29788 14288 29794 14300
rect 25130 14260 25136 14272
rect 21223 14232 24992 14260
rect 25091 14232 25136 14260
rect 21223 14229 21235 14232
rect 21177 14223 21235 14229
rect 25130 14220 25136 14232
rect 25188 14220 25194 14272
rect 27154 14220 27160 14272
rect 27212 14260 27218 14272
rect 27338 14260 27344 14272
rect 27212 14232 27344 14260
rect 27212 14220 27218 14232
rect 27338 14220 27344 14232
rect 27396 14260 27402 14272
rect 29089 14263 29147 14269
rect 29089 14260 29101 14263
rect 27396 14232 29101 14260
rect 27396 14220 27402 14232
rect 29089 14229 29101 14232
rect 29135 14260 29147 14263
rect 30484 14260 30512 14300
rect 31754 14288 31760 14300
rect 31812 14288 31818 14340
rect 29135 14232 30512 14260
rect 29135 14229 29147 14232
rect 29089 14223 29147 14229
rect 31662 14220 31668 14272
rect 31720 14260 31726 14272
rect 31864 14260 31892 14359
rect 32490 14356 32496 14368
rect 32548 14356 32554 14408
rect 57974 14396 57980 14408
rect 57935 14368 57980 14396
rect 57974 14356 57980 14368
rect 58032 14356 58038 14408
rect 32309 14331 32367 14337
rect 32309 14297 32321 14331
rect 32355 14328 32367 14331
rect 33226 14328 33232 14340
rect 32355 14300 33232 14328
rect 32355 14297 32367 14300
rect 32309 14291 32367 14297
rect 33226 14288 33232 14300
rect 33284 14328 33290 14340
rect 34146 14328 34152 14340
rect 33284 14300 34152 14328
rect 33284 14288 33290 14300
rect 34146 14288 34152 14300
rect 34204 14288 34210 14340
rect 31720 14232 31892 14260
rect 31720 14220 31726 14232
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 14918 14016 14924 14068
rect 14976 14056 14982 14068
rect 15197 14059 15255 14065
rect 15197 14056 15209 14059
rect 14976 14028 15209 14056
rect 14976 14016 14982 14028
rect 15197 14025 15209 14028
rect 15243 14025 15255 14059
rect 15197 14019 15255 14025
rect 15838 14016 15844 14068
rect 15896 14056 15902 14068
rect 20346 14056 20352 14068
rect 15896 14028 19564 14056
rect 20307 14028 20352 14056
rect 15896 14016 15902 14028
rect 19536 13988 19564 14028
rect 20346 14016 20352 14028
rect 20404 14016 20410 14068
rect 22462 14056 22468 14068
rect 22066 14028 22468 14056
rect 22066 13988 22094 14028
rect 22462 14016 22468 14028
rect 22520 14016 22526 14068
rect 23385 14059 23443 14065
rect 23385 14025 23397 14059
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 19076 13960 19334 13988
rect 19536 13960 22094 13988
rect 23400 13988 23428 14019
rect 26878 14016 26884 14068
rect 26936 14056 26942 14068
rect 28537 14059 28595 14065
rect 28537 14056 28549 14059
rect 26936 14028 28549 14056
rect 26936 14016 26942 14028
rect 28537 14025 28549 14028
rect 28583 14025 28595 14059
rect 28537 14019 28595 14025
rect 28626 14016 28632 14068
rect 28684 14056 28690 14068
rect 28684 14028 29408 14056
rect 28684 14016 28690 14028
rect 27246 13988 27252 14000
rect 23400 13960 27108 13988
rect 27159 13960 27252 13988
rect 14001 13923 14059 13929
rect 14001 13889 14013 13923
rect 14047 13920 14059 13923
rect 15930 13920 15936 13932
rect 14047 13892 15936 13920
rect 14047 13889 14059 13892
rect 14001 13883 14059 13889
rect 15930 13880 15936 13892
rect 15988 13880 15994 13932
rect 19076 13920 19104 13960
rect 16868 13892 19104 13920
rect 14642 13812 14648 13864
rect 14700 13852 14706 13864
rect 16868 13861 16896 13892
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 19306 13920 19334 13960
rect 19426 13920 19432 13932
rect 19208 13892 19253 13920
rect 19306 13892 19432 13920
rect 19208 13880 19214 13892
rect 19426 13880 19432 13892
rect 19484 13920 19490 13932
rect 19610 13920 19616 13932
rect 19484 13892 19616 13920
rect 19484 13880 19490 13892
rect 19610 13880 19616 13892
rect 19668 13920 19674 13932
rect 22002 13920 22008 13932
rect 19668 13892 22008 13920
rect 19668 13880 19674 13892
rect 22002 13880 22008 13892
rect 22060 13880 22066 13932
rect 22278 13929 22284 13932
rect 22272 13883 22284 13929
rect 22336 13920 22342 13932
rect 22336 13892 22372 13920
rect 22278 13880 22284 13883
rect 22336 13880 22342 13892
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 24029 13923 24087 13929
rect 24029 13920 24041 13923
rect 23532 13892 24041 13920
rect 23532 13880 23538 13892
rect 24029 13889 24041 13892
rect 24075 13889 24087 13923
rect 24029 13883 24087 13889
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 14700 13824 16865 13852
rect 14700 13812 14706 13824
rect 16853 13821 16865 13824
rect 16899 13821 16911 13855
rect 17126 13852 17132 13864
rect 17087 13824 17132 13852
rect 16853 13815 16911 13821
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 18506 13852 18512 13864
rect 18467 13824 18512 13852
rect 18506 13812 18512 13824
rect 18564 13812 18570 13864
rect 23658 13812 23664 13864
rect 23716 13852 23722 13864
rect 25133 13855 25191 13861
rect 25133 13852 25145 13855
rect 23716 13824 25145 13852
rect 23716 13812 23722 13824
rect 25133 13821 25145 13824
rect 25179 13821 25191 13855
rect 27080 13852 27108 13960
rect 27172 13929 27200 13960
rect 27246 13948 27252 13960
rect 27304 13988 27310 14000
rect 28902 13988 28908 14000
rect 27304 13960 28908 13988
rect 27304 13948 27310 13960
rect 28902 13948 28908 13960
rect 28960 13948 28966 14000
rect 29380 13997 29408 14028
rect 30834 14016 30840 14068
rect 30892 14056 30898 14068
rect 30892 14028 31340 14056
rect 30892 14016 30898 14028
rect 29365 13991 29423 13997
rect 29365 13957 29377 13991
rect 29411 13957 29423 13991
rect 31312 13988 31340 14028
rect 32306 14016 32312 14068
rect 32364 14056 32370 14068
rect 32401 14059 32459 14065
rect 32401 14056 32413 14059
rect 32364 14028 32413 14056
rect 32364 14016 32370 14028
rect 32401 14025 32413 14028
rect 32447 14025 32459 14059
rect 32401 14019 32459 14025
rect 39942 14016 39948 14068
rect 40000 14056 40006 14068
rect 40037 14059 40095 14065
rect 40037 14056 40049 14059
rect 40000 14028 40049 14056
rect 40000 14016 40006 14028
rect 40037 14025 40049 14028
rect 40083 14025 40095 14059
rect 40037 14019 40095 14025
rect 33781 13991 33839 13997
rect 29365 13951 29423 13957
rect 30404 13960 31248 13988
rect 31312 13960 31432 13988
rect 27430 13929 27436 13932
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 27424 13920 27436 13929
rect 27391 13892 27436 13920
rect 27157 13883 27215 13889
rect 27424 13883 27436 13892
rect 27430 13880 27436 13883
rect 27488 13880 27494 13932
rect 30404 13920 30432 13960
rect 28644 13892 30432 13920
rect 30469 13923 30527 13929
rect 27080 13824 27200 13852
rect 25133 13815 25191 13821
rect 17862 13744 17868 13796
rect 17920 13784 17926 13796
rect 21818 13784 21824 13796
rect 17920 13756 21824 13784
rect 17920 13744 17926 13756
rect 21818 13744 21824 13756
rect 21876 13744 21882 13796
rect 17586 13676 17592 13728
rect 17644 13716 17650 13728
rect 21450 13716 21456 13728
rect 17644 13688 21456 13716
rect 17644 13676 17650 13688
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 27172 13716 27200 13824
rect 28644 13784 28672 13892
rect 30469 13889 30481 13923
rect 30515 13920 30527 13923
rect 30515 13892 30880 13920
rect 30515 13889 30527 13892
rect 30469 13883 30527 13889
rect 28718 13812 28724 13864
rect 28776 13852 28782 13864
rect 29457 13855 29515 13861
rect 29457 13852 29469 13855
rect 28776 13824 29469 13852
rect 28776 13812 28782 13824
rect 29457 13821 29469 13824
rect 29503 13821 29515 13855
rect 29457 13815 29515 13821
rect 29641 13855 29699 13861
rect 29641 13821 29653 13855
rect 29687 13821 29699 13855
rect 29641 13815 29699 13821
rect 28092 13756 28672 13784
rect 29656 13784 29684 13815
rect 30006 13812 30012 13864
rect 30064 13852 30070 13864
rect 30742 13852 30748 13864
rect 30064 13824 30748 13852
rect 30064 13812 30070 13824
rect 30742 13812 30748 13824
rect 30800 13812 30806 13864
rect 30852 13852 30880 13892
rect 30926 13880 30932 13932
rect 30984 13920 30990 13932
rect 31220 13920 31248 13960
rect 31404 13929 31432 13960
rect 33781 13957 33793 13991
rect 33827 13988 33839 13991
rect 34146 13988 34152 14000
rect 33827 13960 34152 13988
rect 33827 13957 33839 13960
rect 33781 13951 33839 13957
rect 34146 13948 34152 13960
rect 34204 13948 34210 14000
rect 31297 13923 31355 13929
rect 31297 13920 31309 13923
rect 30984 13892 31029 13920
rect 31220 13892 31309 13920
rect 30984 13880 30990 13892
rect 31297 13889 31309 13892
rect 31343 13889 31355 13923
rect 31297 13883 31355 13889
rect 31389 13923 31447 13929
rect 31389 13889 31401 13923
rect 31435 13920 31447 13923
rect 32122 13920 32128 13932
rect 31435 13892 32128 13920
rect 31435 13889 31447 13892
rect 31389 13883 31447 13889
rect 31312 13852 31340 13883
rect 32122 13880 32128 13892
rect 32180 13920 32186 13932
rect 32309 13923 32367 13929
rect 32309 13920 32321 13923
rect 32180 13892 32321 13920
rect 32180 13880 32186 13892
rect 32309 13889 32321 13892
rect 32355 13889 32367 13923
rect 32309 13883 32367 13889
rect 32398 13880 32404 13932
rect 32456 13920 32462 13932
rect 32493 13923 32551 13929
rect 32493 13920 32505 13923
rect 32456 13892 32505 13920
rect 32456 13880 32462 13892
rect 32493 13889 32505 13892
rect 32539 13889 32551 13923
rect 32493 13883 32551 13889
rect 33965 13923 34023 13929
rect 33965 13889 33977 13923
rect 34011 13889 34023 13923
rect 33965 13883 34023 13889
rect 33980 13852 34008 13883
rect 34422 13880 34428 13932
rect 34480 13920 34486 13932
rect 37090 13920 37096 13932
rect 34480 13892 37096 13920
rect 34480 13880 34486 13892
rect 37090 13880 37096 13892
rect 37148 13880 37154 13932
rect 38749 13923 38807 13929
rect 38749 13889 38761 13923
rect 38795 13920 38807 13923
rect 50706 13920 50712 13932
rect 38795 13892 50712 13920
rect 38795 13889 38807 13892
rect 38749 13883 38807 13889
rect 50706 13880 50712 13892
rect 50764 13880 50770 13932
rect 57057 13923 57115 13929
rect 57057 13889 57069 13923
rect 57103 13920 57115 13923
rect 58250 13920 58256 13932
rect 57103 13892 58256 13920
rect 57103 13889 57115 13892
rect 57057 13883 57115 13889
rect 58250 13880 58256 13892
rect 58308 13880 58314 13932
rect 34238 13852 34244 13864
rect 30852 13824 31248 13852
rect 31312 13824 34244 13852
rect 30190 13784 30196 13796
rect 29656 13756 30196 13784
rect 28092 13728 28120 13756
rect 30190 13744 30196 13756
rect 30248 13744 30254 13796
rect 30561 13787 30619 13793
rect 30561 13753 30573 13787
rect 30607 13784 30619 13787
rect 31110 13784 31116 13796
rect 30607 13756 31116 13784
rect 30607 13753 30619 13756
rect 30561 13747 30619 13753
rect 31110 13744 31116 13756
rect 31168 13744 31174 13796
rect 28074 13716 28080 13728
rect 27172 13688 28080 13716
rect 28074 13676 28080 13688
rect 28132 13676 28138 13728
rect 28994 13716 29000 13728
rect 28955 13688 29000 13716
rect 28994 13676 29000 13688
rect 29052 13676 29058 13728
rect 31220 13716 31248 13824
rect 34238 13812 34244 13824
rect 34296 13812 34302 13864
rect 57330 13852 57336 13864
rect 57291 13824 57336 13852
rect 57330 13812 57336 13824
rect 57388 13812 57394 13864
rect 31662 13744 31668 13796
rect 31720 13784 31726 13796
rect 44818 13784 44824 13796
rect 31720 13756 32536 13784
rect 31720 13744 31726 13756
rect 31846 13716 31852 13728
rect 31220 13688 31852 13716
rect 31846 13676 31852 13688
rect 31904 13676 31910 13728
rect 32508 13716 32536 13756
rect 32692 13756 44824 13784
rect 32692 13716 32720 13756
rect 44818 13744 44824 13756
rect 44876 13744 44882 13796
rect 34146 13716 34152 13728
rect 32508 13688 32720 13716
rect 34107 13688 34152 13716
rect 34146 13676 34152 13688
rect 34204 13676 34210 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 17218 13472 17224 13524
rect 17276 13512 17282 13524
rect 20165 13515 20223 13521
rect 20165 13512 20177 13515
rect 17276 13484 20177 13512
rect 17276 13472 17282 13484
rect 20165 13481 20177 13484
rect 20211 13512 20223 13515
rect 22094 13512 22100 13524
rect 20211 13484 22100 13512
rect 20211 13481 20223 13484
rect 20165 13475 20223 13481
rect 22094 13472 22100 13484
rect 22152 13472 22158 13524
rect 22278 13512 22284 13524
rect 22239 13484 22284 13512
rect 22278 13472 22284 13484
rect 22336 13472 22342 13524
rect 23842 13512 23848 13524
rect 23803 13484 23848 13512
rect 23842 13472 23848 13484
rect 23900 13472 23906 13524
rect 34238 13512 34244 13524
rect 25240 13484 34100 13512
rect 34199 13484 34244 13512
rect 18874 13404 18880 13456
rect 18932 13444 18938 13456
rect 25240 13444 25268 13484
rect 18932 13416 25268 13444
rect 18932 13404 18938 13416
rect 31110 13404 31116 13456
rect 31168 13444 31174 13456
rect 32214 13444 32220 13456
rect 31168 13416 32220 13444
rect 31168 13404 31174 13416
rect 32214 13404 32220 13416
rect 32272 13404 32278 13456
rect 34072 13444 34100 13484
rect 34238 13472 34244 13484
rect 34296 13472 34302 13524
rect 58250 13512 58256 13524
rect 58211 13484 58256 13512
rect 58250 13472 58256 13484
rect 58308 13472 58314 13524
rect 39298 13444 39304 13456
rect 34072 13416 39304 13444
rect 39298 13404 39304 13416
rect 39356 13404 39362 13456
rect 14461 13379 14519 13385
rect 14461 13345 14473 13379
rect 14507 13376 14519 13379
rect 14642 13376 14648 13388
rect 14507 13348 14648 13376
rect 14507 13345 14519 13348
rect 14461 13339 14519 13345
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 14737 13379 14795 13385
rect 14737 13345 14749 13379
rect 14783 13376 14795 13379
rect 17681 13379 17739 13385
rect 17681 13376 17693 13379
rect 14783 13348 17693 13376
rect 14783 13345 14795 13348
rect 14737 13339 14795 13345
rect 17681 13345 17693 13348
rect 17727 13345 17739 13379
rect 17681 13339 17739 13345
rect 19334 13336 19340 13388
rect 19392 13376 19398 13388
rect 19797 13379 19855 13385
rect 19797 13376 19809 13379
rect 19392 13348 19809 13376
rect 19392 13336 19398 13348
rect 19797 13345 19809 13348
rect 19843 13376 19855 13379
rect 21818 13376 21824 13388
rect 19843 13348 21824 13376
rect 19843 13345 19855 13348
rect 19797 13339 19855 13345
rect 21818 13336 21824 13348
rect 21876 13336 21882 13388
rect 24762 13376 24768 13388
rect 23860 13348 24768 13376
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 1854 13308 1860 13320
rect 1815 13280 1860 13308
rect 1854 13268 1860 13280
rect 1912 13268 1918 13320
rect 16574 13308 16580 13320
rect 16535 13280 16580 13308
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 18782 13268 18788 13320
rect 18840 13308 18846 13320
rect 19889 13311 19947 13317
rect 19889 13308 19901 13311
rect 18840 13280 19901 13308
rect 18840 13268 18846 13280
rect 19889 13277 19901 13280
rect 19935 13277 19947 13311
rect 21082 13308 21088 13320
rect 21043 13280 21088 13308
rect 19889 13271 19947 13277
rect 21082 13268 21088 13280
rect 21140 13268 21146 13320
rect 23860 13317 23888 13348
rect 24762 13336 24768 13348
rect 24820 13336 24826 13388
rect 25682 13376 25688 13388
rect 25643 13348 25688 13376
rect 25682 13336 25688 13348
rect 25740 13336 25746 13388
rect 27246 13336 27252 13388
rect 27304 13376 27310 13388
rect 27341 13379 27399 13385
rect 27341 13376 27353 13379
rect 27304 13348 27353 13376
rect 27304 13336 27310 13348
rect 27341 13345 27353 13348
rect 27387 13345 27399 13379
rect 32861 13379 32919 13385
rect 32861 13376 32873 13379
rect 27341 13339 27399 13345
rect 31726 13348 32873 13376
rect 23845 13311 23903 13317
rect 23845 13277 23857 13311
rect 23891 13277 23903 13311
rect 23845 13271 23903 13277
rect 24029 13311 24087 13317
rect 24029 13277 24041 13311
rect 24075 13277 24087 13311
rect 24029 13271 24087 13277
rect 24581 13311 24639 13317
rect 24581 13277 24593 13311
rect 24627 13308 24639 13311
rect 25130 13308 25136 13320
rect 24627 13280 25136 13308
rect 24627 13277 24639 13280
rect 24581 13271 24639 13277
rect 17218 13200 17224 13252
rect 17276 13240 17282 13252
rect 17862 13240 17868 13252
rect 17276 13212 17868 13240
rect 17276 13200 17282 13212
rect 17862 13200 17868 13212
rect 17920 13200 17926 13252
rect 19521 13243 19579 13249
rect 19521 13209 19533 13243
rect 19567 13209 19579 13243
rect 19978 13240 19984 13252
rect 19939 13212 19984 13240
rect 19521 13203 19579 13209
rect 16025 13175 16083 13181
rect 16025 13141 16037 13175
rect 16071 13172 16083 13175
rect 18966 13172 18972 13184
rect 16071 13144 18972 13172
rect 16071 13141 16083 13144
rect 16025 13135 16083 13141
rect 18966 13132 18972 13144
rect 19024 13132 19030 13184
rect 19536 13172 19564 13203
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 20622 13240 20628 13252
rect 20088 13212 20628 13240
rect 19886 13172 19892 13184
rect 19536 13144 19892 13172
rect 19886 13132 19892 13144
rect 19944 13172 19950 13184
rect 20088 13172 20116 13212
rect 20622 13200 20628 13212
rect 20680 13200 20686 13252
rect 24044 13240 24072 13271
rect 25130 13268 25136 13280
rect 25188 13268 25194 13320
rect 27608 13311 27666 13317
rect 27608 13277 27620 13311
rect 27654 13308 27666 13311
rect 28994 13308 29000 13320
rect 27654 13280 29000 13308
rect 27654 13277 27666 13280
rect 27608 13271 27666 13277
rect 28994 13268 29000 13280
rect 29052 13268 29058 13320
rect 29733 13311 29791 13317
rect 29733 13277 29745 13311
rect 29779 13308 29791 13311
rect 30282 13308 30288 13320
rect 29779 13280 30288 13308
rect 29779 13277 29791 13280
rect 29733 13271 29791 13277
rect 30282 13268 30288 13280
rect 30340 13308 30346 13320
rect 31726 13308 31754 13348
rect 32861 13345 32873 13348
rect 32907 13345 32919 13379
rect 56870 13376 56876 13388
rect 56831 13348 56876 13376
rect 32861 13339 32919 13345
rect 56870 13336 56876 13348
rect 56928 13336 56934 13388
rect 31846 13308 31852 13320
rect 30340 13280 31754 13308
rect 31807 13280 31852 13308
rect 30340 13268 30346 13280
rect 31846 13268 31852 13280
rect 31904 13268 31910 13320
rect 31938 13268 31944 13320
rect 31996 13308 32002 13320
rect 32125 13311 32183 13317
rect 31996 13280 32041 13308
rect 31996 13268 32002 13280
rect 32125 13277 32137 13311
rect 32171 13277 32183 13311
rect 32125 13271 32183 13277
rect 25038 13240 25044 13252
rect 24044 13212 25044 13240
rect 25038 13200 25044 13212
rect 25096 13200 25102 13252
rect 30000 13243 30058 13249
rect 30000 13209 30012 13243
rect 30046 13240 30058 13243
rect 30834 13240 30840 13252
rect 30046 13212 30840 13240
rect 30046 13209 30058 13212
rect 30000 13203 30058 13209
rect 30834 13200 30840 13212
rect 30892 13200 30898 13252
rect 31754 13200 31760 13252
rect 31812 13240 31818 13252
rect 32140 13240 32168 13271
rect 32214 13268 32220 13320
rect 32272 13308 32278 13320
rect 32272 13280 32317 13308
rect 32272 13268 32278 13280
rect 31812 13212 32168 13240
rect 33128 13243 33186 13249
rect 31812 13200 31818 13212
rect 33128 13209 33140 13243
rect 33174 13240 33186 13243
rect 33686 13240 33692 13252
rect 33174 13212 33692 13240
rect 33174 13209 33186 13212
rect 33128 13203 33186 13209
rect 33686 13200 33692 13212
rect 33744 13200 33750 13252
rect 46198 13240 46204 13252
rect 34164 13212 46204 13240
rect 19944 13144 20116 13172
rect 19944 13132 19950 13144
rect 21450 13132 21456 13184
rect 21508 13172 21514 13184
rect 28718 13172 28724 13184
rect 21508 13144 28724 13172
rect 21508 13132 21514 13144
rect 28718 13132 28724 13144
rect 28776 13132 28782 13184
rect 31110 13172 31116 13184
rect 31071 13144 31116 13172
rect 31110 13132 31116 13144
rect 31168 13132 31174 13184
rect 31665 13175 31723 13181
rect 31665 13141 31677 13175
rect 31711 13172 31723 13175
rect 34164 13172 34192 13212
rect 46198 13200 46204 13212
rect 46256 13200 46262 13252
rect 56778 13200 56784 13252
rect 56836 13240 56842 13252
rect 57118 13243 57176 13249
rect 57118 13240 57130 13243
rect 56836 13212 57130 13240
rect 56836 13200 56842 13212
rect 57118 13209 57130 13212
rect 57164 13209 57176 13243
rect 57118 13203 57176 13209
rect 31711 13144 34192 13172
rect 31711 13141 31723 13144
rect 31665 13135 31723 13141
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 1578 12928 1584 12980
rect 1636 12968 1642 12980
rect 1636 12940 16988 12968
rect 1636 12928 1642 12940
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12832 1639 12835
rect 12342 12832 12348 12844
rect 1627 12804 12348 12832
rect 1627 12801 1639 12804
rect 1581 12795 1639 12801
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 14642 12832 14648 12844
rect 14603 12804 14648 12832
rect 14642 12792 14648 12804
rect 14700 12792 14706 12844
rect 1762 12764 1768 12776
rect 1723 12736 1768 12764
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 14921 12767 14979 12773
rect 14921 12733 14933 12767
rect 14967 12764 14979 12767
rect 15102 12764 15108 12776
rect 14967 12736 15108 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 16960 12696 16988 12940
rect 18138 12928 18144 12980
rect 18196 12968 18202 12980
rect 18693 12971 18751 12977
rect 18693 12968 18705 12971
rect 18196 12940 18705 12968
rect 18196 12928 18202 12940
rect 18693 12937 18705 12940
rect 18739 12937 18751 12971
rect 18693 12931 18751 12937
rect 18966 12928 18972 12980
rect 19024 12968 19030 12980
rect 22189 12971 22247 12977
rect 19024 12940 22048 12968
rect 19024 12928 19030 12940
rect 20898 12900 20904 12912
rect 20859 12872 20904 12900
rect 20898 12860 20904 12872
rect 20956 12860 20962 12912
rect 17494 12832 17500 12844
rect 17455 12804 17500 12832
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 20714 12832 20720 12844
rect 20675 12804 20720 12832
rect 20714 12792 20720 12804
rect 20772 12792 20778 12844
rect 20993 12767 21051 12773
rect 20993 12733 21005 12767
rect 21039 12764 21051 12767
rect 21634 12764 21640 12776
rect 21039 12736 21640 12764
rect 21039 12733 21051 12736
rect 20993 12727 21051 12733
rect 21634 12724 21640 12736
rect 21692 12724 21698 12776
rect 22020 12764 22048 12940
rect 22189 12937 22201 12971
rect 22235 12968 22247 12971
rect 22278 12968 22284 12980
rect 22235 12940 22284 12968
rect 22235 12937 22247 12940
rect 22189 12931 22247 12937
rect 22278 12928 22284 12940
rect 22336 12928 22342 12980
rect 25866 12968 25872 12980
rect 23400 12940 25872 12968
rect 22094 12860 22100 12912
rect 22152 12900 22158 12912
rect 22373 12903 22431 12909
rect 22373 12900 22385 12903
rect 22152 12872 22385 12900
rect 22152 12860 22158 12872
rect 22373 12869 22385 12872
rect 22419 12869 22431 12903
rect 23400 12900 23428 12940
rect 25866 12928 25872 12940
rect 25924 12928 25930 12980
rect 26234 12928 26240 12980
rect 26292 12968 26298 12980
rect 27249 12971 27307 12977
rect 27249 12968 27261 12971
rect 26292 12940 27261 12968
rect 26292 12928 26298 12940
rect 27249 12937 27261 12940
rect 27295 12937 27307 12971
rect 30834 12968 30840 12980
rect 30795 12940 30840 12968
rect 27249 12931 27307 12937
rect 30834 12928 30840 12940
rect 30892 12928 30898 12980
rect 31202 12968 31208 12980
rect 31163 12940 31208 12968
rect 31202 12928 31208 12940
rect 31260 12928 31266 12980
rect 33686 12968 33692 12980
rect 33647 12940 33692 12968
rect 33686 12928 33692 12940
rect 33744 12928 33750 12980
rect 46198 12928 46204 12980
rect 46256 12968 46262 12980
rect 58253 12971 58311 12977
rect 58253 12968 58265 12971
rect 46256 12940 56916 12968
rect 46256 12928 46262 12940
rect 22373 12863 22431 12869
rect 23308 12872 23428 12900
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12832 22339 12835
rect 22646 12832 22652 12844
rect 22327 12804 22652 12832
rect 22327 12801 22339 12804
rect 22281 12795 22339 12801
rect 22646 12792 22652 12804
rect 22704 12832 22710 12844
rect 23308 12832 23336 12872
rect 23934 12860 23940 12912
rect 23992 12900 23998 12912
rect 26329 12903 26387 12909
rect 23992 12872 26280 12900
rect 23992 12860 23998 12872
rect 22704 12804 23336 12832
rect 23385 12835 23443 12841
rect 22704 12792 22710 12804
rect 23385 12801 23397 12835
rect 23431 12832 23443 12835
rect 23750 12832 23756 12844
rect 23431 12804 23756 12832
rect 23431 12801 23443 12804
rect 23385 12795 23443 12801
rect 23750 12792 23756 12804
rect 23808 12792 23814 12844
rect 24118 12792 24124 12844
rect 24176 12832 24182 12844
rect 26142 12832 26148 12844
rect 24176 12804 24992 12832
rect 26103 12804 26148 12832
rect 24176 12792 24182 12804
rect 22554 12764 22560 12776
rect 22020 12736 22416 12764
rect 22515 12736 22560 12764
rect 21542 12696 21548 12708
rect 16960 12668 21548 12696
rect 21542 12656 21548 12668
rect 21600 12656 21606 12708
rect 22005 12699 22063 12705
rect 22005 12665 22017 12699
rect 22051 12665 22063 12699
rect 22388 12696 22416 12736
rect 22554 12724 22560 12736
rect 22612 12764 22618 12776
rect 23198 12764 23204 12776
rect 22612 12736 23204 12764
rect 22612 12724 22618 12736
rect 23198 12724 23204 12736
rect 23256 12724 23262 12776
rect 24854 12764 24860 12776
rect 24815 12736 24860 12764
rect 24854 12724 24860 12736
rect 24912 12724 24918 12776
rect 24964 12764 24992 12804
rect 26142 12792 26148 12804
rect 26200 12792 26206 12844
rect 26252 12832 26280 12872
rect 26329 12869 26341 12903
rect 26375 12900 26387 12903
rect 29086 12900 29092 12912
rect 26375 12872 29092 12900
rect 26375 12869 26387 12872
rect 26329 12863 26387 12869
rect 29086 12860 29092 12872
rect 29144 12860 29150 12912
rect 33410 12900 33416 12912
rect 29196 12872 33416 12900
rect 26421 12835 26479 12841
rect 26421 12832 26433 12835
rect 26252 12804 26433 12832
rect 26421 12801 26433 12804
rect 26467 12801 26479 12835
rect 26421 12795 26479 12801
rect 26510 12792 26516 12844
rect 26568 12832 26574 12844
rect 27062 12832 27068 12844
rect 26568 12804 27068 12832
rect 26568 12792 26574 12804
rect 27062 12792 27068 12804
rect 27120 12832 27126 12844
rect 27157 12835 27215 12841
rect 27157 12832 27169 12835
rect 27120 12804 27169 12832
rect 27120 12792 27126 12804
rect 27157 12801 27169 12804
rect 27203 12801 27215 12835
rect 27338 12832 27344 12844
rect 27299 12804 27344 12832
rect 27157 12795 27215 12801
rect 27338 12792 27344 12804
rect 27396 12792 27402 12844
rect 28074 12832 28080 12844
rect 28035 12804 28080 12832
rect 28074 12792 28080 12804
rect 28132 12792 28138 12844
rect 29196 12764 29224 12872
rect 33410 12860 33416 12872
rect 33468 12860 33474 12912
rect 36538 12900 36544 12912
rect 33980 12872 36544 12900
rect 31202 12792 31208 12844
rect 31260 12832 31266 12844
rect 33980 12841 34008 12872
rect 36538 12860 36544 12872
rect 36596 12900 36602 12912
rect 37182 12900 37188 12912
rect 36596 12872 37188 12900
rect 36596 12860 36602 12872
rect 37182 12860 37188 12872
rect 37240 12860 37246 12912
rect 46842 12860 46848 12912
rect 46900 12900 46906 12912
rect 49421 12903 49479 12909
rect 49421 12900 49433 12903
rect 46900 12872 49433 12900
rect 46900 12860 46906 12872
rect 49421 12869 49433 12872
rect 49467 12869 49479 12903
rect 49421 12863 49479 12869
rect 33965 12835 34023 12841
rect 31260 12804 33916 12832
rect 31260 12792 31266 12804
rect 24964 12736 29224 12764
rect 30190 12724 30196 12776
rect 30248 12764 30254 12776
rect 31110 12764 31116 12776
rect 30248 12736 31116 12764
rect 30248 12724 30254 12736
rect 31110 12724 31116 12736
rect 31168 12764 31174 12776
rect 31297 12767 31355 12773
rect 31297 12764 31309 12767
rect 31168 12736 31309 12764
rect 31168 12724 31174 12736
rect 31297 12733 31309 12736
rect 31343 12733 31355 12767
rect 31297 12727 31355 12733
rect 31389 12767 31447 12773
rect 31389 12733 31401 12767
rect 31435 12764 31447 12767
rect 32582 12764 32588 12776
rect 31435 12736 32588 12764
rect 31435 12733 31447 12736
rect 31389 12727 31447 12733
rect 22462 12696 22468 12708
rect 22388 12668 22468 12696
rect 22005 12659 22063 12665
rect 16022 12628 16028 12640
rect 15983 12600 16028 12628
rect 16022 12588 16028 12600
rect 16080 12588 16086 12640
rect 20438 12628 20444 12640
rect 20399 12600 20444 12628
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 22020 12628 22048 12659
rect 22462 12656 22468 12668
rect 22520 12656 22526 12708
rect 26145 12699 26203 12705
rect 26145 12665 26157 12699
rect 26191 12696 26203 12699
rect 26326 12696 26332 12708
rect 26191 12668 26332 12696
rect 26191 12665 26203 12668
rect 26145 12659 26203 12665
rect 26326 12656 26332 12668
rect 26384 12656 26390 12708
rect 28994 12656 29000 12708
rect 29052 12696 29058 12708
rect 31404 12696 31432 12727
rect 32582 12724 32588 12736
rect 32640 12724 32646 12776
rect 33888 12764 33916 12804
rect 33965 12801 33977 12835
rect 34011 12801 34023 12835
rect 33965 12795 34023 12801
rect 34057 12835 34115 12841
rect 34057 12801 34069 12835
rect 34103 12801 34115 12835
rect 34057 12795 34115 12801
rect 34072 12764 34100 12795
rect 34146 12792 34152 12844
rect 34204 12832 34210 12844
rect 34333 12835 34391 12841
rect 34204 12804 34249 12832
rect 34204 12792 34210 12804
rect 34333 12801 34345 12835
rect 34379 12801 34391 12835
rect 34333 12795 34391 12801
rect 33888 12736 34100 12764
rect 29052 12668 31432 12696
rect 29052 12656 29058 12668
rect 31478 12656 31484 12708
rect 31536 12696 31542 12708
rect 34348 12696 34376 12795
rect 56594 12792 56600 12844
rect 56652 12832 56658 12844
rect 56781 12835 56839 12841
rect 56781 12832 56793 12835
rect 56652 12804 56793 12832
rect 56652 12792 56658 12804
rect 56781 12801 56793 12804
rect 56827 12801 56839 12835
rect 56888 12832 56916 12940
rect 56980 12940 58265 12968
rect 56980 12909 57008 12940
rect 58253 12937 58265 12940
rect 58299 12937 58311 12971
rect 58253 12931 58311 12937
rect 56965 12903 57023 12909
rect 56965 12869 56977 12903
rect 57011 12869 57023 12903
rect 56965 12863 57023 12869
rect 57057 12835 57115 12841
rect 57057 12832 57069 12835
rect 56888 12804 57069 12832
rect 56781 12795 56839 12801
rect 57057 12801 57069 12804
rect 57103 12801 57115 12835
rect 57057 12795 57115 12801
rect 58069 12835 58127 12841
rect 58069 12801 58081 12835
rect 58115 12801 58127 12835
rect 58250 12832 58256 12844
rect 58211 12804 58256 12832
rect 58069 12795 58127 12801
rect 56410 12724 56416 12776
rect 56468 12764 56474 12776
rect 57882 12764 57888 12776
rect 56468 12736 57888 12764
rect 56468 12724 56474 12736
rect 57882 12724 57888 12736
rect 57940 12764 57946 12776
rect 58084 12764 58112 12795
rect 58250 12792 58256 12804
rect 58308 12792 58314 12844
rect 57940 12736 58112 12764
rect 57940 12724 57946 12736
rect 56778 12696 56784 12708
rect 31536 12668 34376 12696
rect 56739 12668 56784 12696
rect 31536 12656 31542 12668
rect 56778 12656 56784 12668
rect 56836 12656 56842 12708
rect 23106 12628 23112 12640
rect 22020 12600 23112 12628
rect 23106 12588 23112 12600
rect 23164 12628 23170 12640
rect 29273 12631 29331 12637
rect 29273 12628 29285 12631
rect 23164 12600 29285 12628
rect 23164 12588 23170 12600
rect 29273 12597 29285 12600
rect 29319 12597 29331 12631
rect 29273 12591 29331 12597
rect 30650 12588 30656 12640
rect 30708 12628 30714 12640
rect 31662 12628 31668 12640
rect 30708 12600 31668 12628
rect 30708 12588 30714 12600
rect 31662 12588 31668 12600
rect 31720 12588 31726 12640
rect 32766 12588 32772 12640
rect 32824 12628 32830 12640
rect 37458 12628 37464 12640
rect 32824 12600 37464 12628
rect 32824 12588 32830 12600
rect 37458 12588 37464 12600
rect 37516 12588 37522 12640
rect 40770 12588 40776 12640
rect 40828 12628 40834 12640
rect 43254 12628 43260 12640
rect 40828 12600 43260 12628
rect 40828 12588 40834 12600
rect 43254 12588 43260 12600
rect 43312 12588 43318 12640
rect 50893 12631 50951 12637
rect 50893 12597 50905 12631
rect 50939 12628 50951 12631
rect 56870 12628 56876 12640
rect 50939 12600 56876 12628
rect 50939 12597 50951 12600
rect 50893 12591 50951 12597
rect 56870 12588 56876 12600
rect 56928 12588 56934 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 12400 12396 13093 12424
rect 12400 12384 12406 12396
rect 13081 12393 13093 12396
rect 13127 12393 13139 12427
rect 13081 12387 13139 12393
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 16666 12424 16672 12436
rect 13872 12396 16672 12424
rect 13872 12384 13878 12396
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 17126 12384 17132 12436
rect 17184 12424 17190 12436
rect 17773 12427 17831 12433
rect 17773 12424 17785 12427
rect 17184 12396 17785 12424
rect 17184 12384 17190 12396
rect 17773 12393 17785 12396
rect 17819 12393 17831 12427
rect 17773 12387 17831 12393
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19981 12427 20039 12433
rect 19981 12424 19993 12427
rect 19484 12396 19993 12424
rect 19484 12384 19490 12396
rect 19981 12393 19993 12396
rect 20027 12393 20039 12427
rect 19981 12387 20039 12393
rect 21818 12384 21824 12436
rect 21876 12424 21882 12436
rect 27249 12427 27307 12433
rect 27249 12424 27261 12427
rect 21876 12396 27261 12424
rect 21876 12384 21882 12396
rect 27249 12393 27261 12396
rect 27295 12393 27307 12427
rect 27249 12387 27307 12393
rect 31021 12427 31079 12433
rect 31021 12393 31033 12427
rect 31067 12424 31079 12427
rect 31938 12424 31944 12436
rect 31067 12396 31944 12424
rect 31067 12393 31079 12396
rect 31021 12387 31079 12393
rect 31938 12384 31944 12396
rect 31996 12384 32002 12436
rect 19886 12356 19892 12368
rect 13372 12328 19892 12356
rect 13372 12297 13400 12328
rect 19886 12316 19892 12328
rect 19944 12316 19950 12368
rect 20990 12316 20996 12368
rect 21048 12356 21054 12368
rect 30190 12356 30196 12368
rect 21048 12328 30196 12356
rect 21048 12316 21054 12328
rect 30190 12316 30196 12328
rect 30248 12316 30254 12368
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12257 13415 12291
rect 13357 12251 13415 12257
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12288 13507 12291
rect 13814 12288 13820 12300
rect 13495 12260 13820 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 13814 12248 13820 12260
rect 13872 12248 13878 12300
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12288 15899 12291
rect 17034 12288 17040 12300
rect 15887 12260 17040 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 17126 12248 17132 12300
rect 17184 12288 17190 12300
rect 20349 12291 20407 12297
rect 20349 12288 20361 12291
rect 17184 12260 20361 12288
rect 17184 12248 17190 12260
rect 20349 12257 20361 12260
rect 20395 12257 20407 12291
rect 20349 12251 20407 12257
rect 25225 12291 25283 12297
rect 25225 12257 25237 12291
rect 25271 12288 25283 12291
rect 27154 12288 27160 12300
rect 25271 12260 27160 12288
rect 25271 12257 25283 12260
rect 25225 12251 25283 12257
rect 27154 12248 27160 12260
rect 27212 12288 27218 12300
rect 30282 12288 30288 12300
rect 27212 12260 30288 12288
rect 27212 12248 27218 12260
rect 30282 12248 30288 12260
rect 30340 12248 30346 12300
rect 1581 12223 1639 12229
rect 1581 12189 1593 12223
rect 1627 12220 1639 12223
rect 12986 12220 12992 12232
rect 1627 12192 12992 12220
rect 1627 12189 1639 12192
rect 1581 12183 1639 12189
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 13262 12220 13268 12232
rect 13223 12192 13268 12220
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 13538 12180 13544 12232
rect 13596 12220 13602 12232
rect 15749 12223 15807 12229
rect 13596 12192 13641 12220
rect 13596 12180 13602 12192
rect 15749 12189 15761 12223
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 1854 12152 1860 12164
rect 1815 12124 1860 12152
rect 1854 12112 1860 12124
rect 1912 12112 1918 12164
rect 15764 12152 15792 12183
rect 16114 12180 16120 12232
rect 16172 12220 16178 12232
rect 16577 12223 16635 12229
rect 16577 12220 16589 12223
rect 16172 12192 16589 12220
rect 16172 12180 16178 12192
rect 16577 12189 16589 12192
rect 16623 12189 16635 12223
rect 16577 12183 16635 12189
rect 16666 12180 16672 12232
rect 16724 12220 16730 12232
rect 18414 12220 18420 12232
rect 16724 12192 18420 12220
rect 16724 12180 16730 12192
rect 18414 12180 18420 12192
rect 18472 12220 18478 12232
rect 20533 12223 20591 12229
rect 20533 12220 20545 12223
rect 18472 12192 20545 12220
rect 18472 12180 18478 12192
rect 20533 12189 20545 12192
rect 20579 12189 20591 12223
rect 20533 12183 20591 12189
rect 21729 12223 21787 12229
rect 21729 12189 21741 12223
rect 21775 12220 21787 12223
rect 25498 12220 25504 12232
rect 21775 12192 25504 12220
rect 21775 12189 21787 12192
rect 21729 12183 21787 12189
rect 25498 12180 25504 12192
rect 25556 12180 25562 12232
rect 26050 12220 26056 12232
rect 26011 12192 26056 12220
rect 26050 12180 26056 12192
rect 26108 12180 26114 12232
rect 30098 12220 30104 12232
rect 30059 12192 30104 12220
rect 30098 12180 30104 12192
rect 30156 12180 30162 12232
rect 30929 12223 30987 12229
rect 30929 12189 30941 12223
rect 30975 12189 30987 12223
rect 30929 12183 30987 12189
rect 17954 12152 17960 12164
rect 15764 12124 17960 12152
rect 17954 12112 17960 12124
rect 18012 12112 18018 12164
rect 20438 12152 20444 12164
rect 20399 12124 20444 12152
rect 20438 12112 20444 12124
rect 20496 12112 20502 12164
rect 20806 12112 20812 12164
rect 20864 12152 20870 12164
rect 20990 12152 20996 12164
rect 20864 12124 20996 12152
rect 20864 12112 20870 12124
rect 20990 12112 20996 12124
rect 21048 12112 21054 12164
rect 22186 12112 22192 12164
rect 22244 12152 22250 12164
rect 23198 12152 23204 12164
rect 22244 12124 23204 12152
rect 22244 12112 22250 12124
rect 23198 12112 23204 12124
rect 23256 12112 23262 12164
rect 24949 12155 25007 12161
rect 24949 12121 24961 12155
rect 24995 12152 25007 12155
rect 28166 12152 28172 12164
rect 24995 12124 28172 12152
rect 24995 12121 25007 12124
rect 24949 12115 25007 12121
rect 28166 12112 28172 12124
rect 28224 12112 28230 12164
rect 29086 12112 29092 12164
rect 29144 12152 29150 12164
rect 30944 12152 30972 12183
rect 33870 12180 33876 12232
rect 33928 12220 33934 12232
rect 40034 12220 40040 12232
rect 33928 12192 40040 12220
rect 33928 12180 33934 12192
rect 40034 12180 40040 12192
rect 40092 12180 40098 12232
rect 56965 12223 57023 12229
rect 56965 12189 56977 12223
rect 57011 12220 57023 12223
rect 57974 12220 57980 12232
rect 57011 12192 57836 12220
rect 57935 12192 57980 12220
rect 57011 12189 57023 12192
rect 56965 12183 57023 12189
rect 38286 12152 38292 12164
rect 29144 12124 30972 12152
rect 31726 12124 38292 12152
rect 29144 12112 29150 12124
rect 16114 12084 16120 12096
rect 16075 12056 16120 12084
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16482 12044 16488 12096
rect 16540 12084 16546 12096
rect 22278 12084 22284 12096
rect 16540 12056 22284 12084
rect 16540 12044 16546 12056
rect 22278 12044 22284 12056
rect 22336 12044 22342 12096
rect 22370 12044 22376 12096
rect 22428 12084 22434 12096
rect 23014 12084 23020 12096
rect 22428 12056 23020 12084
rect 22428 12044 22434 12056
rect 23014 12044 23020 12056
rect 23072 12084 23078 12096
rect 23109 12087 23167 12093
rect 23109 12084 23121 12087
rect 23072 12056 23121 12084
rect 23072 12044 23078 12056
rect 23109 12053 23121 12056
rect 23155 12053 23167 12087
rect 23109 12047 23167 12053
rect 23934 12044 23940 12096
rect 23992 12084 23998 12096
rect 24581 12087 24639 12093
rect 24581 12084 24593 12087
rect 23992 12056 24593 12084
rect 23992 12044 23998 12056
rect 24581 12053 24593 12056
rect 24627 12053 24639 12087
rect 25038 12084 25044 12096
rect 24999 12056 25044 12084
rect 24581 12047 24639 12053
rect 25038 12044 25044 12056
rect 25096 12044 25102 12096
rect 27890 12044 27896 12096
rect 27948 12084 27954 12096
rect 28442 12084 28448 12096
rect 27948 12056 28448 12084
rect 27948 12044 27954 12056
rect 28442 12044 28448 12056
rect 28500 12044 28506 12096
rect 29730 12084 29736 12096
rect 29691 12056 29736 12084
rect 29730 12044 29736 12056
rect 29788 12044 29794 12096
rect 30190 12084 30196 12096
rect 30151 12056 30196 12084
rect 30190 12044 30196 12056
rect 30248 12044 30254 12096
rect 30282 12044 30288 12096
rect 30340 12084 30346 12096
rect 31726 12084 31754 12124
rect 38286 12112 38292 12124
rect 38344 12112 38350 12164
rect 57238 12152 57244 12164
rect 57199 12124 57244 12152
rect 57238 12112 57244 12124
rect 57296 12112 57302 12164
rect 57808 12152 57836 12192
rect 57974 12180 57980 12192
rect 58032 12180 58038 12232
rect 58250 12152 58256 12164
rect 57808 12124 58256 12152
rect 58250 12112 58256 12124
rect 58308 12112 58314 12164
rect 30340 12056 31754 12084
rect 30340 12044 30346 12056
rect 32674 12044 32680 12096
rect 32732 12084 32738 12096
rect 35434 12084 35440 12096
rect 32732 12056 35440 12084
rect 32732 12044 32738 12056
rect 35434 12044 35440 12056
rect 35492 12044 35498 12096
rect 37182 12044 37188 12096
rect 37240 12084 37246 12096
rect 58069 12087 58127 12093
rect 58069 12084 58081 12087
rect 37240 12056 58081 12084
rect 37240 12044 37246 12056
rect 58069 12053 58081 12056
rect 58115 12053 58127 12087
rect 58069 12047 58127 12053
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 12986 11880 12992 11892
rect 12947 11852 12992 11880
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 15930 11880 15936 11892
rect 15891 11852 15936 11880
rect 15930 11840 15936 11852
rect 15988 11840 15994 11892
rect 16022 11840 16028 11892
rect 16080 11880 16086 11892
rect 16482 11880 16488 11892
rect 16080 11852 16488 11880
rect 16080 11840 16086 11852
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 17034 11880 17040 11892
rect 16995 11852 17040 11880
rect 17034 11840 17040 11852
rect 17092 11840 17098 11892
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 17589 11883 17647 11889
rect 17589 11880 17601 11883
rect 17552 11852 17601 11880
rect 17552 11840 17558 11852
rect 17589 11849 17601 11852
rect 17635 11849 17647 11883
rect 17589 11843 17647 11849
rect 17770 11840 17776 11892
rect 17828 11880 17834 11892
rect 19058 11880 19064 11892
rect 17828 11852 19064 11880
rect 17828 11840 17834 11852
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 19426 11840 19432 11892
rect 19484 11880 19490 11892
rect 19484 11852 21680 11880
rect 19484 11840 19490 11852
rect 13262 11812 13268 11824
rect 13175 11784 13268 11812
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11744 1639 11747
rect 11054 11744 11060 11756
rect 1627 11716 11060 11744
rect 1627 11713 1639 11716
rect 1581 11707 1639 11713
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 13188 11753 13216 11784
rect 13262 11772 13268 11784
rect 13320 11812 13326 11824
rect 17402 11812 17408 11824
rect 13320 11784 17408 11812
rect 13320 11772 13326 11784
rect 17402 11772 17408 11784
rect 17460 11772 17466 11824
rect 19334 11812 19340 11824
rect 17880 11784 19340 11812
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11744 13415 11747
rect 13814 11744 13820 11756
rect 13403 11716 13820 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 15378 11704 15384 11756
rect 15436 11744 15442 11756
rect 15565 11747 15623 11753
rect 15565 11744 15577 11747
rect 15436 11716 15577 11744
rect 15436 11704 15442 11716
rect 15565 11713 15577 11716
rect 15611 11713 15623 11747
rect 15746 11744 15752 11756
rect 15707 11716 15752 11744
rect 15565 11707 15623 11713
rect 15746 11704 15752 11716
rect 15804 11704 15810 11756
rect 17880 11753 17908 11784
rect 19334 11772 19340 11784
rect 19392 11772 19398 11824
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11744 17187 11747
rect 17865 11747 17923 11753
rect 17865 11744 17877 11747
rect 17175 11716 17877 11744
rect 17175 11713 17187 11716
rect 17129 11707 17187 11713
rect 17865 11713 17877 11716
rect 17911 11713 17923 11747
rect 18782 11744 18788 11756
rect 17865 11707 17923 11713
rect 17972 11716 18788 11744
rect 1762 11676 1768 11688
rect 1723 11648 1768 11676
rect 1762 11636 1768 11648
rect 1820 11636 1826 11688
rect 13265 11679 13323 11685
rect 13265 11645 13277 11679
rect 13311 11645 13323 11679
rect 13265 11639 13323 11645
rect 13280 11608 13308 11639
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 16960 11676 16988 11707
rect 17972 11688 18000 11716
rect 18782 11704 18788 11716
rect 18840 11704 18846 11756
rect 19613 11747 19671 11753
rect 19613 11713 19625 11747
rect 19659 11744 19671 11747
rect 20806 11744 20812 11756
rect 19659 11716 20812 11744
rect 19659 11713 19671 11716
rect 19613 11707 19671 11713
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 17773 11679 17831 11685
rect 17773 11676 17785 11679
rect 13504 11648 13549 11676
rect 16960 11648 17785 11676
rect 13504 11636 13510 11648
rect 17773 11645 17785 11648
rect 17819 11645 17831 11679
rect 17954 11676 17960 11688
rect 17915 11648 17960 11676
rect 17773 11639 17831 11645
rect 17678 11608 17684 11620
rect 13280 11580 17684 11608
rect 17678 11568 17684 11580
rect 17736 11568 17742 11620
rect 17788 11608 17816 11639
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11676 18107 11679
rect 18598 11676 18604 11688
rect 18095 11648 18276 11676
rect 18559 11648 18604 11676
rect 18095 11645 18107 11648
rect 18049 11639 18107 11645
rect 18138 11608 18144 11620
rect 17788 11580 18144 11608
rect 18138 11568 18144 11580
rect 18196 11568 18202 11620
rect 18248 11540 18276 11648
rect 18598 11636 18604 11648
rect 18656 11676 18662 11688
rect 19794 11676 19800 11688
rect 18656 11648 19800 11676
rect 18656 11636 18662 11648
rect 19794 11636 19800 11648
rect 19852 11636 19858 11688
rect 21652 11676 21680 11852
rect 21726 11840 21732 11892
rect 21784 11880 21790 11892
rect 22649 11883 22707 11889
rect 22649 11880 22661 11883
rect 21784 11852 22661 11880
rect 21784 11840 21790 11852
rect 22649 11849 22661 11852
rect 22695 11849 22707 11883
rect 23750 11880 23756 11892
rect 23711 11852 23756 11880
rect 22649 11843 22707 11849
rect 23750 11840 23756 11852
rect 23808 11840 23814 11892
rect 25498 11880 25504 11892
rect 25459 11852 25504 11880
rect 25498 11840 25504 11852
rect 25556 11840 25562 11892
rect 26050 11840 26056 11892
rect 26108 11880 26114 11892
rect 30469 11883 30527 11889
rect 30469 11880 30481 11883
rect 26108 11852 30481 11880
rect 26108 11840 26114 11852
rect 30469 11849 30481 11852
rect 30515 11849 30527 11883
rect 30469 11843 30527 11849
rect 32858 11840 32864 11892
rect 32916 11880 32922 11892
rect 34146 11880 34152 11892
rect 32916 11852 34152 11880
rect 32916 11840 32922 11852
rect 34146 11840 34152 11852
rect 34204 11880 34210 11892
rect 35161 11883 35219 11889
rect 34204 11852 34468 11880
rect 34204 11840 34210 11852
rect 22278 11772 22284 11824
rect 22336 11812 22342 11824
rect 27700 11815 27758 11821
rect 22336 11784 27660 11812
rect 22336 11772 22342 11784
rect 22094 11704 22100 11756
rect 22152 11744 22158 11756
rect 22833 11747 22891 11753
rect 22833 11744 22845 11747
rect 22152 11716 22845 11744
rect 22152 11704 22158 11716
rect 22833 11713 22845 11716
rect 22879 11713 22891 11747
rect 23106 11744 23112 11756
rect 23067 11716 23112 11744
rect 22833 11707 22891 11713
rect 23106 11704 23112 11716
rect 23164 11704 23170 11756
rect 23658 11744 23664 11756
rect 23619 11716 23664 11744
rect 23658 11704 23664 11716
rect 23716 11704 23722 11756
rect 23842 11744 23848 11756
rect 23803 11716 23848 11744
rect 23842 11704 23848 11716
rect 23900 11704 23906 11756
rect 24320 11753 24348 11784
rect 24305 11747 24363 11753
rect 24305 11713 24317 11747
rect 24351 11713 24363 11747
rect 24305 11707 24363 11713
rect 27246 11704 27252 11756
rect 27304 11744 27310 11756
rect 27433 11747 27491 11753
rect 27433 11744 27445 11747
rect 27304 11716 27445 11744
rect 27304 11704 27310 11716
rect 27433 11713 27445 11716
rect 27479 11713 27491 11747
rect 27632 11744 27660 11784
rect 27700 11781 27712 11815
rect 27746 11812 27758 11815
rect 29730 11812 29736 11824
rect 27746 11784 29736 11812
rect 27746 11781 27758 11784
rect 27700 11775 27758 11781
rect 29730 11772 29736 11784
rect 29788 11772 29794 11824
rect 29822 11772 29828 11824
rect 29880 11812 29886 11824
rect 30282 11812 30288 11824
rect 29880 11784 30288 11812
rect 29880 11772 29886 11784
rect 30282 11772 30288 11784
rect 30340 11772 30346 11824
rect 34065 11815 34123 11821
rect 34065 11781 34077 11815
rect 34111 11812 34123 11815
rect 34330 11812 34336 11824
rect 34111 11784 34336 11812
rect 34111 11781 34123 11784
rect 34065 11775 34123 11781
rect 34330 11772 34336 11784
rect 34388 11772 34394 11824
rect 28166 11744 28172 11756
rect 27632 11716 28172 11744
rect 27433 11707 27491 11713
rect 28166 11704 28172 11716
rect 28224 11704 28230 11756
rect 29270 11744 29276 11756
rect 29183 11716 29276 11744
rect 29270 11704 29276 11716
rect 29328 11744 29334 11756
rect 30098 11744 30104 11756
rect 29328 11716 30104 11744
rect 29328 11704 29334 11716
rect 30098 11704 30104 11716
rect 30156 11704 30162 11756
rect 33686 11744 33692 11756
rect 33647 11716 33692 11744
rect 33686 11704 33692 11716
rect 33744 11704 33750 11756
rect 33870 11753 33876 11756
rect 33837 11747 33876 11753
rect 33837 11713 33849 11747
rect 33837 11707 33876 11713
rect 33870 11704 33876 11707
rect 33928 11704 33934 11756
rect 33962 11704 33968 11756
rect 34020 11744 34026 11756
rect 34146 11744 34152 11756
rect 34204 11753 34210 11756
rect 34020 11716 34065 11744
rect 34112 11716 34152 11744
rect 34020 11704 34026 11716
rect 34146 11704 34152 11716
rect 34204 11707 34212 11753
rect 34440 11744 34468 11852
rect 35161 11849 35173 11883
rect 35207 11880 35219 11883
rect 35710 11880 35716 11892
rect 35207 11852 35716 11880
rect 35207 11849 35219 11852
rect 35161 11843 35219 11849
rect 35710 11840 35716 11852
rect 35768 11840 35774 11892
rect 34606 11772 34612 11824
rect 34664 11812 34670 11824
rect 47854 11812 47860 11824
rect 34664 11784 47860 11812
rect 34664 11772 34670 11784
rect 47854 11772 47860 11784
rect 47912 11772 47918 11824
rect 36078 11744 36084 11756
rect 34440 11716 36084 11744
rect 34204 11704 34210 11707
rect 36078 11704 36084 11716
rect 36136 11704 36142 11756
rect 37918 11704 37924 11756
rect 37976 11744 37982 11756
rect 38197 11747 38255 11753
rect 38197 11744 38209 11747
rect 37976 11716 38209 11744
rect 37976 11704 37982 11716
rect 38197 11713 38209 11716
rect 38243 11713 38255 11747
rect 38197 11707 38255 11713
rect 42702 11704 42708 11756
rect 42760 11744 42766 11756
rect 43438 11744 43444 11756
rect 42760 11716 43444 11744
rect 42760 11704 42766 11716
rect 43438 11704 43444 11716
rect 43496 11704 43502 11756
rect 47670 11704 47676 11756
rect 47728 11744 47734 11756
rect 51442 11744 51448 11756
rect 47728 11716 51448 11744
rect 47728 11704 47734 11716
rect 51442 11704 51448 11716
rect 51500 11704 51506 11756
rect 57146 11744 57152 11756
rect 57107 11716 57152 11744
rect 57146 11704 57152 11716
rect 57204 11704 57210 11756
rect 22925 11679 22983 11685
rect 21652 11648 21956 11676
rect 18322 11568 18328 11620
rect 18380 11608 18386 11620
rect 18877 11611 18935 11617
rect 18877 11608 18889 11611
rect 18380 11580 18889 11608
rect 18380 11568 18386 11580
rect 18877 11577 18889 11580
rect 18923 11577 18935 11611
rect 19978 11608 19984 11620
rect 18877 11571 18935 11577
rect 18984 11580 19984 11608
rect 18984 11540 19012 11580
rect 19978 11568 19984 11580
rect 20036 11568 20042 11620
rect 21818 11608 21824 11620
rect 20088 11580 21824 11608
rect 18248 11512 19012 11540
rect 19058 11500 19064 11552
rect 19116 11540 19122 11552
rect 20088 11540 20116 11580
rect 21818 11568 21824 11580
rect 21876 11568 21882 11620
rect 21928 11608 21956 11648
rect 22925 11645 22937 11679
rect 22971 11645 22983 11679
rect 22925 11639 22983 11645
rect 22940 11608 22968 11639
rect 23014 11636 23020 11688
rect 23072 11676 23078 11688
rect 23072 11648 23117 11676
rect 23072 11636 23078 11648
rect 34054 11636 34060 11688
rect 34112 11676 34118 11688
rect 35253 11679 35311 11685
rect 35253 11676 35265 11679
rect 34112 11648 35265 11676
rect 34112 11636 34118 11648
rect 35253 11645 35265 11648
rect 35299 11645 35311 11679
rect 35253 11639 35311 11645
rect 35345 11679 35403 11685
rect 35345 11645 35357 11679
rect 35391 11676 35403 11679
rect 38378 11676 38384 11688
rect 35391 11648 38384 11676
rect 35391 11645 35403 11648
rect 35345 11639 35403 11645
rect 25590 11608 25596 11620
rect 21928 11580 25596 11608
rect 25590 11568 25596 11580
rect 25648 11568 25654 11620
rect 28442 11568 28448 11620
rect 28500 11608 28506 11620
rect 33962 11608 33968 11620
rect 28500 11580 33968 11608
rect 28500 11568 28506 11580
rect 33962 11568 33968 11580
rect 34020 11568 34026 11620
rect 34606 11568 34612 11620
rect 34664 11608 34670 11620
rect 35360 11608 35388 11639
rect 38378 11636 38384 11648
rect 38436 11636 38442 11688
rect 34664 11580 35388 11608
rect 34664 11568 34670 11580
rect 19116 11512 20116 11540
rect 19116 11500 19122 11512
rect 21726 11500 21732 11552
rect 21784 11540 21790 11552
rect 28813 11543 28871 11549
rect 28813 11540 28825 11543
rect 21784 11512 28825 11540
rect 21784 11500 21790 11512
rect 28813 11509 28825 11512
rect 28859 11540 28871 11543
rect 30190 11540 30196 11552
rect 28859 11512 30196 11540
rect 28859 11509 28871 11512
rect 28813 11503 28871 11509
rect 30190 11500 30196 11512
rect 30248 11500 30254 11552
rect 34330 11500 34336 11552
rect 34388 11540 34394 11552
rect 34790 11540 34796 11552
rect 34388 11512 34433 11540
rect 34751 11512 34796 11540
rect 34388 11500 34394 11512
rect 34790 11500 34796 11512
rect 34848 11500 34854 11552
rect 57238 11540 57244 11552
rect 57199 11512 57244 11540
rect 57238 11500 57244 11512
rect 57296 11500 57302 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 13449 11339 13507 11345
rect 13449 11305 13461 11339
rect 13495 11336 13507 11339
rect 13538 11336 13544 11348
rect 13495 11308 13544 11336
rect 13495 11305 13507 11308
rect 13449 11299 13507 11305
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 17678 11296 17684 11348
rect 17736 11336 17742 11348
rect 17736 11308 20392 11336
rect 17736 11296 17742 11308
rect 9122 11228 9128 11280
rect 9180 11268 9186 11280
rect 13265 11271 13323 11277
rect 13265 11268 13277 11271
rect 9180 11240 13277 11268
rect 9180 11228 9186 11240
rect 13265 11237 13277 11240
rect 13311 11237 13323 11271
rect 13265 11231 13323 11237
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 19426 11268 19432 11280
rect 16264 11240 19432 11268
rect 16264 11228 16270 11240
rect 19426 11228 19432 11240
rect 19484 11228 19490 11280
rect 20364 11268 20392 11308
rect 20438 11296 20444 11348
rect 20496 11336 20502 11348
rect 20622 11336 20628 11348
rect 20496 11308 20628 11336
rect 20496 11296 20502 11308
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 20806 11336 20812 11348
rect 20767 11308 20812 11336
rect 20806 11296 20812 11308
rect 20864 11296 20870 11348
rect 21266 11336 21272 11348
rect 21227 11308 21272 11336
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 22554 11296 22560 11348
rect 22612 11296 22618 11348
rect 23017 11339 23075 11345
rect 23017 11305 23029 11339
rect 23063 11336 23075 11339
rect 23842 11336 23848 11348
rect 23063 11308 23848 11336
rect 23063 11305 23075 11308
rect 23017 11299 23075 11305
rect 23842 11296 23848 11308
rect 23900 11296 23906 11348
rect 24578 11336 24584 11348
rect 24539 11308 24584 11336
rect 24578 11296 24584 11308
rect 24636 11296 24642 11348
rect 25498 11296 25504 11348
rect 25556 11336 25562 11348
rect 25556 11308 28948 11336
rect 25556 11296 25562 11308
rect 21450 11268 21456 11280
rect 20364 11240 21456 11268
rect 21450 11228 21456 11240
rect 21508 11228 21514 11280
rect 12802 11160 12808 11212
rect 12860 11200 12866 11212
rect 17126 11200 17132 11212
rect 12860 11172 17132 11200
rect 12860 11160 12866 11172
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 18138 11160 18144 11212
rect 18196 11200 18202 11212
rect 18233 11203 18291 11209
rect 18233 11200 18245 11203
rect 18196 11172 18245 11200
rect 18196 11160 18202 11172
rect 18233 11169 18245 11172
rect 18279 11200 18291 11203
rect 19150 11200 19156 11212
rect 18279 11172 19156 11200
rect 18279 11169 18291 11172
rect 18233 11163 18291 11169
rect 19150 11160 19156 11172
rect 19208 11160 19214 11212
rect 21729 11203 21787 11209
rect 21729 11200 21741 11203
rect 20824 11172 21741 11200
rect 14826 11092 14832 11144
rect 14884 11132 14890 11144
rect 16022 11132 16028 11144
rect 14884 11104 16028 11132
rect 14884 11092 14890 11104
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11132 18015 11135
rect 18598 11132 18604 11144
rect 18003 11104 18604 11132
rect 18003 11101 18015 11104
rect 17957 11095 18015 11101
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 19426 11132 19432 11144
rect 19339 11104 19432 11132
rect 19426 11092 19432 11104
rect 19484 11132 19490 11144
rect 20622 11132 20628 11144
rect 19484 11104 20628 11132
rect 19484 11092 19490 11104
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 12989 11067 13047 11073
rect 12989 11033 13001 11067
rect 13035 11064 13047 11067
rect 17494 11064 17500 11076
rect 13035 11036 17500 11064
rect 13035 11033 13047 11036
rect 12989 11027 13047 11033
rect 17494 11024 17500 11036
rect 17552 11024 17558 11076
rect 19674 11067 19732 11073
rect 19674 11064 19686 11067
rect 17604 11036 19686 11064
rect 17604 11005 17632 11036
rect 19674 11033 19686 11036
rect 19720 11033 19732 11067
rect 19674 11027 19732 11033
rect 20346 11024 20352 11076
rect 20404 11064 20410 11076
rect 20824 11064 20852 11172
rect 21729 11169 21741 11172
rect 21775 11169 21787 11203
rect 21729 11163 21787 11169
rect 21913 11203 21971 11209
rect 21913 11169 21925 11203
rect 21959 11200 21971 11203
rect 22572 11200 22600 11296
rect 22649 11203 22707 11209
rect 22649 11200 22661 11203
rect 21959 11172 22094 11200
rect 22572 11172 22661 11200
rect 21959 11169 21971 11172
rect 21913 11163 21971 11169
rect 20898 11092 20904 11144
rect 20956 11132 20962 11144
rect 21450 11132 21456 11144
rect 20956 11104 21456 11132
rect 20956 11092 20962 11104
rect 21450 11092 21456 11104
rect 21508 11132 21514 11144
rect 21637 11135 21695 11141
rect 21637 11132 21649 11135
rect 21508 11104 21649 11132
rect 21508 11092 21514 11104
rect 21637 11101 21649 11104
rect 21683 11101 21695 11135
rect 22066 11132 22094 11172
rect 22649 11169 22661 11172
rect 22695 11169 22707 11203
rect 22649 11163 22707 11169
rect 26418 11160 26424 11212
rect 26476 11200 26482 11212
rect 28920 11209 28948 11308
rect 33226 11296 33232 11348
rect 33284 11336 33290 11348
rect 33686 11336 33692 11348
rect 33284 11308 33692 11336
rect 33284 11296 33290 11308
rect 33686 11296 33692 11308
rect 33744 11296 33750 11348
rect 34054 11296 34060 11348
rect 34112 11336 34118 11348
rect 36265 11339 36323 11345
rect 36265 11336 36277 11339
rect 34112 11308 36277 11336
rect 34112 11296 34118 11308
rect 36265 11305 36277 11308
rect 36311 11305 36323 11339
rect 58250 11336 58256 11348
rect 58211 11308 58256 11336
rect 36265 11299 36323 11305
rect 58250 11296 58256 11308
rect 58308 11296 58314 11348
rect 32582 11228 32588 11280
rect 32640 11268 32646 11280
rect 34606 11268 34612 11280
rect 32640 11240 34612 11268
rect 32640 11228 32646 11240
rect 28905 11203 28963 11209
rect 26476 11172 28580 11200
rect 26476 11160 26482 11172
rect 22554 11132 22560 11144
rect 22066 11104 22560 11132
rect 21637 11095 21695 11101
rect 22554 11092 22560 11104
rect 22612 11092 22618 11144
rect 22833 11135 22891 11141
rect 22833 11101 22845 11135
rect 22879 11132 22891 11135
rect 23290 11132 23296 11144
rect 22879 11104 23296 11132
rect 22879 11101 22891 11104
rect 22833 11095 22891 11101
rect 23290 11092 23296 11104
rect 23348 11092 23354 11144
rect 23382 11092 23388 11144
rect 23440 11132 23446 11144
rect 24210 11132 24216 11144
rect 23440 11104 24216 11132
rect 23440 11092 23446 11104
rect 24210 11092 24216 11104
rect 24268 11092 24274 11144
rect 24581 11135 24639 11141
rect 24581 11101 24593 11135
rect 24627 11132 24639 11135
rect 24670 11132 24676 11144
rect 24627 11104 24676 11132
rect 24627 11101 24639 11104
rect 24581 11095 24639 11101
rect 24670 11092 24676 11104
rect 24728 11092 24734 11144
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11101 24823 11135
rect 25590 11132 25596 11144
rect 25503 11104 25596 11132
rect 24765 11095 24823 11101
rect 20404 11036 20852 11064
rect 20404 11024 20410 11036
rect 20990 11024 20996 11076
rect 21048 11064 21054 11076
rect 24780 11064 24808 11095
rect 25590 11092 25596 11104
rect 25648 11132 25654 11144
rect 28442 11132 28448 11144
rect 25648 11104 28448 11132
rect 25648 11092 25654 11104
rect 28442 11092 28448 11104
rect 28500 11092 28506 11144
rect 28552 11132 28580 11172
rect 28905 11169 28917 11203
rect 28951 11169 28963 11203
rect 28905 11163 28963 11169
rect 28994 11160 29000 11212
rect 29052 11200 29058 11212
rect 34054 11200 34060 11212
rect 29052 11172 34060 11200
rect 29052 11160 29058 11172
rect 34054 11160 34060 11172
rect 34112 11160 34118 11212
rect 34256 11209 34284 11240
rect 34606 11228 34612 11240
rect 34664 11228 34670 11280
rect 34241 11203 34299 11209
rect 34241 11169 34253 11203
rect 34287 11169 34299 11203
rect 34241 11163 34299 11169
rect 34790 11160 34796 11212
rect 34848 11200 34854 11212
rect 34848 11172 35020 11200
rect 34848 11160 34854 11172
rect 32953 11135 33011 11141
rect 32953 11132 32965 11135
rect 28552 11104 32965 11132
rect 32953 11101 32965 11104
rect 32999 11101 33011 11135
rect 32953 11095 33011 11101
rect 33226 11092 33232 11144
rect 33284 11132 33290 11144
rect 34882 11132 34888 11144
rect 33284 11104 33916 11132
rect 34843 11104 34888 11132
rect 33284 11092 33290 11104
rect 21048 11036 24808 11064
rect 21048 11024 21054 11036
rect 28258 11024 28264 11076
rect 28316 11064 28322 11076
rect 28813 11067 28871 11073
rect 28813 11064 28825 11067
rect 28316 11036 28825 11064
rect 28316 11024 28322 11036
rect 28813 11033 28825 11036
rect 28859 11064 28871 11067
rect 29454 11064 29460 11076
rect 28859 11036 29460 11064
rect 28859 11033 28871 11036
rect 28813 11027 28871 11033
rect 29454 11024 29460 11036
rect 29512 11024 29518 11076
rect 32398 11064 32404 11076
rect 32359 11036 32404 11064
rect 32398 11024 32404 11036
rect 32456 11024 32462 11076
rect 32582 11064 32588 11076
rect 32543 11036 32588 11064
rect 32582 11024 32588 11036
rect 32640 11024 32646 11076
rect 32687 11067 32745 11073
rect 32687 11033 32699 11067
rect 32733 11064 32745 11067
rect 33778 11064 33784 11076
rect 32733 11036 33784 11064
rect 32733 11033 32745 11036
rect 32687 11027 32745 11033
rect 33778 11024 33784 11036
rect 33836 11024 33842 11076
rect 33888 11064 33916 11104
rect 34882 11092 34888 11104
rect 34940 11092 34946 11144
rect 34992 11132 35020 11172
rect 36538 11160 36544 11212
rect 36596 11200 36602 11212
rect 36998 11200 37004 11212
rect 36596 11172 37004 11200
rect 36596 11160 36602 11172
rect 36998 11160 37004 11172
rect 37056 11160 37062 11212
rect 37918 11160 37924 11212
rect 37976 11200 37982 11212
rect 38657 11203 38715 11209
rect 38657 11200 38669 11203
rect 37976 11172 38669 11200
rect 37976 11160 37982 11172
rect 38657 11169 38669 11172
rect 38703 11169 38715 11203
rect 56870 11200 56876 11212
rect 56831 11172 56876 11200
rect 38657 11163 38715 11169
rect 56870 11160 56876 11172
rect 56928 11160 56934 11212
rect 35141 11135 35199 11141
rect 35141 11132 35153 11135
rect 34992 11104 35153 11132
rect 35141 11101 35153 11104
rect 35187 11101 35199 11135
rect 35141 11095 35199 11101
rect 36630 11092 36636 11144
rect 36688 11132 36694 11144
rect 36725 11135 36783 11141
rect 36725 11132 36737 11135
rect 36688 11104 36737 11132
rect 36688 11092 36694 11104
rect 36725 11101 36737 11104
rect 36771 11132 36783 11135
rect 38381 11135 38439 11141
rect 36771 11104 38240 11132
rect 36771 11101 36783 11104
rect 36725 11095 36783 11101
rect 34057 11067 34115 11073
rect 34057 11064 34069 11067
rect 33888 11036 34069 11064
rect 34057 11033 34069 11036
rect 34103 11033 34115 11067
rect 34057 11027 34115 11033
rect 34146 11024 34152 11076
rect 34204 11064 34210 11076
rect 34606 11064 34612 11076
rect 34204 11036 34612 11064
rect 34204 11024 34210 11036
rect 34606 11024 34612 11036
rect 34664 11024 34670 11076
rect 35894 11024 35900 11076
rect 35952 11064 35958 11076
rect 37461 11067 37519 11073
rect 37461 11064 37473 11067
rect 35952 11036 37473 11064
rect 35952 11024 35958 11036
rect 37461 11033 37473 11036
rect 37507 11033 37519 11067
rect 38212 11064 38240 11104
rect 38381 11101 38393 11135
rect 38427 11132 38439 11135
rect 39114 11132 39120 11144
rect 38427 11104 39120 11132
rect 38427 11101 38439 11104
rect 38381 11095 38439 11101
rect 39114 11092 39120 11104
rect 39172 11092 39178 11144
rect 40402 11064 40408 11076
rect 38212 11036 40408 11064
rect 37461 11027 37519 11033
rect 40402 11024 40408 11036
rect 40460 11024 40466 11076
rect 56778 11024 56784 11076
rect 56836 11064 56842 11076
rect 57118 11067 57176 11073
rect 57118 11064 57130 11067
rect 56836 11036 57130 11064
rect 56836 11024 56842 11036
rect 57118 11033 57130 11036
rect 57164 11033 57176 11067
rect 57118 11027 57176 11033
rect 17589 10999 17647 11005
rect 17589 10965 17601 10999
rect 17635 10965 17647 10999
rect 17589 10959 17647 10965
rect 18046 10956 18052 11008
rect 18104 10996 18110 11008
rect 18104 10968 18149 10996
rect 18104 10956 18110 10968
rect 19978 10956 19984 11008
rect 20036 10996 20042 11008
rect 25774 10996 25780 11008
rect 20036 10968 25780 10996
rect 20036 10956 20042 10968
rect 25774 10956 25780 10968
rect 25832 10956 25838 11008
rect 25866 10956 25872 11008
rect 25924 10996 25930 11008
rect 26789 10999 26847 11005
rect 26789 10996 26801 10999
rect 25924 10968 26801 10996
rect 25924 10956 25930 10968
rect 26789 10965 26801 10968
rect 26835 10965 26847 10999
rect 28350 10996 28356 11008
rect 28311 10968 28356 10996
rect 26789 10959 26847 10965
rect 28350 10956 28356 10968
rect 28408 10956 28414 11008
rect 28721 10999 28779 11005
rect 28721 10965 28733 10999
rect 28767 10996 28779 10999
rect 29086 10996 29092 11008
rect 28767 10968 29092 10996
rect 28767 10965 28779 10968
rect 28721 10959 28779 10965
rect 29086 10956 29092 10968
rect 29144 10956 29150 11008
rect 32766 10996 32772 11008
rect 32727 10968 32772 10996
rect 32766 10956 32772 10968
rect 32824 10956 32830 11008
rect 33597 10999 33655 11005
rect 33597 10965 33609 10999
rect 33643 10996 33655 10999
rect 33870 10996 33876 11008
rect 33643 10968 33876 10996
rect 33643 10965 33655 10968
rect 33597 10959 33655 10965
rect 33870 10956 33876 10968
rect 33928 10956 33934 11008
rect 33965 10999 34023 11005
rect 33965 10965 33977 10999
rect 34011 10996 34023 10999
rect 36446 10996 36452 11008
rect 34011 10968 36452 10996
rect 34011 10965 34023 10968
rect 33965 10959 34023 10965
rect 36446 10956 36452 10968
rect 36504 10956 36510 11008
rect 40126 10956 40132 11008
rect 40184 10996 40190 11008
rect 41690 10996 41696 11008
rect 40184 10968 41696 10996
rect 40184 10956 40190 10968
rect 41690 10956 41696 10968
rect 41748 10956 41754 11008
rect 49234 10956 49240 11008
rect 49292 10996 49298 11008
rect 51258 10996 51264 11008
rect 49292 10968 51264 10996
rect 49292 10956 49298 10968
rect 51258 10956 51264 10968
rect 51316 10956 51322 11008
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 14737 10795 14795 10801
rect 14737 10792 14749 10795
rect 11112 10764 14749 10792
rect 11112 10752 11118 10764
rect 14737 10761 14749 10764
rect 14783 10761 14795 10795
rect 21450 10792 21456 10804
rect 14737 10755 14795 10761
rect 16592 10764 20760 10792
rect 21411 10764 21456 10792
rect 16592 10724 16620 10764
rect 2746 10696 16620 10724
rect 1581 10659 1639 10665
rect 1581 10625 1593 10659
rect 1627 10656 1639 10659
rect 2409 10659 2467 10665
rect 2409 10656 2421 10659
rect 1627 10628 2421 10656
rect 1627 10625 1639 10628
rect 1581 10619 1639 10625
rect 2409 10625 2421 10628
rect 2455 10656 2467 10659
rect 2746 10656 2774 10696
rect 17126 10684 17132 10736
rect 17184 10724 17190 10736
rect 17184 10696 17908 10724
rect 17184 10684 17190 10696
rect 13078 10656 13084 10668
rect 2455 10628 2774 10656
rect 13039 10628 13084 10656
rect 2455 10625 2467 10628
rect 2409 10619 2467 10625
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 13265 10659 13323 10665
rect 13265 10625 13277 10659
rect 13311 10656 13323 10659
rect 13998 10656 14004 10668
rect 13311 10628 14004 10656
rect 13311 10625 13323 10628
rect 13265 10619 13323 10625
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 17681 10659 17739 10665
rect 17681 10656 17693 10659
rect 14108 10628 15424 10656
rect 1762 10588 1768 10600
rect 1723 10560 1768 10588
rect 1762 10548 1768 10560
rect 1820 10548 1826 10600
rect 12986 10548 12992 10600
rect 13044 10588 13050 10600
rect 13173 10591 13231 10597
rect 13173 10588 13185 10591
rect 13044 10560 13185 10588
rect 13044 10548 13050 10560
rect 13173 10557 13185 10560
rect 13219 10557 13231 10591
rect 13173 10551 13231 10557
rect 13354 10548 13360 10600
rect 13412 10588 13418 10600
rect 13412 10560 13457 10588
rect 13412 10548 13418 10560
rect 5994 10480 6000 10532
rect 6052 10520 6058 10532
rect 14108 10520 14136 10628
rect 14918 10588 14924 10600
rect 14879 10560 14924 10588
rect 14918 10548 14924 10560
rect 14976 10548 14982 10600
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 15105 10591 15163 10597
rect 15105 10557 15117 10591
rect 15151 10557 15163 10591
rect 15105 10551 15163 10557
rect 6052 10492 14136 10520
rect 6052 10480 6058 10492
rect 12894 10452 12900 10464
rect 12855 10424 12900 10452
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 15028 10452 15056 10551
rect 15120 10520 15148 10551
rect 15194 10548 15200 10600
rect 15252 10588 15258 10600
rect 15396 10588 15424 10628
rect 17328 10628 17693 10656
rect 17328 10588 17356 10628
rect 17681 10625 17693 10628
rect 17727 10625 17739 10659
rect 17681 10619 17739 10625
rect 17770 10588 17776 10600
rect 15252 10560 15297 10588
rect 15396 10560 17356 10588
rect 17731 10560 17776 10588
rect 15252 10548 15258 10560
rect 17770 10548 17776 10560
rect 17828 10548 17834 10600
rect 17880 10597 17908 10696
rect 18506 10684 18512 10736
rect 18564 10724 18570 10736
rect 18874 10724 18880 10736
rect 18564 10696 18880 10724
rect 18564 10684 18570 10696
rect 18874 10684 18880 10696
rect 18932 10684 18938 10736
rect 20622 10724 20628 10736
rect 20088 10696 20628 10724
rect 20088 10665 20116 10696
rect 20622 10684 20628 10696
rect 20680 10684 20686 10736
rect 20732 10724 20760 10764
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 21634 10752 21640 10804
rect 21692 10792 21698 10804
rect 21910 10792 21916 10804
rect 21692 10764 21916 10792
rect 21692 10752 21698 10764
rect 21910 10752 21916 10764
rect 21968 10792 21974 10804
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 21968 10764 22385 10792
rect 21968 10752 21974 10764
rect 22373 10761 22385 10764
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 23584 10764 28488 10792
rect 23584 10724 23612 10764
rect 24578 10724 24584 10736
rect 20732 10696 23612 10724
rect 23676 10696 24584 10724
rect 20073 10659 20131 10665
rect 20073 10625 20085 10659
rect 20119 10625 20131 10659
rect 20073 10619 20131 10625
rect 20340 10659 20398 10665
rect 20340 10625 20352 10659
rect 20386 10656 20398 10659
rect 21266 10656 21272 10668
rect 20386 10628 21272 10656
rect 20386 10625 20398 10628
rect 20340 10619 20398 10625
rect 21266 10616 21272 10628
rect 21324 10616 21330 10668
rect 21634 10656 21640 10668
rect 21376 10628 21640 10656
rect 17865 10591 17923 10597
rect 17865 10557 17877 10591
rect 17911 10588 17923 10591
rect 18506 10588 18512 10600
rect 17911 10560 18512 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 18506 10548 18512 10560
rect 18564 10548 18570 10600
rect 21376 10588 21404 10628
rect 21634 10616 21640 10628
rect 21692 10616 21698 10668
rect 22278 10616 22284 10668
rect 22336 10656 22342 10668
rect 22830 10656 22836 10668
rect 22336 10628 22836 10656
rect 22336 10616 22342 10628
rect 22830 10616 22836 10628
rect 22888 10616 22894 10668
rect 23676 10665 23704 10696
rect 24578 10684 24584 10696
rect 24636 10724 24642 10736
rect 24636 10696 27200 10724
rect 24636 10684 24642 10696
rect 23934 10665 23940 10668
rect 23661 10659 23719 10665
rect 23661 10625 23673 10659
rect 23707 10625 23719 10659
rect 23928 10656 23940 10665
rect 23895 10628 23940 10656
rect 23661 10619 23719 10625
rect 23928 10619 23940 10628
rect 23934 10616 23940 10619
rect 23992 10616 23998 10668
rect 27172 10665 27200 10696
rect 26421 10659 26479 10665
rect 26421 10625 26433 10659
rect 26467 10625 26479 10659
rect 26421 10619 26479 10625
rect 27157 10659 27215 10665
rect 27157 10625 27169 10659
rect 27203 10625 27215 10659
rect 28350 10656 28356 10668
rect 27157 10619 27215 10625
rect 27264 10628 28356 10656
rect 21192 10560 21404 10588
rect 17126 10520 17132 10532
rect 15120 10492 17132 10520
rect 17126 10480 17132 10492
rect 17184 10480 17190 10532
rect 17313 10523 17371 10529
rect 17313 10489 17325 10523
rect 17359 10520 17371 10523
rect 18046 10520 18052 10532
rect 17359 10492 18052 10520
rect 17359 10489 17371 10492
rect 17313 10483 17371 10489
rect 18046 10480 18052 10492
rect 18104 10480 18110 10532
rect 21192 10452 21220 10560
rect 21450 10548 21456 10600
rect 21508 10588 21514 10600
rect 22002 10588 22008 10600
rect 21508 10560 22008 10588
rect 21508 10548 21514 10560
rect 22002 10548 22008 10560
rect 22060 10548 22066 10600
rect 22186 10548 22192 10600
rect 22244 10588 22250 10600
rect 22465 10591 22523 10597
rect 22465 10588 22477 10591
rect 22244 10560 22477 10588
rect 22244 10548 22250 10560
rect 22465 10557 22477 10560
rect 22511 10557 22523 10591
rect 22646 10588 22652 10600
rect 22607 10560 22652 10588
rect 22465 10551 22523 10557
rect 22646 10548 22652 10560
rect 22704 10548 22710 10600
rect 26237 10591 26295 10597
rect 26237 10557 26249 10591
rect 26283 10557 26295 10591
rect 26436 10588 26464 10619
rect 27264 10588 27292 10628
rect 28350 10616 28356 10628
rect 28408 10616 28414 10668
rect 27430 10588 27436 10600
rect 26436 10560 27292 10588
rect 27391 10560 27436 10588
rect 26237 10551 26295 10557
rect 21542 10480 21548 10532
rect 21600 10520 21606 10532
rect 26252 10520 26280 10551
rect 27430 10548 27436 10560
rect 27488 10548 27494 10600
rect 28460 10588 28488 10764
rect 28534 10752 28540 10804
rect 28592 10792 28598 10804
rect 47670 10792 47676 10804
rect 28592 10764 35020 10792
rect 28592 10752 28598 10764
rect 28626 10684 28632 10736
rect 28684 10724 28690 10736
rect 33778 10724 33784 10736
rect 28684 10696 33784 10724
rect 28684 10684 28690 10696
rect 33778 10684 33784 10696
rect 33836 10684 33842 10736
rect 34882 10724 34888 10736
rect 33888 10696 34888 10724
rect 29270 10656 29276 10668
rect 29231 10628 29276 10656
rect 29270 10616 29276 10628
rect 29328 10616 29334 10668
rect 29454 10656 29460 10668
rect 29415 10628 29460 10656
rect 29454 10616 29460 10628
rect 29512 10616 29518 10668
rect 30926 10616 30932 10668
rect 30984 10656 30990 10668
rect 33888 10665 33916 10696
rect 34882 10684 34888 10696
rect 34940 10684 34946 10736
rect 33873 10659 33931 10665
rect 33873 10656 33885 10659
rect 30984 10628 33885 10656
rect 30984 10616 30990 10628
rect 33873 10625 33885 10628
rect 33919 10625 33931 10659
rect 33873 10619 33931 10625
rect 33962 10616 33968 10668
rect 34020 10656 34026 10668
rect 34129 10659 34187 10665
rect 34129 10656 34141 10659
rect 34020 10628 34141 10656
rect 34020 10616 34026 10628
rect 34129 10625 34141 10628
rect 34175 10625 34187 10659
rect 34129 10619 34187 10625
rect 28460 10560 31754 10588
rect 26970 10520 26976 10532
rect 21600 10492 23704 10520
rect 26252 10492 26976 10520
rect 21600 10480 21606 10492
rect 15028 10424 21220 10452
rect 21266 10412 21272 10464
rect 21324 10452 21330 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21324 10424 22017 10452
rect 21324 10412 21330 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 23676 10452 23704 10492
rect 26970 10480 26976 10492
rect 27028 10480 27034 10532
rect 28166 10480 28172 10532
rect 28224 10520 28230 10532
rect 28537 10523 28595 10529
rect 28537 10520 28549 10523
rect 28224 10492 28549 10520
rect 28224 10480 28230 10492
rect 28537 10489 28549 10492
rect 28583 10489 28595 10523
rect 31726 10520 31754 10560
rect 32398 10520 32404 10532
rect 31726 10492 32404 10520
rect 28537 10483 28595 10489
rect 32398 10480 32404 10492
rect 32456 10480 32462 10532
rect 34992 10520 35020 10764
rect 35728 10764 47676 10792
rect 35728 10665 35756 10764
rect 47670 10752 47676 10764
rect 47728 10752 47734 10804
rect 57146 10792 57152 10804
rect 56796 10764 57152 10792
rect 35986 10724 35992 10736
rect 35947 10696 35992 10724
rect 35986 10684 35992 10696
rect 36044 10684 36050 10736
rect 56594 10684 56600 10736
rect 56652 10724 56658 10736
rect 56796 10733 56824 10764
rect 57146 10752 57152 10764
rect 57204 10752 57210 10804
rect 56781 10727 56839 10733
rect 56781 10724 56793 10727
rect 56652 10696 56793 10724
rect 56652 10684 56658 10696
rect 56781 10693 56793 10696
rect 56827 10693 56839 10727
rect 56781 10687 56839 10693
rect 56965 10727 57023 10733
rect 56965 10693 56977 10727
rect 57011 10724 57023 10727
rect 58161 10727 58219 10733
rect 58161 10724 58173 10727
rect 57011 10696 58173 10724
rect 57011 10693 57023 10696
rect 56965 10687 57023 10693
rect 58161 10693 58173 10696
rect 58207 10693 58219 10727
rect 58161 10687 58219 10693
rect 35713 10659 35771 10665
rect 35713 10625 35725 10659
rect 35759 10625 35771 10659
rect 35894 10656 35900 10668
rect 35855 10628 35900 10656
rect 35713 10619 35771 10625
rect 35894 10616 35900 10628
rect 35952 10616 35958 10668
rect 36078 10656 36084 10668
rect 36039 10628 36084 10656
rect 36078 10616 36084 10628
rect 36136 10616 36142 10668
rect 37734 10665 37740 10668
rect 37728 10619 37740 10665
rect 37792 10656 37798 10668
rect 57057 10659 57115 10665
rect 37792 10628 37828 10656
rect 37734 10616 37740 10619
rect 37792 10616 37798 10628
rect 57057 10625 57069 10659
rect 57103 10625 57115 10659
rect 57057 10619 57115 10625
rect 35066 10548 35072 10600
rect 35124 10588 35130 10600
rect 37461 10591 37519 10597
rect 37461 10588 37473 10591
rect 35124 10560 37473 10588
rect 35124 10548 35130 10560
rect 37461 10557 37473 10560
rect 37507 10557 37519 10591
rect 37461 10551 37519 10557
rect 56594 10548 56600 10600
rect 56652 10588 56658 10600
rect 57072 10588 57100 10619
rect 57882 10616 57888 10668
rect 57940 10656 57946 10668
rect 58069 10659 58127 10665
rect 58069 10656 58081 10659
rect 57940 10628 58081 10656
rect 57940 10616 57946 10628
rect 58069 10625 58081 10628
rect 58115 10625 58127 10659
rect 58250 10656 58256 10668
rect 58211 10628 58256 10656
rect 58069 10619 58127 10625
rect 58250 10616 58256 10628
rect 58308 10616 58314 10668
rect 56652 10560 57100 10588
rect 56652 10548 56658 10560
rect 36814 10520 36820 10532
rect 34992 10492 36820 10520
rect 36814 10480 36820 10492
rect 36872 10480 36878 10532
rect 56778 10520 56784 10532
rect 56739 10492 56784 10520
rect 56778 10480 56784 10492
rect 56836 10480 56842 10532
rect 23842 10452 23848 10464
rect 23676 10424 23848 10452
rect 22005 10415 22063 10421
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 25038 10452 25044 10464
rect 24999 10424 25044 10452
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 26602 10452 26608 10464
rect 26563 10424 26608 10452
rect 26602 10412 26608 10424
rect 26660 10412 26666 10464
rect 26786 10412 26792 10464
rect 26844 10452 26850 10464
rect 29086 10452 29092 10464
rect 26844 10424 29092 10452
rect 26844 10412 26850 10424
rect 29086 10412 29092 10424
rect 29144 10412 29150 10464
rect 29362 10452 29368 10464
rect 29323 10424 29368 10452
rect 29362 10412 29368 10424
rect 29420 10412 29426 10464
rect 29730 10412 29736 10464
rect 29788 10452 29794 10464
rect 32306 10452 32312 10464
rect 29788 10424 32312 10452
rect 29788 10412 29794 10424
rect 32306 10412 32312 10424
rect 32364 10412 32370 10464
rect 33226 10412 33232 10464
rect 33284 10452 33290 10464
rect 35253 10455 35311 10461
rect 35253 10452 35265 10455
rect 33284 10424 35265 10452
rect 33284 10412 33290 10424
rect 35253 10421 35265 10424
rect 35299 10421 35311 10455
rect 36262 10452 36268 10464
rect 36223 10424 36268 10452
rect 35253 10415 35311 10421
rect 36262 10412 36268 10424
rect 36320 10412 36326 10464
rect 38838 10452 38844 10464
rect 38799 10424 38844 10452
rect 38838 10412 38844 10424
rect 38896 10412 38902 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 13265 10251 13323 10257
rect 13265 10217 13277 10251
rect 13311 10248 13323 10251
rect 13446 10248 13452 10260
rect 13311 10220 13452 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 17770 10208 17776 10260
rect 17828 10248 17834 10260
rect 21542 10248 21548 10260
rect 17828 10220 21548 10248
rect 17828 10208 17834 10220
rect 21542 10208 21548 10220
rect 21600 10208 21606 10260
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 22060 10208 22094 10248
rect 22646 10208 22652 10260
rect 22704 10248 22710 10260
rect 23937 10251 23995 10257
rect 23937 10248 23949 10251
rect 22704 10220 23949 10248
rect 22704 10208 22710 10220
rect 23937 10217 23949 10220
rect 23983 10217 23995 10251
rect 25774 10248 25780 10260
rect 23937 10211 23995 10217
rect 24044 10220 24808 10248
rect 25735 10220 25780 10248
rect 8938 10140 8944 10192
rect 8996 10180 9002 10192
rect 13081 10183 13139 10189
rect 13081 10180 13093 10183
rect 8996 10152 13093 10180
rect 8996 10140 9002 10152
rect 13081 10149 13093 10152
rect 13127 10149 13139 10183
rect 13081 10143 13139 10149
rect 14553 10183 14611 10189
rect 14553 10149 14565 10183
rect 14599 10149 14611 10183
rect 14553 10143 14611 10149
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 14568 10112 14596 10143
rect 14918 10140 14924 10192
rect 14976 10180 14982 10192
rect 20070 10180 20076 10192
rect 14976 10152 20076 10180
rect 14976 10140 14982 10152
rect 20070 10140 20076 10152
rect 20128 10140 20134 10192
rect 21910 10180 21916 10192
rect 21871 10152 21916 10180
rect 21910 10140 21916 10152
rect 21968 10140 21974 10192
rect 22066 10180 22094 10208
rect 24044 10180 24072 10220
rect 22066 10152 24072 10180
rect 24780 10180 24808 10220
rect 25774 10208 25780 10220
rect 25832 10208 25838 10260
rect 28626 10248 28632 10260
rect 25884 10220 28632 10248
rect 25884 10180 25912 10220
rect 28626 10208 28632 10220
rect 28684 10208 28690 10260
rect 30466 10248 30472 10260
rect 29104 10220 30472 10248
rect 24780 10152 25912 10180
rect 8444 10084 14596 10112
rect 8444 10072 8450 10084
rect 22462 10072 22468 10124
rect 22520 10112 22526 10124
rect 22520 10084 23971 10112
rect 22520 10072 22526 10084
rect 1581 10047 1639 10053
rect 1581 10013 1593 10047
rect 1627 10044 1639 10047
rect 12894 10044 12900 10056
rect 1627 10016 12900 10044
rect 1627 10013 1639 10016
rect 1581 10007 1639 10013
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 12986 10004 12992 10056
rect 13044 10044 13050 10056
rect 20533 10047 20591 10053
rect 13044 10016 20484 10044
rect 13044 10004 13050 10016
rect 1854 9976 1860 9988
rect 1815 9948 1860 9976
rect 1854 9936 1860 9948
rect 1912 9936 1918 9988
rect 12805 9979 12863 9985
rect 12805 9945 12817 9979
rect 12851 9976 12863 9979
rect 13998 9976 14004 9988
rect 12851 9948 14004 9976
rect 12851 9945 12863 9948
rect 12805 9939 12863 9945
rect 13998 9936 14004 9948
rect 14056 9976 14062 9988
rect 14277 9979 14335 9985
rect 14277 9976 14289 9979
rect 14056 9948 14289 9976
rect 14056 9936 14062 9948
rect 14277 9945 14289 9948
rect 14323 9945 14335 9979
rect 20456 9976 20484 10016
rect 20533 10013 20545 10047
rect 20579 10044 20591 10047
rect 20622 10044 20628 10056
rect 20579 10016 20628 10044
rect 20579 10013 20591 10016
rect 20533 10007 20591 10013
rect 20622 10004 20628 10016
rect 20680 10004 20686 10056
rect 20800 10047 20858 10053
rect 20800 10013 20812 10047
rect 20846 10044 20858 10047
rect 21266 10044 21272 10056
rect 20846 10016 21272 10044
rect 20846 10013 20858 10016
rect 20800 10007 20858 10013
rect 21266 10004 21272 10016
rect 21324 10004 21330 10056
rect 21634 10004 21640 10056
rect 21692 10044 21698 10056
rect 21692 10016 21864 10044
rect 21692 10004 21698 10016
rect 21726 9976 21732 9988
rect 20456 9948 21732 9976
rect 14277 9939 14335 9945
rect 21726 9936 21732 9948
rect 21784 9936 21790 9988
rect 21836 9976 21864 10016
rect 22094 10004 22100 10056
rect 22152 10044 22158 10056
rect 23658 10044 23664 10056
rect 22152 10016 23664 10044
rect 22152 10004 22158 10016
rect 23658 10004 23664 10016
rect 23716 10004 23722 10056
rect 23750 10004 23756 10056
rect 23808 10044 23814 10056
rect 23943 10044 23971 10084
rect 24210 10044 24216 10056
rect 23808 10016 23853 10044
rect 23943 10016 24216 10044
rect 23808 10004 23814 10016
rect 24210 10004 24216 10016
rect 24268 10044 24274 10056
rect 24581 10047 24639 10053
rect 24268 10038 24532 10044
rect 24581 10038 24593 10047
rect 24268 10016 24593 10038
rect 24268 10004 24274 10016
rect 24504 10013 24593 10016
rect 24627 10013 24639 10047
rect 24504 10010 24639 10013
rect 24581 10007 24639 10010
rect 25866 10004 25872 10056
rect 25924 10044 25930 10056
rect 27614 10044 27620 10056
rect 25924 10016 27620 10044
rect 25924 10004 25930 10016
rect 27614 10004 27620 10016
rect 27672 10004 27678 10056
rect 27709 10047 27767 10053
rect 27709 10013 27721 10047
rect 27755 10044 27767 10047
rect 29104 10044 29132 10220
rect 30466 10208 30472 10220
rect 30524 10208 30530 10260
rect 31662 10208 31668 10260
rect 31720 10248 31726 10260
rect 31720 10220 36308 10248
rect 31720 10208 31726 10220
rect 29178 10140 29184 10192
rect 29236 10180 29242 10192
rect 30742 10180 30748 10192
rect 29236 10152 29960 10180
rect 29236 10140 29242 10152
rect 27755 10016 29132 10044
rect 27755 10013 27767 10016
rect 27709 10007 27767 10013
rect 29730 10004 29736 10056
rect 29788 10044 29794 10056
rect 29932 10053 29960 10152
rect 30392 10152 30748 10180
rect 30392 10112 30420 10152
rect 30742 10140 30748 10152
rect 30800 10140 30806 10192
rect 30116 10084 30420 10112
rect 30116 10053 30144 10084
rect 30466 10072 30472 10124
rect 30524 10112 30530 10124
rect 30926 10112 30932 10124
rect 30524 10084 30932 10112
rect 30524 10072 30530 10084
rect 30926 10072 30932 10084
rect 30984 10072 30990 10124
rect 31662 10112 31668 10124
rect 31036 10084 31668 10112
rect 29917 10047 29975 10053
rect 29788 10016 29833 10044
rect 29788 10004 29794 10016
rect 29917 10013 29929 10047
rect 29963 10013 29975 10047
rect 29917 10007 29975 10013
rect 30009 10047 30067 10053
rect 30009 10013 30021 10047
rect 30055 10013 30067 10047
rect 30009 10007 30067 10013
rect 30101 10047 30159 10053
rect 30101 10013 30113 10047
rect 30147 10013 30159 10047
rect 30285 10047 30343 10053
rect 30285 10044 30297 10047
rect 30101 10007 30159 10013
rect 30208 10016 30297 10044
rect 21836 9948 26556 9976
rect 14737 9911 14795 9917
rect 14737 9877 14749 9911
rect 14783 9908 14795 9911
rect 26418 9908 26424 9920
rect 14783 9880 26424 9908
rect 14783 9877 14795 9880
rect 14737 9871 14795 9877
rect 26418 9868 26424 9880
rect 26476 9868 26482 9920
rect 26528 9908 26556 9948
rect 26602 9936 26608 9988
rect 26660 9976 26666 9988
rect 27954 9979 28012 9985
rect 27954 9976 27966 9979
rect 26660 9948 27966 9976
rect 26660 9936 26666 9948
rect 27954 9945 27966 9948
rect 28000 9945 28012 9979
rect 27954 9939 28012 9945
rect 29638 9936 29644 9988
rect 29696 9976 29702 9988
rect 30024 9976 30052 10007
rect 29696 9948 30052 9976
rect 29696 9936 29702 9948
rect 28534 9908 28540 9920
rect 26528 9880 28540 9908
rect 28534 9868 28540 9880
rect 28592 9868 28598 9920
rect 29086 9908 29092 9920
rect 29047 9880 29092 9908
rect 29086 9868 29092 9880
rect 29144 9868 29150 9920
rect 29454 9868 29460 9920
rect 29512 9908 29518 9920
rect 30208 9908 30236 10016
rect 30285 10013 30297 10016
rect 30331 10013 30343 10047
rect 30285 10007 30343 10013
rect 30374 10004 30380 10056
rect 30432 10044 30438 10056
rect 31036 10044 31064 10084
rect 31662 10072 31668 10084
rect 31720 10072 31726 10124
rect 36280 10112 36308 10220
rect 37734 10208 37740 10260
rect 37792 10248 37798 10260
rect 37829 10251 37887 10257
rect 37829 10248 37841 10251
rect 37792 10220 37841 10248
rect 37792 10208 37798 10220
rect 37829 10217 37841 10220
rect 37875 10217 37887 10251
rect 37829 10211 37887 10217
rect 38838 10180 38844 10192
rect 38304 10152 38844 10180
rect 38304 10121 38332 10152
rect 38838 10140 38844 10152
rect 38896 10140 38902 10192
rect 57241 10183 57299 10189
rect 57241 10180 57253 10183
rect 41386 10152 57253 10180
rect 38289 10115 38347 10121
rect 38289 10112 38301 10115
rect 36280 10084 38301 10112
rect 38289 10081 38301 10084
rect 38335 10081 38347 10115
rect 38289 10075 38347 10081
rect 38378 10072 38384 10124
rect 38436 10112 38442 10124
rect 41386 10112 41414 10152
rect 57241 10149 57253 10152
rect 57287 10149 57299 10183
rect 57241 10143 57299 10149
rect 58158 10112 58164 10124
rect 38436 10084 38481 10112
rect 38764 10084 41414 10112
rect 58119 10084 58164 10112
rect 38436 10072 38442 10084
rect 31202 10044 31208 10056
rect 30432 10016 31064 10044
rect 31163 10016 31208 10044
rect 30432 10004 30438 10016
rect 31202 10004 31208 10016
rect 31260 10004 31266 10056
rect 35894 10004 35900 10056
rect 35952 10044 35958 10056
rect 36354 10044 36360 10056
rect 35952 10016 36360 10044
rect 35952 10004 35958 10016
rect 36354 10004 36360 10016
rect 36412 10004 36418 10056
rect 38197 10047 38255 10053
rect 38197 10013 38209 10047
rect 38243 10044 38255 10047
rect 38654 10044 38660 10056
rect 38243 10016 38660 10044
rect 38243 10013 38255 10016
rect 38197 10007 38255 10013
rect 38654 10004 38660 10016
rect 38712 10004 38718 10056
rect 34882 9936 34888 9988
rect 34940 9976 34946 9988
rect 38764 9976 38792 10084
rect 58158 10072 58164 10084
rect 58216 10072 58222 10124
rect 40221 10047 40279 10053
rect 40221 10013 40233 10047
rect 40267 10044 40279 10047
rect 42150 10044 42156 10056
rect 40267 10016 42156 10044
rect 40267 10013 40279 10016
rect 40221 10007 40279 10013
rect 42150 10004 42156 10016
rect 42208 10004 42214 10056
rect 53834 10004 53840 10056
rect 53892 10044 53898 10056
rect 57885 10047 57943 10053
rect 57885 10044 57897 10047
rect 53892 10016 57897 10044
rect 53892 10004 53898 10016
rect 57885 10013 57897 10016
rect 57931 10013 57943 10047
rect 57885 10007 57943 10013
rect 34940 9948 38792 9976
rect 34940 9936 34946 9948
rect 39942 9936 39948 9988
rect 40000 9976 40006 9988
rect 40497 9979 40555 9985
rect 40497 9976 40509 9979
rect 40000 9948 40509 9976
rect 40000 9936 40006 9948
rect 40497 9945 40509 9948
rect 40543 9945 40555 9979
rect 45094 9976 45100 9988
rect 40497 9939 40555 9945
rect 41386 9948 45100 9976
rect 29512 9880 30236 9908
rect 30469 9911 30527 9917
rect 29512 9868 29518 9880
rect 30469 9877 30481 9911
rect 30515 9908 30527 9911
rect 31294 9908 31300 9920
rect 30515 9880 31300 9908
rect 30515 9877 30527 9880
rect 30469 9871 30527 9877
rect 31294 9868 31300 9880
rect 31352 9868 31358 9920
rect 32030 9868 32036 9920
rect 32088 9908 32094 9920
rect 32309 9911 32367 9917
rect 32309 9908 32321 9911
rect 32088 9880 32321 9908
rect 32088 9868 32094 9880
rect 32309 9877 32321 9880
rect 32355 9877 32367 9911
rect 32309 9871 32367 9877
rect 32950 9868 32956 9920
rect 33008 9908 33014 9920
rect 41386 9908 41414 9948
rect 45094 9936 45100 9948
rect 45152 9936 45158 9988
rect 57054 9976 57060 9988
rect 57015 9948 57060 9976
rect 57054 9936 57060 9948
rect 57112 9936 57118 9988
rect 33008 9880 41414 9908
rect 33008 9868 33014 9880
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 23566 9704 23572 9716
rect 10560 9676 23572 9704
rect 10560 9664 10566 9676
rect 23566 9664 23572 9676
rect 23624 9664 23630 9716
rect 23658 9664 23664 9716
rect 23716 9704 23722 9716
rect 23716 9676 25728 9704
rect 23716 9664 23722 9676
rect 12437 9639 12495 9645
rect 12437 9605 12449 9639
rect 12483 9636 12495 9639
rect 13998 9636 14004 9648
rect 12483 9608 14004 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 1581 9571 1639 9577
rect 1581 9537 1593 9571
rect 1627 9568 1639 9571
rect 1627 9540 2774 9568
rect 1627 9537 1639 9540
rect 1581 9531 1639 9537
rect 1762 9500 1768 9512
rect 1723 9472 1768 9500
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 2746 9432 2774 9540
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 12544 9500 12572 9608
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 25700 9636 25728 9676
rect 25774 9664 25780 9716
rect 25832 9704 25838 9716
rect 27157 9707 27215 9713
rect 25832 9676 27108 9704
rect 25832 9664 25838 9676
rect 25866 9636 25872 9648
rect 25700 9608 25872 9636
rect 25866 9596 25872 9608
rect 25924 9596 25930 9648
rect 27080 9636 27108 9676
rect 27157 9673 27169 9707
rect 27203 9704 27215 9707
rect 27430 9704 27436 9716
rect 27203 9676 27436 9704
rect 27203 9673 27215 9676
rect 27157 9667 27215 9673
rect 27430 9664 27436 9676
rect 27488 9664 27494 9716
rect 30374 9704 30380 9716
rect 27540 9676 30380 9704
rect 27540 9636 27568 9676
rect 30374 9664 30380 9676
rect 30432 9664 30438 9716
rect 30745 9707 30803 9713
rect 30745 9673 30757 9707
rect 30791 9704 30803 9707
rect 31202 9704 31208 9716
rect 30791 9676 31208 9704
rect 30791 9673 30803 9676
rect 30745 9667 30803 9673
rect 31202 9664 31208 9676
rect 31260 9664 31266 9716
rect 31386 9664 31392 9716
rect 31444 9704 31450 9716
rect 44818 9704 44824 9716
rect 31444 9676 44824 9704
rect 31444 9664 31450 9676
rect 44818 9664 44824 9676
rect 44876 9664 44882 9716
rect 29362 9636 29368 9648
rect 27080 9608 27568 9636
rect 27724 9608 29368 9636
rect 19797 9571 19855 9577
rect 19797 9537 19809 9571
rect 19843 9568 19855 9571
rect 25682 9568 25688 9580
rect 19843 9540 25688 9568
rect 19843 9537 19855 9540
rect 19797 9531 19855 9537
rect 25682 9528 25688 9540
rect 25740 9528 25746 9580
rect 27410 9568 27416 9580
rect 27371 9540 27416 9568
rect 27410 9528 27416 9540
rect 27468 9528 27474 9580
rect 27525 9571 27583 9577
rect 27525 9537 27537 9571
rect 27571 9537 27583 9571
rect 27525 9531 27583 9537
rect 27638 9571 27696 9577
rect 27638 9537 27650 9571
rect 27684 9568 27696 9571
rect 27724 9568 27752 9608
rect 29362 9596 29368 9608
rect 29420 9596 29426 9648
rect 29546 9596 29552 9648
rect 29604 9636 29610 9648
rect 29917 9639 29975 9645
rect 29917 9636 29929 9639
rect 29604 9608 29929 9636
rect 29604 9596 29610 9608
rect 29917 9605 29929 9608
rect 29963 9636 29975 9639
rect 30006 9636 30012 9648
rect 29963 9608 30012 9636
rect 29963 9605 29975 9608
rect 29917 9599 29975 9605
rect 30006 9596 30012 9608
rect 30064 9596 30070 9648
rect 33870 9596 33876 9648
rect 33928 9636 33934 9648
rect 34882 9636 34888 9648
rect 33928 9608 34888 9636
rect 33928 9596 33934 9608
rect 34882 9596 34888 9608
rect 34940 9596 34946 9648
rect 57238 9636 57244 9648
rect 36556 9608 57244 9636
rect 27684 9540 27752 9568
rect 27801 9571 27859 9577
rect 27684 9537 27696 9540
rect 27638 9531 27696 9537
rect 27801 9537 27813 9571
rect 27847 9568 27859 9571
rect 27847 9540 27936 9568
rect 27847 9537 27859 9540
rect 27801 9531 27859 9537
rect 12216 9472 12572 9500
rect 12897 9503 12955 9509
rect 12216 9460 12222 9472
rect 12897 9469 12909 9503
rect 12943 9500 12955 9503
rect 13354 9500 13360 9512
rect 12943 9472 13360 9500
rect 12943 9469 12955 9472
rect 12897 9463 12955 9469
rect 13354 9460 13360 9472
rect 13412 9460 13418 9512
rect 14461 9503 14519 9509
rect 14461 9469 14473 9503
rect 14507 9500 14519 9503
rect 15194 9500 15200 9512
rect 14507 9472 15200 9500
rect 14507 9469 14519 9472
rect 14461 9463 14519 9469
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 19889 9503 19947 9509
rect 19889 9500 19901 9503
rect 18196 9472 19901 9500
rect 18196 9460 18202 9472
rect 19889 9469 19901 9472
rect 19935 9469 19947 9503
rect 19889 9463 19947 9469
rect 20073 9503 20131 9509
rect 20073 9469 20085 9503
rect 20119 9500 20131 9503
rect 20622 9500 20628 9512
rect 20119 9472 20628 9500
rect 20119 9469 20131 9472
rect 20073 9463 20131 9469
rect 12526 9432 12532 9444
rect 2746 9404 12532 9432
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 12710 9432 12716 9444
rect 12671 9404 12716 9432
rect 12710 9392 12716 9404
rect 12768 9392 12774 9444
rect 12986 9392 12992 9444
rect 13044 9432 13050 9444
rect 14277 9435 14335 9441
rect 14277 9432 14289 9435
rect 13044 9404 14289 9432
rect 13044 9392 13050 9404
rect 14277 9401 14289 9404
rect 14323 9401 14335 9435
rect 14277 9395 14335 9401
rect 15746 9392 15752 9444
rect 15804 9432 15810 9444
rect 19904 9432 19932 9463
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 27062 9460 27068 9512
rect 27120 9500 27126 9512
rect 27540 9500 27568 9531
rect 27120 9472 27660 9500
rect 27120 9460 27126 9472
rect 27632 9444 27660 9472
rect 20806 9432 20812 9444
rect 15804 9404 19840 9432
rect 19904 9404 20812 9432
rect 15804 9392 15810 9404
rect 19426 9364 19432 9376
rect 19387 9336 19432 9364
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 19812 9364 19840 9404
rect 20806 9392 20812 9404
rect 20864 9392 20870 9444
rect 23106 9392 23112 9444
rect 23164 9432 23170 9444
rect 26694 9432 26700 9444
rect 23164 9404 26700 9432
rect 23164 9392 23170 9404
rect 26694 9392 26700 9404
rect 26752 9392 26758 9444
rect 27614 9392 27620 9444
rect 27672 9392 27678 9444
rect 27706 9392 27712 9444
rect 27764 9432 27770 9444
rect 27908 9432 27936 9540
rect 28166 9528 28172 9580
rect 28224 9568 28230 9580
rect 28261 9571 28319 9577
rect 28261 9568 28273 9571
rect 28224 9540 28273 9568
rect 28224 9528 28230 9540
rect 28261 9537 28273 9540
rect 28307 9537 28319 9571
rect 28261 9531 28319 9537
rect 28353 9571 28411 9577
rect 28353 9537 28365 9571
rect 28399 9568 28411 9571
rect 29454 9568 29460 9580
rect 28399 9540 29460 9568
rect 28399 9537 28411 9540
rect 28353 9531 28411 9537
rect 29454 9528 29460 9540
rect 29512 9528 29518 9580
rect 30098 9568 30104 9580
rect 30059 9540 30104 9568
rect 30098 9528 30104 9540
rect 30156 9528 30162 9580
rect 30190 9528 30196 9580
rect 30248 9568 30254 9580
rect 30975 9574 31033 9577
rect 30852 9571 31033 9574
rect 30852 9568 30987 9571
rect 30248 9546 30987 9568
rect 30248 9540 30880 9546
rect 30248 9528 30254 9540
rect 30975 9537 30987 9546
rect 31021 9537 31033 9571
rect 31110 9568 31116 9580
rect 31071 9540 31116 9568
rect 30975 9531 31033 9537
rect 31110 9528 31116 9540
rect 31168 9528 31174 9580
rect 31202 9534 31208 9586
rect 31260 9574 31266 9586
rect 31260 9546 31305 9574
rect 31389 9571 31447 9577
rect 31260 9534 31266 9546
rect 31389 9537 31401 9571
rect 31435 9568 31447 9571
rect 31478 9568 31484 9580
rect 31435 9540 31484 9568
rect 31435 9537 31447 9540
rect 31389 9531 31447 9537
rect 31478 9528 31484 9540
rect 31536 9528 31542 9580
rect 34330 9528 34336 9580
rect 34388 9568 34394 9580
rect 34977 9571 35035 9577
rect 34977 9568 34989 9571
rect 34388 9540 34989 9568
rect 34388 9528 34394 9540
rect 34977 9537 34989 9540
rect 35023 9537 35035 9571
rect 34977 9531 35035 9537
rect 35066 9528 35072 9580
rect 35124 9568 35130 9580
rect 35253 9571 35311 9577
rect 35124 9540 35169 9568
rect 35124 9528 35130 9540
rect 35253 9537 35265 9571
rect 35299 9568 35311 9571
rect 35710 9568 35716 9580
rect 35299 9540 35716 9568
rect 35299 9537 35311 9540
rect 35253 9531 35311 9537
rect 35710 9528 35716 9540
rect 35768 9528 35774 9580
rect 30282 9500 30288 9512
rect 30243 9472 30288 9500
rect 30282 9460 30288 9472
rect 30340 9460 30346 9512
rect 31125 9500 31153 9528
rect 34514 9500 34520 9512
rect 31125 9472 34520 9500
rect 34514 9460 34520 9472
rect 34572 9460 34578 9512
rect 35437 9503 35495 9509
rect 35437 9469 35449 9503
rect 35483 9469 35495 9503
rect 35437 9463 35495 9469
rect 27764 9404 27936 9432
rect 27764 9392 27770 9404
rect 30098 9392 30104 9444
rect 30156 9432 30162 9444
rect 32030 9432 32036 9444
rect 30156 9404 32036 9432
rect 30156 9392 30162 9404
rect 32030 9392 32036 9404
rect 32088 9392 32094 9444
rect 32582 9392 32588 9444
rect 32640 9432 32646 9444
rect 35452 9432 35480 9463
rect 32640 9404 35480 9432
rect 32640 9392 32646 9404
rect 28074 9364 28080 9376
rect 19812 9336 28080 9364
rect 28074 9324 28080 9336
rect 28132 9324 28138 9376
rect 28166 9324 28172 9376
rect 28224 9364 28230 9376
rect 29546 9364 29552 9376
rect 28224 9336 29552 9364
rect 28224 9324 28230 9336
rect 29546 9324 29552 9336
rect 29604 9364 29610 9376
rect 36556 9364 36584 9608
rect 57238 9596 57244 9608
rect 57296 9596 57302 9648
rect 57422 9636 57428 9648
rect 57348 9608 57428 9636
rect 37550 9528 37556 9580
rect 37608 9568 37614 9580
rect 37921 9571 37979 9577
rect 37921 9568 37933 9571
rect 37608 9540 37933 9568
rect 37608 9528 37614 9540
rect 37921 9537 37933 9540
rect 37967 9537 37979 9571
rect 37921 9531 37979 9537
rect 38105 9571 38163 9577
rect 38105 9537 38117 9571
rect 38151 9537 38163 9571
rect 38105 9531 38163 9537
rect 37642 9460 37648 9512
rect 37700 9500 37706 9512
rect 38120 9500 38148 9531
rect 38286 9528 38292 9580
rect 38344 9568 38350 9580
rect 38654 9568 38660 9580
rect 38344 9540 38660 9568
rect 38344 9528 38350 9540
rect 38654 9528 38660 9540
rect 38712 9568 38718 9580
rect 39577 9571 39635 9577
rect 39577 9568 39589 9571
rect 38712 9540 39589 9568
rect 38712 9528 38718 9540
rect 39577 9537 39589 9540
rect 39623 9568 39635 9571
rect 39942 9568 39948 9580
rect 39623 9540 39948 9568
rect 39623 9537 39635 9540
rect 39577 9531 39635 9537
rect 39942 9528 39948 9540
rect 40000 9528 40006 9580
rect 40494 9568 40500 9580
rect 40455 9540 40500 9568
rect 40494 9528 40500 9540
rect 40552 9528 40558 9580
rect 40764 9571 40822 9577
rect 40764 9537 40776 9571
rect 40810 9568 40822 9571
rect 41046 9568 41052 9580
rect 40810 9540 41052 9568
rect 40810 9537 40822 9540
rect 40764 9531 40822 9537
rect 41046 9528 41052 9540
rect 41104 9528 41110 9580
rect 56318 9568 56324 9580
rect 45526 9540 56324 9568
rect 37700 9472 38148 9500
rect 37700 9460 37706 9472
rect 39666 9460 39672 9512
rect 39724 9500 39730 9512
rect 39853 9503 39911 9509
rect 39853 9500 39865 9503
rect 39724 9472 39865 9500
rect 39724 9460 39730 9472
rect 39853 9469 39865 9472
rect 39899 9500 39911 9503
rect 40126 9500 40132 9512
rect 39899 9472 40132 9500
rect 39899 9469 39911 9472
rect 39853 9463 39911 9469
rect 40126 9460 40132 9472
rect 40184 9460 40190 9512
rect 40310 9460 40316 9512
rect 40368 9460 40374 9512
rect 36630 9392 36636 9444
rect 36688 9432 36694 9444
rect 39942 9432 39948 9444
rect 36688 9404 39948 9432
rect 36688 9392 36694 9404
rect 39942 9392 39948 9404
rect 40000 9392 40006 9444
rect 40328 9432 40356 9460
rect 40494 9432 40500 9444
rect 40328 9404 40500 9432
rect 40494 9392 40500 9404
rect 40552 9392 40558 9444
rect 41598 9392 41604 9444
rect 41656 9432 41662 9444
rect 45526 9432 45554 9540
rect 56318 9528 56324 9540
rect 56376 9528 56382 9580
rect 57348 9577 57376 9608
rect 57422 9596 57428 9608
rect 57480 9636 57486 9648
rect 57882 9636 57888 9648
rect 57480 9608 57888 9636
rect 57480 9596 57486 9608
rect 57882 9596 57888 9608
rect 57940 9596 57946 9648
rect 57333 9571 57391 9577
rect 57333 9537 57345 9571
rect 57379 9537 57391 9571
rect 57514 9568 57520 9580
rect 57475 9540 57520 9568
rect 57333 9531 57391 9537
rect 57514 9528 57520 9540
rect 57572 9528 57578 9580
rect 50062 9460 50068 9512
rect 50120 9500 50126 9512
rect 50798 9500 50804 9512
rect 50120 9472 50804 9500
rect 50120 9460 50126 9472
rect 50798 9460 50804 9472
rect 50856 9460 50862 9512
rect 41656 9404 45554 9432
rect 41656 9392 41662 9404
rect 29604 9336 36584 9364
rect 29604 9324 29610 9336
rect 37274 9324 37280 9376
rect 37332 9364 37338 9376
rect 37826 9364 37832 9376
rect 37332 9336 37832 9364
rect 37332 9324 37338 9336
rect 37826 9324 37832 9336
rect 37884 9324 37890 9376
rect 38010 9364 38016 9376
rect 37971 9336 38016 9364
rect 38010 9324 38016 9336
rect 38068 9324 38074 9376
rect 40310 9324 40316 9376
rect 40368 9364 40374 9376
rect 41877 9367 41935 9373
rect 41877 9364 41889 9367
rect 40368 9336 41889 9364
rect 40368 9324 40374 9336
rect 41877 9333 41889 9336
rect 41923 9364 41935 9367
rect 53834 9364 53840 9376
rect 41923 9336 53840 9364
rect 41923 9333 41935 9336
rect 41877 9327 41935 9333
rect 53834 9324 53840 9336
rect 53892 9324 53898 9376
rect 57425 9367 57483 9373
rect 57425 9333 57437 9367
rect 57471 9364 57483 9367
rect 58250 9364 58256 9376
rect 57471 9336 58256 9364
rect 57471 9333 57483 9336
rect 57425 9327 57483 9333
rect 58250 9324 58256 9336
rect 58308 9324 58314 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 18230 9120 18236 9172
rect 18288 9160 18294 9172
rect 20806 9160 20812 9172
rect 18288 9132 20668 9160
rect 20767 9132 20812 9160
rect 18288 9120 18294 9132
rect 19426 9052 19432 9104
rect 19484 9052 19490 9104
rect 20640 9092 20668 9132
rect 20806 9120 20812 9132
rect 20864 9120 20870 9172
rect 27798 9160 27804 9172
rect 22066 9132 27804 9160
rect 22066 9092 22094 9132
rect 27798 9120 27804 9132
rect 27856 9120 27862 9172
rect 28074 9120 28080 9172
rect 28132 9160 28138 9172
rect 30374 9160 30380 9172
rect 28132 9132 30380 9160
rect 28132 9120 28138 9132
rect 30374 9120 30380 9132
rect 30432 9120 30438 9172
rect 30466 9120 30472 9172
rect 30524 9160 30530 9172
rect 31662 9160 31668 9172
rect 30524 9132 31668 9160
rect 30524 9120 30530 9132
rect 31662 9120 31668 9132
rect 31720 9160 31726 9172
rect 31846 9160 31852 9172
rect 31720 9132 31852 9160
rect 31720 9120 31726 9132
rect 31846 9120 31852 9132
rect 31904 9160 31910 9172
rect 37274 9160 37280 9172
rect 31904 9132 37280 9160
rect 31904 9120 31910 9132
rect 37274 9120 37280 9132
rect 37332 9120 37338 9172
rect 37369 9163 37427 9169
rect 37369 9129 37381 9163
rect 37415 9160 37427 9163
rect 37458 9160 37464 9172
rect 37415 9132 37464 9160
rect 37415 9129 37427 9132
rect 37369 9123 37427 9129
rect 37458 9120 37464 9132
rect 37516 9120 37522 9172
rect 37826 9120 37832 9172
rect 37884 9160 37890 9172
rect 38102 9160 38108 9172
rect 37884 9132 38108 9160
rect 37884 9120 37890 9132
rect 38102 9120 38108 9132
rect 38160 9120 38166 9172
rect 38286 9120 38292 9172
rect 38344 9160 38350 9172
rect 39025 9163 39083 9169
rect 39025 9160 39037 9163
rect 38344 9132 39037 9160
rect 38344 9120 38350 9132
rect 39025 9129 39037 9132
rect 39071 9160 39083 9163
rect 39758 9160 39764 9172
rect 39071 9132 39764 9160
rect 39071 9129 39083 9132
rect 39025 9123 39083 9129
rect 39758 9120 39764 9132
rect 39816 9120 39822 9172
rect 39942 9120 39948 9172
rect 40000 9160 40006 9172
rect 40000 9132 40908 9160
rect 40000 9120 40006 9132
rect 34606 9092 34612 9104
rect 20640 9064 22094 9092
rect 25608 9064 34612 9092
rect 19444 9024 19472 9052
rect 19444 8996 19564 9024
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8956 1639 8959
rect 11790 8956 11796 8968
rect 1627 8928 11796 8956
rect 1627 8925 1639 8928
rect 1581 8919 1639 8925
rect 11790 8916 11796 8928
rect 11848 8916 11854 8968
rect 19426 8956 19432 8968
rect 19387 8928 19432 8956
rect 19426 8916 19432 8928
rect 19484 8916 19490 8968
rect 19536 8956 19564 8996
rect 23658 8984 23664 9036
rect 23716 9024 23722 9036
rect 23753 9027 23811 9033
rect 23753 9024 23765 9027
rect 23716 8996 23765 9024
rect 23716 8984 23722 8996
rect 23753 8993 23765 8996
rect 23799 8993 23811 9027
rect 24578 9024 24584 9036
rect 24539 8996 24584 9024
rect 23753 8987 23811 8993
rect 24578 8984 24584 8996
rect 24636 8984 24642 9036
rect 19685 8959 19743 8965
rect 19685 8956 19697 8959
rect 19536 8928 19697 8956
rect 19685 8925 19697 8928
rect 19731 8925 19743 8959
rect 23566 8956 23572 8968
rect 23527 8928 23572 8956
rect 19685 8919 19743 8925
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 25608 8956 25636 9064
rect 34606 9052 34612 9064
rect 34664 9092 34670 9104
rect 34977 9095 35035 9101
rect 34977 9092 34989 9095
rect 34664 9064 34989 9092
rect 34664 9052 34670 9064
rect 34977 9061 34989 9064
rect 35023 9061 35035 9095
rect 34977 9055 35035 9061
rect 35360 9064 36400 9092
rect 30653 9027 30711 9033
rect 30653 8993 30665 9027
rect 30699 9024 30711 9027
rect 35360 9024 35388 9064
rect 36262 9024 36268 9036
rect 30699 8996 35388 9024
rect 35452 8996 36268 9024
rect 30699 8993 30711 8996
rect 30653 8987 30711 8993
rect 23768 8928 25636 8956
rect 1854 8888 1860 8900
rect 1815 8860 1860 8888
rect 1854 8848 1860 8860
rect 1912 8848 1918 8900
rect 16482 8848 16488 8900
rect 16540 8888 16546 8900
rect 23768 8888 23796 8928
rect 30466 8916 30472 8968
rect 30524 8956 30530 8968
rect 30837 8959 30895 8965
rect 30837 8956 30849 8959
rect 30524 8928 30849 8956
rect 30524 8916 30530 8928
rect 30837 8925 30849 8928
rect 30883 8925 30895 8959
rect 30837 8919 30895 8925
rect 30929 8959 30987 8965
rect 30929 8925 30941 8959
rect 30975 8925 30987 8959
rect 30929 8919 30987 8925
rect 31113 8959 31171 8965
rect 31113 8925 31125 8959
rect 31159 8925 31171 8959
rect 31113 8919 31171 8925
rect 31205 8959 31263 8965
rect 31205 8925 31217 8959
rect 31251 8956 31263 8959
rect 31294 8956 31300 8968
rect 31251 8928 31300 8956
rect 31251 8925 31263 8928
rect 31205 8919 31263 8925
rect 16540 8860 23796 8888
rect 24848 8891 24906 8897
rect 16540 8848 16546 8860
rect 24848 8857 24860 8891
rect 24894 8888 24906 8891
rect 25866 8888 25872 8900
rect 24894 8860 25872 8888
rect 24894 8857 24906 8860
rect 24848 8851 24906 8857
rect 25866 8848 25872 8860
rect 25924 8848 25930 8900
rect 29730 8848 29736 8900
rect 29788 8888 29794 8900
rect 30944 8888 30972 8919
rect 29788 8860 30972 8888
rect 31128 8888 31156 8919
rect 31294 8916 31300 8928
rect 31352 8916 31358 8968
rect 31662 8916 31668 8968
rect 31720 8956 31726 8968
rect 31849 8959 31907 8965
rect 31849 8956 31861 8959
rect 31720 8928 31861 8956
rect 31720 8916 31726 8928
rect 31849 8925 31861 8928
rect 31895 8925 31907 8959
rect 32030 8956 32036 8968
rect 31991 8928 32036 8956
rect 31849 8919 31907 8925
rect 31478 8888 31484 8900
rect 31128 8860 31484 8888
rect 29788 8848 29794 8860
rect 31478 8848 31484 8860
rect 31536 8888 31542 8900
rect 31754 8888 31760 8900
rect 31536 8860 31760 8888
rect 31536 8848 31542 8860
rect 31754 8848 31760 8860
rect 31812 8848 31818 8900
rect 31864 8888 31892 8919
rect 32030 8916 32036 8928
rect 32088 8916 32094 8968
rect 32122 8916 32128 8968
rect 32180 8956 32186 8968
rect 32585 8959 32643 8965
rect 32180 8928 32225 8956
rect 32180 8916 32186 8928
rect 32585 8925 32597 8959
rect 32631 8925 32643 8959
rect 32585 8919 32643 8925
rect 32769 8959 32827 8965
rect 32769 8925 32781 8959
rect 32815 8925 32827 8959
rect 32769 8919 32827 8925
rect 32398 8888 32404 8900
rect 31864 8860 32404 8888
rect 32398 8848 32404 8860
rect 32456 8848 32462 8900
rect 17954 8780 17960 8832
rect 18012 8820 18018 8832
rect 19978 8820 19984 8832
rect 18012 8792 19984 8820
rect 18012 8780 18018 8792
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 25958 8820 25964 8832
rect 25919 8792 25964 8820
rect 25958 8780 25964 8792
rect 26016 8780 26022 8832
rect 31202 8780 31208 8832
rect 31260 8820 31266 8832
rect 31665 8823 31723 8829
rect 31665 8820 31677 8823
rect 31260 8792 31677 8820
rect 31260 8780 31266 8792
rect 31665 8789 31677 8792
rect 31711 8789 31723 8823
rect 31665 8783 31723 8789
rect 31938 8780 31944 8832
rect 31996 8820 32002 8832
rect 32600 8820 32628 8919
rect 32784 8888 32812 8919
rect 34790 8916 34796 8968
rect 34848 8956 34854 8968
rect 35452 8965 35480 8996
rect 36262 8984 36268 8996
rect 36320 8984 36326 9036
rect 36372 9024 36400 9064
rect 36446 9052 36452 9104
rect 36504 9092 36510 9104
rect 39390 9092 39396 9104
rect 36504 9064 39396 9092
rect 36504 9052 36510 9064
rect 39390 9052 39396 9064
rect 39448 9052 39454 9104
rect 40126 9052 40132 9104
rect 40184 9092 40190 9104
rect 40880 9092 40908 9132
rect 41046 9120 41052 9172
rect 41104 9160 41110 9172
rect 41417 9163 41475 9169
rect 41417 9160 41429 9163
rect 41104 9132 41429 9160
rect 41104 9120 41110 9132
rect 41417 9129 41429 9132
rect 41463 9129 41475 9163
rect 58342 9160 58348 9172
rect 41417 9123 41475 9129
rect 45526 9132 58348 9160
rect 45526 9092 45554 9132
rect 58342 9120 58348 9132
rect 58400 9120 58406 9172
rect 40184 9064 40807 9092
rect 40880 9064 45554 9092
rect 40184 9052 40190 9064
rect 40779 9024 40807 9064
rect 41046 9024 41052 9036
rect 36372 8996 40724 9024
rect 40779 8996 41052 9024
rect 35161 8959 35219 8965
rect 35161 8956 35173 8959
rect 34848 8928 35173 8956
rect 34848 8916 34854 8928
rect 35161 8925 35173 8928
rect 35207 8925 35219 8959
rect 35161 8919 35219 8925
rect 35253 8959 35311 8965
rect 35253 8925 35265 8959
rect 35299 8925 35311 8959
rect 35253 8919 35311 8925
rect 35437 8959 35495 8965
rect 35437 8925 35449 8959
rect 35483 8925 35495 8959
rect 35437 8919 35495 8925
rect 32858 8888 32864 8900
rect 32784 8860 32864 8888
rect 32858 8848 32864 8860
rect 32916 8888 32922 8900
rect 34882 8888 34888 8900
rect 32916 8860 34888 8888
rect 32916 8848 32922 8860
rect 34882 8848 34888 8860
rect 34940 8848 34946 8900
rect 35268 8888 35296 8919
rect 35526 8916 35532 8968
rect 35584 8956 35590 8968
rect 37274 8956 37280 8968
rect 35584 8928 35629 8956
rect 37235 8928 37280 8956
rect 35584 8916 35590 8928
rect 37274 8916 37280 8928
rect 37332 8916 37338 8968
rect 37737 8959 37795 8965
rect 37737 8925 37749 8959
rect 37783 8956 37795 8959
rect 38562 8956 38568 8968
rect 37783 8928 38568 8956
rect 37783 8925 37795 8928
rect 37737 8919 37795 8925
rect 38562 8916 38568 8928
rect 38620 8916 38626 8968
rect 38746 8916 38752 8968
rect 38804 8956 38810 8968
rect 40037 8959 40095 8965
rect 40037 8956 40049 8959
rect 38804 8928 40049 8956
rect 38804 8916 38810 8928
rect 40037 8925 40049 8928
rect 40083 8925 40095 8959
rect 40310 8956 40316 8968
rect 40271 8928 40316 8956
rect 40037 8919 40095 8925
rect 40310 8916 40316 8928
rect 40368 8916 40374 8968
rect 40405 8959 40463 8965
rect 40405 8925 40417 8959
rect 40451 8956 40463 8959
rect 40494 8956 40500 8968
rect 40451 8928 40500 8956
rect 40451 8925 40463 8928
rect 40405 8919 40463 8925
rect 40494 8916 40500 8928
rect 40552 8916 40558 8968
rect 40696 8956 40724 8996
rect 41046 8984 41052 8996
rect 41104 8984 41110 9036
rect 43346 9024 43352 9036
rect 41156 8996 43352 9024
rect 41156 8956 41184 8996
rect 43346 8984 43352 8996
rect 43404 8984 43410 9036
rect 56870 9024 56876 9036
rect 56831 8996 56876 9024
rect 56870 8984 56876 8996
rect 56928 8984 56934 9036
rect 40696 8928 41184 8956
rect 41233 8959 41291 8965
rect 41233 8925 41245 8959
rect 41279 8925 41291 8959
rect 50062 8956 50068 8968
rect 41233 8919 41291 8925
rect 41340 8928 50068 8956
rect 37090 8888 37096 8900
rect 35268 8860 37096 8888
rect 37090 8848 37096 8860
rect 37148 8848 37154 8900
rect 38013 8891 38071 8897
rect 38013 8857 38025 8891
rect 38059 8888 38071 8891
rect 38102 8888 38108 8900
rect 38059 8860 38108 8888
rect 38059 8857 38071 8860
rect 38013 8851 38071 8857
rect 38102 8848 38108 8860
rect 38160 8848 38166 8900
rect 38194 8848 38200 8900
rect 38252 8888 38258 8900
rect 38473 8891 38531 8897
rect 38473 8888 38485 8891
rect 38252 8860 38485 8888
rect 38252 8848 38258 8860
rect 38473 8857 38485 8860
rect 38519 8888 38531 8891
rect 38841 8891 38899 8897
rect 38841 8888 38853 8891
rect 38519 8860 38853 8888
rect 38519 8857 38531 8860
rect 38473 8851 38531 8857
rect 38841 8857 38853 8860
rect 38887 8888 38899 8891
rect 40218 8888 40224 8900
rect 38887 8860 40080 8888
rect 40179 8860 40224 8888
rect 38887 8857 38899 8860
rect 38841 8851 38899 8857
rect 31996 8792 32628 8820
rect 32677 8823 32735 8829
rect 31996 8780 32002 8792
rect 32677 8789 32689 8823
rect 32723 8820 32735 8823
rect 34422 8820 34428 8832
rect 32723 8792 34428 8820
rect 32723 8789 32735 8792
rect 32677 8783 32735 8789
rect 34422 8780 34428 8792
rect 34480 8780 34486 8832
rect 37826 8780 37832 8832
rect 37884 8820 37890 8832
rect 38746 8820 38752 8832
rect 37884 8792 38752 8820
rect 37884 8780 37890 8792
rect 38746 8780 38752 8792
rect 38804 8780 38810 8832
rect 39022 8780 39028 8832
rect 39080 8829 39086 8832
rect 39080 8823 39099 8829
rect 39087 8789 39099 8823
rect 39206 8820 39212 8832
rect 39167 8792 39212 8820
rect 39080 8783 39099 8789
rect 39080 8780 39086 8783
rect 39206 8780 39212 8792
rect 39264 8780 39270 8832
rect 40052 8820 40080 8860
rect 40218 8848 40224 8860
rect 40276 8848 40282 8900
rect 41248 8888 41276 8919
rect 40604 8860 41276 8888
rect 40310 8820 40316 8832
rect 40052 8792 40316 8820
rect 40310 8780 40316 8792
rect 40368 8780 40374 8832
rect 40604 8829 40632 8860
rect 40589 8823 40647 8829
rect 40589 8789 40601 8823
rect 40635 8789 40647 8823
rect 40589 8783 40647 8789
rect 41046 8780 41052 8832
rect 41104 8820 41110 8832
rect 41340 8820 41368 8928
rect 50062 8916 50068 8928
rect 50120 8916 50126 8968
rect 57140 8891 57198 8897
rect 57140 8857 57152 8891
rect 57186 8888 57198 8891
rect 58066 8888 58072 8900
rect 57186 8860 58072 8888
rect 57186 8857 57198 8860
rect 57140 8851 57198 8857
rect 58066 8848 58072 8860
rect 58124 8848 58130 8900
rect 41104 8792 41368 8820
rect 41104 8780 41110 8792
rect 43346 8780 43352 8832
rect 43404 8820 43410 8832
rect 56594 8820 56600 8832
rect 43404 8792 56600 8820
rect 43404 8780 43410 8792
rect 56594 8780 56600 8792
rect 56652 8780 56658 8832
rect 57514 8780 57520 8832
rect 57572 8820 57578 8832
rect 58253 8823 58311 8829
rect 58253 8820 58265 8823
rect 57572 8792 58265 8820
rect 57572 8780 57578 8792
rect 58253 8789 58265 8792
rect 58299 8789 58311 8823
rect 58253 8783 58311 8789
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 11790 8616 11796 8628
rect 11751 8588 11796 8616
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 12406 8588 19564 8616
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8480 12127 8483
rect 12406 8480 12434 8588
rect 13078 8548 13084 8560
rect 13004 8520 13084 8548
rect 13004 8489 13032 8520
rect 13078 8508 13084 8520
rect 13136 8508 13142 8560
rect 18233 8551 18291 8557
rect 18233 8517 18245 8551
rect 18279 8548 18291 8551
rect 18322 8548 18328 8560
rect 18279 8520 18328 8548
rect 18279 8517 18291 8520
rect 18233 8511 18291 8517
rect 18322 8508 18328 8520
rect 18380 8508 18386 8560
rect 19426 8548 19432 8560
rect 19076 8520 19432 8548
rect 12115 8452 12434 8480
rect 12989 8483 13047 8489
rect 12115 8449 12127 8452
rect 12069 8443 12127 8449
rect 12989 8449 13001 8483
rect 13035 8449 13047 8483
rect 18138 8480 18144 8492
rect 12989 8443 13047 8449
rect 13096 8452 18144 8480
rect 11974 8412 11980 8424
rect 11935 8384 11980 8412
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12158 8412 12164 8424
rect 12119 8384 12164 8412
rect 12158 8372 12164 8384
rect 12216 8372 12222 8424
rect 12250 8372 12256 8424
rect 12308 8412 12314 8424
rect 12308 8384 12353 8412
rect 12308 8372 12314 8384
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 13096 8421 13124 8452
rect 18138 8440 18144 8452
rect 18196 8440 18202 8492
rect 19076 8489 19104 8520
rect 19426 8508 19432 8520
rect 19484 8508 19490 8560
rect 19536 8548 19564 8588
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 24305 8619 24363 8625
rect 24305 8616 24317 8619
rect 20036 8588 24317 8616
rect 20036 8576 20042 8588
rect 24305 8585 24317 8588
rect 24351 8585 24363 8619
rect 25866 8616 25872 8628
rect 25827 8588 25872 8616
rect 24305 8579 24363 8585
rect 25866 8576 25872 8588
rect 25924 8576 25930 8628
rect 26237 8619 26295 8625
rect 26237 8585 26249 8619
rect 26283 8616 26295 8619
rect 26510 8616 26516 8628
rect 26283 8588 26516 8616
rect 26283 8585 26295 8588
rect 26237 8579 26295 8585
rect 26510 8576 26516 8588
rect 26568 8576 26574 8628
rect 29730 8616 29736 8628
rect 26620 8588 29040 8616
rect 29691 8588 29736 8616
rect 25958 8548 25964 8560
rect 19536 8520 25964 8548
rect 25958 8508 25964 8520
rect 26016 8548 26022 8560
rect 26329 8551 26387 8557
rect 26329 8548 26341 8551
rect 26016 8520 26341 8548
rect 26016 8508 26022 8520
rect 26329 8517 26341 8520
rect 26375 8517 26387 8551
rect 26329 8511 26387 8517
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8449 19119 8483
rect 19317 8483 19375 8489
rect 19317 8480 19329 8483
rect 19061 8443 19119 8449
rect 19168 8452 19329 8480
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12584 8384 12817 8412
rect 12584 8372 12590 8384
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 13081 8415 13139 8421
rect 13081 8381 13093 8415
rect 13127 8381 13139 8415
rect 13081 8375 13139 8381
rect 13173 8415 13231 8421
rect 13173 8381 13185 8415
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 12176 8344 12204 8372
rect 13188 8344 13216 8375
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13320 8384 13365 8412
rect 13320 8372 13326 8384
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18325 8415 18383 8421
rect 18325 8412 18337 8415
rect 18012 8384 18337 8412
rect 18012 8372 18018 8384
rect 18325 8381 18337 8384
rect 18371 8381 18383 8415
rect 18325 8375 18383 8381
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8412 18567 8415
rect 18598 8412 18604 8424
rect 18555 8384 18604 8412
rect 18555 8381 18567 8384
rect 18509 8375 18567 8381
rect 18598 8372 18604 8384
rect 18656 8412 18662 8424
rect 18966 8412 18972 8424
rect 18656 8384 18972 8412
rect 18656 8372 18662 8384
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 19168 8412 19196 8452
rect 19317 8449 19329 8452
rect 19363 8449 19375 8483
rect 19317 8443 19375 8449
rect 23109 8483 23167 8489
rect 23109 8449 23121 8483
rect 23155 8480 23167 8483
rect 24762 8480 24768 8492
rect 23155 8452 24768 8480
rect 23155 8449 23167 8452
rect 23109 8443 23167 8449
rect 24762 8440 24768 8452
rect 24820 8440 24826 8492
rect 26620 8480 26648 8588
rect 29012 8557 29040 8588
rect 29730 8576 29736 8588
rect 29788 8576 29794 8628
rect 30742 8576 30748 8628
rect 30800 8616 30806 8628
rect 31570 8616 31576 8628
rect 30800 8588 31576 8616
rect 30800 8576 30806 8588
rect 31570 8576 31576 8588
rect 31628 8576 31634 8628
rect 34977 8619 35035 8625
rect 34977 8585 34989 8619
rect 35023 8616 35035 8619
rect 40218 8616 40224 8628
rect 35023 8588 40224 8616
rect 35023 8585 35035 8588
rect 34977 8579 35035 8585
rect 40218 8576 40224 8588
rect 40276 8576 40282 8628
rect 56318 8616 56324 8628
rect 56279 8588 56324 8616
rect 56318 8576 56324 8588
rect 56376 8576 56382 8628
rect 57146 8576 57152 8628
rect 57204 8616 57210 8628
rect 58250 8616 58256 8628
rect 57204 8588 58112 8616
rect 58211 8588 58256 8616
rect 57204 8576 57210 8588
rect 27985 8551 28043 8557
rect 27985 8517 27997 8551
rect 28031 8548 28043 8551
rect 28997 8551 29055 8557
rect 28031 8520 28856 8548
rect 28031 8517 28043 8520
rect 27985 8511 28043 8517
rect 26252 8452 26648 8480
rect 19076 8384 19196 8412
rect 13906 8344 13912 8356
rect 12176 8316 13912 8344
rect 13906 8304 13912 8316
rect 13964 8304 13970 8356
rect 17865 8347 17923 8353
rect 17865 8313 17877 8347
rect 17911 8344 17923 8347
rect 19076 8344 19104 8384
rect 20438 8372 20444 8424
rect 20496 8412 20502 8424
rect 20496 8384 20576 8412
rect 20496 8372 20502 8384
rect 17911 8316 19104 8344
rect 17911 8313 17923 8316
rect 17865 8307 17923 8313
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 19058 8276 19064 8288
rect 12032 8248 19064 8276
rect 12032 8236 12038 8248
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 19702 8236 19708 8288
rect 19760 8276 19766 8288
rect 20441 8279 20499 8285
rect 20441 8276 20453 8279
rect 19760 8248 20453 8276
rect 19760 8236 19766 8248
rect 20441 8245 20453 8248
rect 20487 8245 20499 8279
rect 20548 8276 20576 8384
rect 21818 8372 21824 8424
rect 21876 8412 21882 8424
rect 23014 8412 23020 8424
rect 21876 8384 23020 8412
rect 21876 8372 21882 8384
rect 23014 8372 23020 8384
rect 23072 8372 23078 8424
rect 24210 8372 24216 8424
rect 24268 8412 24274 8424
rect 26252 8412 26280 8452
rect 28074 8440 28080 8492
rect 28132 8480 28138 8492
rect 28828 8489 28856 8520
rect 28997 8517 29009 8551
rect 29043 8548 29055 8551
rect 30006 8548 30012 8560
rect 29043 8520 30012 8548
rect 29043 8517 29055 8520
rect 28997 8511 29055 8517
rect 30006 8508 30012 8520
rect 30064 8548 30070 8560
rect 30653 8551 30711 8557
rect 30653 8548 30665 8551
rect 30064 8520 30665 8548
rect 30064 8508 30070 8520
rect 30653 8517 30665 8520
rect 30699 8517 30711 8551
rect 32122 8548 32128 8560
rect 30653 8511 30711 8517
rect 30760 8520 32128 8548
rect 30760 8492 30788 8520
rect 32122 8508 32128 8520
rect 32180 8508 32186 8560
rect 32398 8508 32404 8560
rect 32456 8548 32462 8560
rect 34606 8548 34612 8560
rect 32456 8520 34376 8548
rect 34567 8520 34612 8548
rect 32456 8508 32462 8520
rect 28169 8483 28227 8489
rect 28169 8480 28181 8483
rect 28132 8452 28181 8480
rect 28132 8440 28138 8452
rect 28169 8449 28181 8452
rect 28215 8449 28227 8483
rect 28169 8443 28227 8449
rect 28813 8483 28871 8489
rect 28813 8449 28825 8483
rect 28859 8480 28871 8483
rect 29454 8480 29460 8492
rect 28859 8452 29460 8480
rect 28859 8449 28871 8452
rect 28813 8443 28871 8449
rect 29454 8440 29460 8452
rect 29512 8440 29518 8492
rect 29641 8483 29699 8489
rect 29641 8449 29653 8483
rect 29687 8449 29699 8483
rect 30466 8480 30472 8492
rect 30427 8452 30472 8480
rect 29641 8443 29699 8449
rect 26418 8412 26424 8424
rect 24268 8384 26280 8412
rect 26379 8384 26424 8412
rect 24268 8372 24274 8384
rect 26418 8372 26424 8384
rect 26476 8372 26482 8424
rect 29656 8412 29684 8443
rect 30466 8440 30472 8452
rect 30524 8440 30530 8492
rect 30742 8480 30748 8492
rect 30655 8452 30748 8480
rect 30742 8440 30748 8452
rect 30800 8440 30806 8492
rect 31294 8440 31300 8492
rect 31352 8480 31358 8492
rect 31481 8483 31539 8489
rect 31481 8480 31493 8483
rect 31352 8452 31493 8480
rect 31352 8440 31358 8452
rect 31481 8449 31493 8452
rect 31527 8449 31539 8483
rect 31481 8443 31539 8449
rect 31570 8440 31576 8492
rect 31628 8480 31634 8492
rect 31628 8452 31673 8480
rect 31628 8440 31634 8452
rect 32306 8440 32312 8492
rect 32364 8480 32370 8492
rect 32585 8483 32643 8489
rect 32585 8480 32597 8483
rect 32364 8452 32597 8480
rect 32364 8440 32370 8452
rect 32585 8449 32597 8452
rect 32631 8449 32643 8483
rect 32766 8480 32772 8492
rect 32727 8452 32772 8480
rect 32585 8443 32643 8449
rect 32766 8440 32772 8452
rect 32824 8440 32830 8492
rect 34348 8489 34376 8520
rect 34606 8508 34612 8520
rect 34664 8508 34670 8560
rect 34698 8508 34704 8560
rect 34756 8548 34762 8560
rect 39206 8548 39212 8560
rect 34756 8520 34801 8548
rect 35360 8520 39212 8548
rect 34756 8508 34762 8520
rect 33413 8483 33471 8489
rect 33413 8449 33425 8483
rect 33459 8480 33471 8483
rect 34333 8483 34391 8489
rect 33459 8452 34284 8480
rect 33459 8449 33471 8452
rect 33413 8443 33471 8449
rect 26528 8384 29684 8412
rect 25498 8304 25504 8356
rect 25556 8344 25562 8356
rect 26528 8344 26556 8384
rect 30374 8372 30380 8424
rect 30432 8412 30438 8424
rect 31389 8415 31447 8421
rect 31389 8412 31401 8415
rect 30432 8384 31401 8412
rect 30432 8372 30438 8384
rect 31389 8381 31401 8384
rect 31435 8381 31447 8415
rect 31662 8412 31668 8424
rect 31623 8384 31668 8412
rect 31389 8375 31447 8381
rect 31662 8372 31668 8384
rect 31720 8372 31726 8424
rect 32677 8415 32735 8421
rect 32677 8381 32689 8415
rect 32723 8412 32735 8415
rect 33318 8412 33324 8424
rect 32723 8384 33324 8412
rect 32723 8381 32735 8384
rect 32677 8375 32735 8381
rect 33318 8372 33324 8384
rect 33376 8372 33382 8424
rect 33686 8412 33692 8424
rect 33647 8384 33692 8412
rect 33686 8372 33692 8384
rect 33744 8412 33750 8424
rect 33962 8412 33968 8424
rect 33744 8384 33968 8412
rect 33744 8372 33750 8384
rect 33962 8372 33968 8384
rect 34020 8372 34026 8424
rect 34256 8412 34284 8452
rect 34333 8449 34345 8483
rect 34379 8449 34391 8483
rect 34333 8443 34391 8449
rect 34422 8440 34428 8492
rect 34480 8480 34486 8492
rect 34882 8489 34888 8492
rect 34839 8483 34888 8489
rect 34480 8452 34525 8480
rect 34480 8440 34486 8452
rect 34839 8449 34851 8483
rect 34885 8449 34888 8483
rect 34839 8443 34888 8449
rect 34882 8440 34888 8443
rect 34940 8440 34946 8492
rect 35360 8412 35388 8520
rect 39206 8508 39212 8520
rect 39264 8508 39270 8560
rect 39390 8508 39396 8560
rect 39448 8548 39454 8560
rect 41598 8548 41604 8560
rect 39448 8520 41604 8548
rect 39448 8508 39454 8520
rect 41598 8508 41604 8520
rect 41656 8508 41662 8560
rect 57330 8548 57336 8560
rect 57291 8520 57336 8548
rect 57330 8508 57336 8520
rect 57388 8508 57394 8560
rect 58084 8557 58112 8588
rect 58250 8576 58256 8588
rect 58308 8576 58314 8628
rect 58069 8551 58127 8557
rect 58069 8517 58081 8551
rect 58115 8517 58127 8551
rect 58069 8511 58127 8517
rect 35437 8483 35495 8489
rect 35437 8449 35449 8483
rect 35483 8480 35495 8483
rect 37553 8483 37611 8489
rect 35483 8452 37412 8480
rect 35483 8449 35495 8452
rect 35437 8443 35495 8449
rect 34256 8384 35388 8412
rect 35526 8372 35532 8424
rect 35584 8412 35590 8424
rect 35621 8415 35679 8421
rect 35621 8412 35633 8415
rect 35584 8384 35633 8412
rect 35584 8372 35590 8384
rect 35621 8381 35633 8384
rect 35667 8381 35679 8415
rect 35621 8375 35679 8381
rect 29178 8344 29184 8356
rect 25556 8316 26556 8344
rect 29139 8316 29184 8344
rect 25556 8304 25562 8316
rect 29178 8304 29184 8316
rect 29236 8304 29242 8356
rect 30285 8347 30343 8353
rect 30285 8313 30297 8347
rect 30331 8313 30343 8347
rect 30285 8307 30343 8313
rect 31205 8347 31263 8353
rect 31205 8313 31217 8347
rect 31251 8344 31263 8347
rect 33410 8344 33416 8356
rect 31251 8316 33416 8344
rect 31251 8313 31263 8316
rect 31205 8307 31263 8313
rect 26786 8276 26792 8288
rect 20548 8248 26792 8276
rect 20441 8239 20499 8245
rect 26786 8236 26792 8248
rect 26844 8236 26850 8288
rect 28350 8276 28356 8288
rect 28311 8248 28356 8276
rect 28350 8236 28356 8248
rect 28408 8236 28414 8288
rect 30300 8276 30328 8307
rect 33410 8304 33416 8316
rect 33468 8304 33474 8356
rect 37384 8344 37412 8452
rect 37553 8449 37565 8483
rect 37599 8480 37611 8483
rect 37734 8480 37740 8492
rect 37599 8452 37740 8480
rect 37599 8449 37611 8452
rect 37553 8443 37611 8449
rect 37734 8440 37740 8452
rect 37792 8480 37798 8492
rect 38102 8480 38108 8492
rect 37792 8452 38108 8480
rect 37792 8440 37798 8452
rect 38102 8440 38108 8452
rect 38160 8440 38166 8492
rect 38289 8483 38347 8489
rect 38289 8449 38301 8483
rect 38335 8449 38347 8483
rect 38289 8443 38347 8449
rect 37458 8372 37464 8424
rect 37516 8412 37522 8424
rect 38304 8412 38332 8443
rect 38654 8440 38660 8492
rect 38712 8480 38718 8492
rect 39761 8483 39819 8489
rect 38712 8452 38757 8480
rect 38712 8440 38718 8452
rect 39761 8449 39773 8483
rect 39807 8480 39819 8483
rect 40126 8480 40132 8492
rect 39807 8452 40132 8480
rect 39807 8449 39819 8452
rect 39761 8443 39819 8449
rect 40126 8440 40132 8452
rect 40184 8440 40190 8492
rect 40310 8440 40316 8492
rect 40368 8480 40374 8492
rect 56226 8480 56232 8492
rect 40368 8452 48314 8480
rect 56187 8452 56232 8480
rect 40368 8440 40374 8452
rect 37516 8384 38332 8412
rect 38672 8412 38700 8440
rect 39206 8412 39212 8424
rect 38672 8384 39212 8412
rect 37516 8372 37522 8384
rect 39206 8372 39212 8384
rect 39264 8372 39270 8424
rect 40037 8415 40095 8421
rect 40037 8381 40049 8415
rect 40083 8412 40095 8415
rect 40494 8412 40500 8424
rect 40083 8384 40500 8412
rect 40083 8381 40095 8384
rect 40037 8375 40095 8381
rect 38930 8344 38936 8356
rect 34440 8316 35296 8344
rect 31386 8276 31392 8288
rect 30300 8248 31392 8276
rect 31386 8236 31392 8248
rect 31444 8236 31450 8288
rect 32306 8236 32312 8288
rect 32364 8276 32370 8288
rect 34440 8276 34468 8316
rect 32364 8248 34468 8276
rect 35268 8276 35296 8316
rect 35728 8316 37320 8344
rect 37384 8316 38936 8344
rect 35728 8276 35756 8316
rect 35268 8248 35756 8276
rect 37292 8276 37320 8316
rect 38930 8304 38936 8316
rect 38988 8304 38994 8356
rect 37642 8276 37648 8288
rect 37292 8248 37648 8276
rect 32364 8236 32370 8248
rect 37642 8236 37648 8248
rect 37700 8236 37706 8288
rect 38102 8236 38108 8288
rect 38160 8276 38166 8288
rect 40052 8276 40080 8375
rect 40494 8372 40500 8384
rect 40552 8372 40558 8424
rect 48286 8412 48314 8452
rect 56226 8440 56232 8452
rect 56284 8440 56290 8492
rect 57057 8483 57115 8489
rect 57057 8449 57069 8483
rect 57103 8480 57115 8483
rect 57514 8480 57520 8492
rect 57103 8452 57520 8480
rect 57103 8449 57115 8452
rect 57057 8443 57115 8449
rect 57514 8440 57520 8452
rect 57572 8440 57578 8492
rect 58342 8480 58348 8492
rect 58303 8452 58348 8480
rect 58342 8440 58348 8452
rect 58400 8440 58406 8492
rect 58526 8412 58532 8424
rect 48286 8384 58532 8412
rect 58526 8372 58532 8384
rect 58584 8372 58590 8424
rect 58066 8344 58072 8356
rect 58027 8316 58072 8344
rect 58066 8304 58072 8316
rect 58124 8304 58130 8356
rect 38160 8248 40080 8276
rect 38160 8236 38166 8248
rect 56134 8236 56140 8288
rect 56192 8276 56198 8288
rect 57146 8276 57152 8288
rect 56192 8248 57152 8276
rect 56192 8236 56198 8248
rect 57146 8236 57152 8248
rect 57204 8236 57210 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 12069 8075 12127 8081
rect 12069 8041 12081 8075
rect 12115 8072 12127 8075
rect 12250 8072 12256 8084
rect 12115 8044 12256 8072
rect 12115 8041 12127 8044
rect 12069 8035 12127 8041
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17126 8072 17132 8084
rect 17000 8044 17132 8072
rect 17000 8032 17006 8044
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 17402 8032 17408 8084
rect 17460 8072 17466 8084
rect 17460 8044 20576 8072
rect 17460 8032 17466 8044
rect 11146 7964 11152 8016
rect 11204 8004 11210 8016
rect 11885 8007 11943 8013
rect 11885 8004 11897 8007
rect 11204 7976 11897 8004
rect 11204 7964 11210 7976
rect 11885 7973 11897 7976
rect 11931 7973 11943 8007
rect 11885 7967 11943 7973
rect 16850 7964 16856 8016
rect 16908 8004 16914 8016
rect 17313 8007 17371 8013
rect 17313 8004 17325 8007
rect 16908 7976 17325 8004
rect 16908 7964 16914 7976
rect 17313 7973 17325 7976
rect 17359 8004 17371 8007
rect 19150 8004 19156 8016
rect 17359 7976 19156 8004
rect 17359 7973 17371 7976
rect 17313 7967 17371 7973
rect 19150 7964 19156 7976
rect 19208 7964 19214 8016
rect 2682 7896 2688 7948
rect 2740 7936 2746 7948
rect 2740 7908 19380 7936
rect 2740 7896 2746 7908
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 11790 7868 11796 7880
rect 1627 7840 11796 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 16761 7871 16819 7877
rect 16761 7837 16773 7871
rect 16807 7837 16819 7871
rect 16761 7831 16819 7837
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7868 18383 7871
rect 19352 7868 19380 7908
rect 19426 7896 19432 7948
rect 19484 7936 19490 7948
rect 19521 7939 19579 7945
rect 19521 7936 19533 7939
rect 19484 7908 19533 7936
rect 19484 7896 19490 7908
rect 19521 7905 19533 7908
rect 19567 7905 19579 7939
rect 20548 7936 20576 8044
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 21450 8072 21456 8084
rect 20772 8044 21456 8072
rect 20772 8032 20778 8044
rect 21450 8032 21456 8044
rect 21508 8072 21514 8084
rect 32030 8072 32036 8084
rect 21508 8044 32036 8072
rect 21508 8032 21514 8044
rect 32030 8032 32036 8044
rect 32088 8032 32094 8084
rect 32122 8032 32128 8084
rect 32180 8072 32186 8084
rect 36630 8072 36636 8084
rect 32180 8044 36636 8072
rect 32180 8032 32186 8044
rect 36630 8032 36636 8044
rect 36688 8032 36694 8084
rect 38010 8032 38016 8084
rect 38068 8072 38074 8084
rect 38381 8075 38439 8081
rect 38381 8072 38393 8075
rect 38068 8044 38393 8072
rect 38068 8032 38074 8044
rect 38381 8041 38393 8044
rect 38427 8072 38439 8075
rect 38746 8072 38752 8084
rect 38427 8044 38752 8072
rect 38427 8041 38439 8044
rect 38381 8035 38439 8041
rect 38746 8032 38752 8044
rect 38804 8032 38810 8084
rect 38841 8075 38899 8081
rect 38841 8041 38853 8075
rect 38887 8072 38899 8075
rect 38930 8072 38936 8084
rect 38887 8044 38936 8072
rect 38887 8041 38899 8044
rect 38841 8035 38899 8041
rect 38930 8032 38936 8044
rect 38988 8032 38994 8084
rect 40126 8072 40132 8084
rect 40087 8044 40132 8072
rect 40126 8032 40132 8044
rect 40184 8032 40190 8084
rect 57238 8072 57244 8084
rect 55600 8044 57244 8072
rect 27154 7964 27160 8016
rect 27212 8004 27218 8016
rect 27522 8004 27528 8016
rect 27212 7976 27528 8004
rect 27212 7964 27218 7976
rect 27522 7964 27528 7976
rect 27580 8004 27586 8016
rect 28445 8007 28503 8013
rect 28445 8004 28457 8007
rect 27580 7976 28457 8004
rect 27580 7964 27586 7976
rect 28445 7973 28457 7976
rect 28491 7973 28503 8007
rect 28445 7967 28503 7973
rect 30745 8007 30803 8013
rect 30745 7973 30757 8007
rect 30791 8004 30803 8007
rect 30791 7976 32996 8004
rect 30791 7973 30803 7976
rect 30745 7967 30803 7973
rect 20548 7908 24072 7936
rect 19521 7899 19579 7905
rect 24044 7877 24072 7908
rect 23477 7871 23535 7877
rect 23477 7868 23489 7871
rect 18371 7840 19288 7868
rect 19352 7840 23489 7868
rect 18371 7837 18383 7840
rect 18325 7831 18383 7837
rect 1854 7800 1860 7812
rect 1815 7772 1860 7800
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 11609 7803 11667 7809
rect 11609 7769 11621 7803
rect 11655 7800 11667 7803
rect 12158 7800 12164 7812
rect 11655 7772 12164 7800
rect 11655 7769 11667 7772
rect 11609 7763 11667 7769
rect 12158 7760 12164 7772
rect 12216 7760 12222 7812
rect 16776 7800 16804 7831
rect 18601 7803 18659 7809
rect 18601 7800 18613 7803
rect 16776 7772 18613 7800
rect 18340 7744 18368 7772
rect 18601 7769 18613 7772
rect 18647 7769 18659 7803
rect 19260 7800 19288 7840
rect 23477 7837 23489 7840
rect 23523 7837 23535 7871
rect 23477 7831 23535 7837
rect 24029 7871 24087 7877
rect 24029 7837 24041 7871
rect 24075 7837 24087 7871
rect 24029 7831 24087 7837
rect 24670 7828 24676 7880
rect 24728 7868 24734 7880
rect 25133 7871 25191 7877
rect 25133 7868 25145 7871
rect 24728 7840 25145 7868
rect 24728 7828 24734 7840
rect 25133 7837 25145 7840
rect 25179 7837 25191 7871
rect 25133 7831 25191 7837
rect 27065 7871 27123 7877
rect 27065 7837 27077 7871
rect 27111 7868 27123 7871
rect 27172 7868 27200 7964
rect 30466 7936 30472 7948
rect 30024 7908 30472 7936
rect 30024 7877 30052 7908
rect 30466 7896 30472 7908
rect 30524 7896 30530 7948
rect 31018 7936 31024 7948
rect 30979 7908 31024 7936
rect 31018 7896 31024 7908
rect 31076 7896 31082 7948
rect 31202 7936 31208 7948
rect 31163 7908 31208 7936
rect 31202 7896 31208 7908
rect 31260 7896 31266 7948
rect 31478 7896 31484 7948
rect 31536 7936 31542 7948
rect 32122 7936 32128 7948
rect 31536 7908 31984 7936
rect 32083 7908 32128 7936
rect 31536 7896 31542 7908
rect 27111 7840 27200 7868
rect 30009 7871 30067 7877
rect 27111 7837 27123 7840
rect 27065 7831 27123 7837
rect 30009 7837 30021 7871
rect 30055 7837 30067 7871
rect 30009 7831 30067 7837
rect 30285 7871 30343 7877
rect 30285 7837 30297 7871
rect 30331 7868 30343 7871
rect 30742 7868 30748 7880
rect 30331 7840 30748 7868
rect 30331 7837 30343 7840
rect 30285 7831 30343 7837
rect 30742 7828 30748 7840
rect 30800 7828 30806 7880
rect 30834 7828 30840 7880
rect 30892 7868 30898 7880
rect 30929 7871 30987 7877
rect 30929 7868 30941 7871
rect 30892 7840 30941 7868
rect 30892 7828 30898 7840
rect 30929 7837 30941 7840
rect 30975 7837 30987 7871
rect 30929 7831 30987 7837
rect 31113 7871 31171 7877
rect 31113 7837 31125 7871
rect 31159 7868 31171 7871
rect 31570 7868 31576 7880
rect 31159 7840 31576 7868
rect 31159 7837 31171 7840
rect 31113 7831 31171 7837
rect 19610 7800 19616 7812
rect 19260 7772 19616 7800
rect 18601 7763 18659 7769
rect 19610 7760 19616 7772
rect 19668 7760 19674 7812
rect 19788 7803 19846 7809
rect 19788 7769 19800 7803
rect 19834 7800 19846 7803
rect 19978 7800 19984 7812
rect 19834 7772 19984 7800
rect 19834 7769 19846 7772
rect 19788 7763 19846 7769
rect 19978 7760 19984 7772
rect 20036 7760 20042 7812
rect 20346 7760 20352 7812
rect 20404 7800 20410 7812
rect 20530 7800 20536 7812
rect 20404 7772 20536 7800
rect 20404 7760 20410 7772
rect 20530 7760 20536 7772
rect 20588 7760 20594 7812
rect 23658 7800 23664 7812
rect 23619 7772 23664 7800
rect 23658 7760 23664 7772
rect 23716 7760 23722 7812
rect 25400 7803 25458 7809
rect 23768 7772 25360 7800
rect 17138 7735 17196 7741
rect 17138 7701 17150 7735
rect 17184 7732 17196 7735
rect 18230 7732 18236 7744
rect 17184 7704 18236 7732
rect 17184 7701 17196 7704
rect 17138 7695 17196 7701
rect 18230 7692 18236 7704
rect 18288 7692 18294 7744
rect 18322 7692 18328 7744
rect 18380 7692 18386 7744
rect 20898 7732 20904 7744
rect 20859 7704 20904 7732
rect 20898 7692 20904 7704
rect 20956 7692 20962 7744
rect 23768 7741 23796 7772
rect 23753 7735 23811 7741
rect 23753 7701 23765 7735
rect 23799 7701 23811 7735
rect 23753 7695 23811 7701
rect 23845 7735 23903 7741
rect 23845 7701 23857 7735
rect 23891 7732 23903 7735
rect 24854 7732 24860 7744
rect 23891 7704 24860 7732
rect 23891 7701 23903 7704
rect 23845 7695 23903 7701
rect 24854 7692 24860 7704
rect 24912 7692 24918 7744
rect 25332 7732 25360 7772
rect 25400 7769 25412 7803
rect 25446 7800 25458 7803
rect 25774 7800 25780 7812
rect 25446 7772 25780 7800
rect 25446 7769 25458 7772
rect 25400 7763 25458 7769
rect 25774 7760 25780 7772
rect 25832 7760 25838 7812
rect 26418 7760 26424 7812
rect 26476 7800 26482 7812
rect 27433 7803 27491 7809
rect 27433 7800 27445 7803
rect 26476 7772 27445 7800
rect 26476 7760 26482 7772
rect 27433 7769 27445 7772
rect 27479 7769 27491 7803
rect 27433 7763 27491 7769
rect 28261 7803 28319 7809
rect 28261 7769 28273 7803
rect 28307 7800 28319 7803
rect 28718 7800 28724 7812
rect 28307 7772 28724 7800
rect 28307 7769 28319 7772
rect 28261 7763 28319 7769
rect 28718 7760 28724 7772
rect 28776 7760 28782 7812
rect 29825 7803 29883 7809
rect 29825 7769 29837 7803
rect 29871 7800 29883 7803
rect 30944 7800 30972 7831
rect 31570 7828 31576 7840
rect 31628 7828 31634 7880
rect 31754 7828 31760 7880
rect 31812 7868 31818 7880
rect 31956 7868 31984 7908
rect 32122 7896 32128 7908
rect 32180 7896 32186 7948
rect 32217 7939 32275 7945
rect 32217 7905 32229 7939
rect 32263 7936 32275 7939
rect 32398 7936 32404 7948
rect 32263 7908 32404 7936
rect 32263 7905 32275 7908
rect 32217 7899 32275 7905
rect 32398 7896 32404 7908
rect 32456 7896 32462 7948
rect 32968 7945 32996 7976
rect 37274 7964 37280 8016
rect 37332 8004 37338 8016
rect 38473 8007 38531 8013
rect 37332 7976 38424 8004
rect 37332 7964 37338 7976
rect 38396 7948 38424 7976
rect 38473 7973 38485 8007
rect 38519 8004 38531 8007
rect 38519 7976 38884 8004
rect 38519 7973 38531 7976
rect 38473 7967 38531 7973
rect 38856 7948 38884 7976
rect 32953 7939 33011 7945
rect 32953 7905 32965 7939
rect 32999 7905 33011 7939
rect 32953 7899 33011 7905
rect 33318 7896 33324 7948
rect 33376 7936 33382 7948
rect 33413 7939 33471 7945
rect 33413 7936 33425 7939
rect 33376 7908 33425 7936
rect 33376 7896 33382 7908
rect 33413 7905 33425 7908
rect 33459 7905 33471 7939
rect 33413 7899 33471 7905
rect 33505 7939 33563 7945
rect 33505 7905 33517 7939
rect 33551 7936 33563 7939
rect 34146 7936 34152 7948
rect 33551 7908 34152 7936
rect 33551 7905 33563 7908
rect 33505 7899 33563 7905
rect 32309 7871 32367 7877
rect 32309 7868 32321 7871
rect 31812 7840 31857 7868
rect 31956 7840 32321 7868
rect 31812 7828 31818 7840
rect 32309 7837 32321 7840
rect 32355 7868 32367 7871
rect 33520 7868 33548 7899
rect 34146 7896 34152 7908
rect 34204 7896 34210 7948
rect 34885 7939 34943 7945
rect 34885 7905 34897 7939
rect 34931 7936 34943 7939
rect 35342 7936 35348 7948
rect 34931 7908 35348 7936
rect 34931 7905 34943 7908
rect 34885 7899 34943 7905
rect 35342 7896 35348 7908
rect 35400 7896 35406 7948
rect 36078 7896 36084 7948
rect 36136 7936 36142 7948
rect 36265 7939 36323 7945
rect 36265 7936 36277 7939
rect 36136 7908 36277 7936
rect 36136 7896 36142 7908
rect 36265 7905 36277 7908
rect 36311 7905 36323 7939
rect 38013 7939 38071 7945
rect 38013 7936 38025 7939
rect 36265 7899 36323 7905
rect 37200 7908 38025 7936
rect 37200 7877 37228 7908
rect 38013 7905 38025 7908
rect 38059 7936 38071 7939
rect 38194 7936 38200 7948
rect 38059 7908 38200 7936
rect 38059 7905 38071 7908
rect 38013 7899 38071 7905
rect 38194 7896 38200 7908
rect 38252 7896 38258 7948
rect 38378 7896 38384 7948
rect 38436 7936 38442 7948
rect 38565 7939 38623 7945
rect 38565 7936 38577 7939
rect 38436 7908 38577 7936
rect 38436 7896 38442 7908
rect 38565 7905 38577 7908
rect 38611 7905 38623 7939
rect 38565 7899 38623 7905
rect 38838 7896 38844 7948
rect 38896 7896 38902 7948
rect 39758 7896 39764 7948
rect 39816 7936 39822 7948
rect 39816 7908 40356 7936
rect 39816 7896 39822 7908
rect 35161 7871 35219 7877
rect 35161 7868 35173 7871
rect 32355 7840 33548 7868
rect 34992 7840 35173 7868
rect 32355 7837 32367 7840
rect 32309 7831 32367 7837
rect 34992 7812 35020 7840
rect 35161 7837 35173 7840
rect 35207 7837 35219 7871
rect 35161 7831 35219 7837
rect 37185 7871 37243 7877
rect 37185 7837 37197 7871
rect 37231 7837 37243 7871
rect 37185 7831 37243 7837
rect 37277 7871 37335 7877
rect 37277 7837 37289 7871
rect 37323 7837 37335 7871
rect 37277 7831 37335 7837
rect 33594 7800 33600 7812
rect 29871 7772 30788 7800
rect 30944 7772 33600 7800
rect 29871 7769 29883 7772
rect 29825 7763 29883 7769
rect 26142 7732 26148 7744
rect 25332 7704 26148 7732
rect 26142 7692 26148 7704
rect 26200 7732 26206 7744
rect 26513 7735 26571 7741
rect 26513 7732 26525 7735
rect 26200 7704 26525 7732
rect 26200 7692 26206 7704
rect 26513 7701 26525 7704
rect 26559 7701 26571 7735
rect 26513 7695 26571 7701
rect 28074 7692 28080 7744
rect 28132 7732 28138 7744
rect 29454 7732 29460 7744
rect 28132 7704 29460 7732
rect 28132 7692 28138 7704
rect 29454 7692 29460 7704
rect 29512 7732 29518 7744
rect 30193 7735 30251 7741
rect 30193 7732 30205 7735
rect 29512 7704 30205 7732
rect 29512 7692 29518 7704
rect 30193 7701 30205 7704
rect 30239 7701 30251 7735
rect 30760 7732 30788 7772
rect 33594 7760 33600 7772
rect 33652 7760 33658 7812
rect 34974 7760 34980 7812
rect 35032 7760 35038 7812
rect 37292 7800 37320 7831
rect 37366 7828 37372 7880
rect 37424 7868 37430 7880
rect 37461 7871 37519 7877
rect 37461 7868 37473 7871
rect 37424 7840 37473 7868
rect 37424 7828 37430 7840
rect 37461 7837 37473 7840
rect 37507 7837 37519 7871
rect 37461 7831 37519 7837
rect 37553 7871 37611 7877
rect 37553 7837 37565 7871
rect 37599 7868 37611 7871
rect 37734 7868 37740 7880
rect 37599 7840 37740 7868
rect 37599 7837 37611 7840
rect 37553 7831 37611 7837
rect 37734 7828 37740 7840
rect 37792 7828 37798 7880
rect 38102 7828 38108 7880
rect 38160 7868 38166 7880
rect 40328 7877 40356 7908
rect 40037 7871 40095 7877
rect 40037 7868 40049 7871
rect 38160 7840 40049 7868
rect 38160 7828 38166 7840
rect 40037 7837 40049 7840
rect 40083 7837 40095 7871
rect 40037 7831 40095 7837
rect 40313 7871 40371 7877
rect 40313 7837 40325 7871
rect 40359 7868 40371 7871
rect 55306 7868 55312 7880
rect 40359 7840 55312 7868
rect 40359 7837 40371 7840
rect 40313 7831 40371 7837
rect 55306 7828 55312 7840
rect 55364 7828 55370 7880
rect 55493 7871 55551 7877
rect 55493 7837 55505 7871
rect 55539 7868 55551 7871
rect 55600 7868 55628 8044
rect 57238 8032 57244 8044
rect 57296 8032 57302 8084
rect 56137 8007 56195 8013
rect 56137 7973 56149 8007
rect 56183 7973 56195 8007
rect 56137 7967 56195 7973
rect 56152 7936 56180 7967
rect 56870 7936 56876 7948
rect 56152 7908 56640 7936
rect 56831 7908 56876 7936
rect 55539 7840 55628 7868
rect 55677 7871 55735 7877
rect 55539 7837 55551 7840
rect 55493 7831 55551 7837
rect 55677 7837 55689 7871
rect 55723 7868 55735 7871
rect 55723 7840 56364 7868
rect 55723 7837 55735 7840
rect 55677 7831 55735 7837
rect 39758 7800 39764 7812
rect 37292 7772 39764 7800
rect 39758 7760 39764 7772
rect 39816 7760 39822 7812
rect 40126 7760 40132 7812
rect 40184 7800 40190 7812
rect 50154 7800 50160 7812
rect 40184 7772 50160 7800
rect 40184 7760 40190 7772
rect 50154 7760 50160 7772
rect 50212 7760 50218 7812
rect 56134 7800 56140 7812
rect 56095 7772 56140 7800
rect 56134 7760 56140 7772
rect 56192 7760 56198 7812
rect 56336 7800 56364 7840
rect 56410 7828 56416 7880
rect 56468 7868 56474 7880
rect 56612 7868 56640 7908
rect 56870 7896 56876 7908
rect 56928 7896 56934 7948
rect 57129 7871 57187 7877
rect 57129 7868 57141 7871
rect 56468 7840 56513 7868
rect 56612 7840 57141 7868
rect 56468 7828 56474 7840
rect 57129 7837 57141 7840
rect 57175 7837 57187 7871
rect 57129 7831 57187 7837
rect 56336 7772 56548 7800
rect 56520 7744 56548 7772
rect 31662 7732 31668 7744
rect 30760 7704 31668 7732
rect 30193 7695 30251 7701
rect 31662 7692 31668 7704
rect 31720 7692 31726 7744
rect 33137 7735 33195 7741
rect 33137 7701 33149 7735
rect 33183 7732 33195 7735
rect 36906 7732 36912 7744
rect 33183 7704 36912 7732
rect 33183 7701 33195 7704
rect 33137 7695 33195 7701
rect 36906 7692 36912 7704
rect 36964 7692 36970 7744
rect 37001 7735 37059 7741
rect 37001 7701 37013 7735
rect 37047 7732 37059 7735
rect 38010 7732 38016 7744
rect 37047 7704 38016 7732
rect 37047 7701 37059 7704
rect 37001 7695 37059 7701
rect 38010 7692 38016 7704
rect 38068 7692 38074 7744
rect 55677 7735 55735 7741
rect 55677 7701 55689 7735
rect 55723 7732 55735 7735
rect 56321 7735 56379 7741
rect 56321 7732 56333 7735
rect 55723 7704 56333 7732
rect 55723 7701 55735 7704
rect 55677 7695 55735 7701
rect 56321 7701 56333 7704
rect 56367 7701 56379 7735
rect 56321 7695 56379 7701
rect 56502 7692 56508 7744
rect 56560 7732 56566 7744
rect 58253 7735 58311 7741
rect 58253 7732 58265 7735
rect 56560 7704 58265 7732
rect 56560 7692 56566 7704
rect 58253 7701 58265 7704
rect 58299 7701 58311 7735
rect 58253 7695 58311 7701
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 11790 7528 11796 7540
rect 11751 7500 11796 7528
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 13262 7528 13268 7540
rect 13223 7500 13268 7528
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 17865 7531 17923 7537
rect 17865 7497 17877 7531
rect 17911 7528 17923 7531
rect 17954 7528 17960 7540
rect 17911 7500 17960 7528
rect 17911 7497 17923 7500
rect 17865 7491 17923 7497
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 19426 7488 19432 7540
rect 19484 7528 19490 7540
rect 23750 7528 23756 7540
rect 19484 7500 23756 7528
rect 19484 7488 19490 7500
rect 23750 7488 23756 7500
rect 23808 7528 23814 7540
rect 24670 7528 24676 7540
rect 23808 7500 24676 7528
rect 23808 7488 23814 7500
rect 24670 7488 24676 7500
rect 24728 7488 24734 7540
rect 24762 7488 24768 7540
rect 24820 7528 24826 7540
rect 28353 7531 28411 7537
rect 28353 7528 28365 7531
rect 24820 7500 28365 7528
rect 24820 7488 24826 7500
rect 28353 7497 28365 7500
rect 28399 7497 28411 7531
rect 28353 7491 28411 7497
rect 30926 7488 30932 7540
rect 30984 7528 30990 7540
rect 31205 7531 31263 7537
rect 31205 7528 31217 7531
rect 30984 7500 31217 7528
rect 30984 7488 30990 7500
rect 31205 7497 31217 7500
rect 31251 7497 31263 7531
rect 32398 7528 32404 7540
rect 32359 7500 32404 7528
rect 31205 7491 31263 7497
rect 32398 7488 32404 7500
rect 32456 7488 32462 7540
rect 33781 7531 33839 7537
rect 33781 7497 33793 7531
rect 33827 7497 33839 7531
rect 34974 7528 34980 7540
rect 34935 7500 34980 7528
rect 33781 7491 33839 7497
rect 7650 7420 7656 7472
rect 7708 7460 7714 7472
rect 18233 7463 18291 7469
rect 18233 7460 18245 7463
rect 7708 7432 18245 7460
rect 7708 7420 7714 7432
rect 18233 7429 18245 7432
rect 18279 7429 18291 7463
rect 18233 7423 18291 7429
rect 18325 7463 18383 7469
rect 18325 7429 18337 7463
rect 18371 7460 18383 7463
rect 23385 7463 23443 7469
rect 18371 7432 22094 7460
rect 18371 7429 18383 7432
rect 18325 7423 18383 7429
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 11054 7392 11060 7404
rect 1627 7364 11060 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 11054 7352 11060 7364
rect 11112 7352 11118 7404
rect 11974 7392 11980 7404
rect 11935 7364 11980 7392
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7392 12219 7395
rect 12805 7395 12863 7401
rect 12805 7392 12817 7395
rect 12207 7364 12817 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 12805 7361 12817 7364
rect 12851 7392 12863 7395
rect 13262 7392 13268 7404
rect 12851 7364 13268 7392
rect 12851 7361 12863 7364
rect 12805 7355 12863 7361
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 20346 7392 20352 7404
rect 20307 7364 20352 7392
rect 20346 7352 20352 7364
rect 20404 7352 20410 7404
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7392 20499 7395
rect 20898 7392 20904 7404
rect 20487 7364 20904 7392
rect 20487 7361 20499 7364
rect 20441 7355 20499 7361
rect 1762 7324 1768 7336
rect 1723 7296 1768 7324
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 12069 7327 12127 7333
rect 12069 7293 12081 7327
rect 12115 7293 12127 7327
rect 12250 7324 12256 7336
rect 12211 7296 12256 7324
rect 12069 7287 12127 7293
rect 12084 7188 12112 7287
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 18506 7324 18512 7336
rect 18467 7296 18512 7324
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 13078 7256 13084 7268
rect 13039 7228 13084 7256
rect 13078 7216 13084 7228
rect 13136 7216 13142 7268
rect 18690 7216 18696 7268
rect 18748 7256 18754 7268
rect 18874 7256 18880 7268
rect 18748 7228 18880 7256
rect 18748 7216 18754 7228
rect 18874 7216 18880 7228
rect 18932 7256 18938 7268
rect 19794 7256 19800 7268
rect 18932 7228 19800 7256
rect 18932 7216 18938 7228
rect 19794 7216 19800 7228
rect 19852 7216 19858 7268
rect 19978 7256 19984 7268
rect 19939 7228 19984 7256
rect 19978 7216 19984 7228
rect 20036 7216 20042 7268
rect 20456 7188 20484 7355
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 22066 7392 22094 7432
rect 23385 7429 23397 7463
rect 23431 7460 23443 7463
rect 29914 7460 29920 7472
rect 23431 7432 29920 7460
rect 23431 7429 23443 7432
rect 23385 7423 23443 7429
rect 29914 7420 29920 7432
rect 29972 7420 29978 7472
rect 33796 7460 33824 7491
rect 34974 7488 34980 7500
rect 35032 7488 35038 7540
rect 35158 7488 35164 7540
rect 35216 7528 35222 7540
rect 36078 7528 36084 7540
rect 35216 7500 36084 7528
rect 35216 7488 35222 7500
rect 36078 7488 36084 7500
rect 36136 7488 36142 7540
rect 36906 7488 36912 7540
rect 36964 7528 36970 7540
rect 36964 7500 38884 7528
rect 36964 7488 36970 7500
rect 38654 7460 38660 7472
rect 32324 7432 33180 7460
rect 33796 7432 38660 7460
rect 32324 7404 32352 7432
rect 25498 7392 25504 7404
rect 22066 7364 25504 7392
rect 25498 7352 25504 7364
rect 25556 7352 25562 7404
rect 27154 7392 27160 7404
rect 27115 7364 27160 7392
rect 27154 7352 27160 7364
rect 27212 7392 27218 7404
rect 28074 7392 28080 7404
rect 27212 7364 28080 7392
rect 27212 7352 27218 7364
rect 28074 7352 28080 7364
rect 28132 7352 28138 7404
rect 32306 7392 32312 7404
rect 32267 7364 32312 7392
rect 32306 7352 32312 7364
rect 32364 7352 32370 7404
rect 32398 7352 32404 7404
rect 32456 7392 32462 7404
rect 33152 7401 33180 7432
rect 38654 7420 38660 7432
rect 38712 7420 38718 7472
rect 32493 7395 32551 7401
rect 32493 7392 32505 7395
rect 32456 7364 32505 7392
rect 32456 7352 32462 7364
rect 32493 7361 32505 7364
rect 32539 7361 32551 7395
rect 32493 7355 32551 7361
rect 33137 7395 33195 7401
rect 33137 7361 33149 7395
rect 33183 7361 33195 7395
rect 33137 7355 33195 7361
rect 33226 7352 33232 7404
rect 33284 7392 33290 7404
rect 33321 7395 33379 7401
rect 33321 7392 33333 7395
rect 33284 7364 33333 7392
rect 33284 7352 33290 7364
rect 33321 7361 33333 7364
rect 33367 7361 33379 7395
rect 33321 7355 33379 7361
rect 33410 7352 33416 7404
rect 33468 7392 33474 7404
rect 33597 7395 33655 7401
rect 33597 7392 33609 7395
rect 33468 7364 33609 7392
rect 33468 7352 33474 7364
rect 33597 7361 33609 7364
rect 33643 7361 33655 7395
rect 34146 7392 34152 7404
rect 34107 7364 34152 7392
rect 33597 7355 33655 7361
rect 34146 7352 34152 7364
rect 34204 7352 34210 7404
rect 34606 7352 34612 7404
rect 34664 7392 34670 7404
rect 35253 7395 35311 7401
rect 35253 7392 35265 7395
rect 34664 7364 35265 7392
rect 34664 7352 34670 7364
rect 35253 7361 35265 7364
rect 35299 7361 35311 7395
rect 35253 7355 35311 7361
rect 35345 7395 35403 7401
rect 35345 7361 35357 7395
rect 35391 7361 35403 7395
rect 35345 7355 35403 7361
rect 20622 7324 20628 7336
rect 20583 7296 20628 7324
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 23198 7284 23204 7336
rect 23256 7324 23262 7336
rect 28534 7324 28540 7336
rect 23256 7296 28540 7324
rect 23256 7284 23262 7296
rect 28534 7284 28540 7296
rect 28592 7284 28598 7336
rect 28626 7284 28632 7336
rect 28684 7324 28690 7336
rect 33778 7324 33784 7336
rect 28684 7296 33784 7324
rect 28684 7284 28690 7296
rect 33778 7284 33784 7296
rect 33836 7284 33842 7336
rect 34057 7327 34115 7333
rect 34057 7293 34069 7327
rect 34103 7293 34115 7327
rect 34057 7287 34115 7293
rect 21358 7216 21364 7268
rect 21416 7256 21422 7268
rect 33137 7259 33195 7265
rect 21416 7228 33088 7256
rect 21416 7216 21422 7228
rect 12084 7160 20484 7188
rect 20530 7148 20536 7200
rect 20588 7188 20594 7200
rect 30834 7188 30840 7200
rect 20588 7160 30840 7188
rect 20588 7148 20594 7160
rect 30834 7148 30840 7160
rect 30892 7148 30898 7200
rect 31202 7148 31208 7200
rect 31260 7188 31266 7200
rect 32582 7188 32588 7200
rect 31260 7160 32588 7188
rect 31260 7148 31266 7160
rect 32582 7148 32588 7160
rect 32640 7148 32646 7200
rect 33060 7188 33088 7228
rect 33137 7225 33149 7259
rect 33183 7256 33195 7259
rect 34072 7256 34100 7287
rect 34514 7284 34520 7336
rect 34572 7324 34578 7336
rect 35360 7324 35388 7355
rect 35434 7352 35440 7404
rect 35492 7392 35498 7404
rect 35621 7395 35679 7401
rect 35492 7364 35537 7392
rect 35492 7352 35498 7364
rect 35621 7361 35633 7395
rect 35667 7392 35679 7395
rect 35894 7392 35900 7404
rect 35667 7364 35900 7392
rect 35667 7361 35679 7364
rect 35621 7355 35679 7361
rect 35894 7352 35900 7364
rect 35952 7352 35958 7404
rect 37550 7392 37556 7404
rect 37511 7364 37556 7392
rect 37550 7352 37556 7364
rect 37608 7352 37614 7404
rect 37645 7395 37703 7401
rect 37645 7361 37657 7395
rect 37691 7392 37703 7395
rect 38286 7392 38292 7404
rect 37691 7364 38292 7392
rect 37691 7361 37703 7364
rect 37645 7355 37703 7361
rect 38286 7352 38292 7364
rect 38344 7352 38350 7404
rect 38746 7392 38752 7404
rect 38707 7364 38752 7392
rect 38746 7352 38752 7364
rect 38804 7352 38810 7404
rect 38856 7392 38884 7500
rect 39316 7500 58388 7528
rect 39025 7395 39083 7401
rect 38856 7364 38976 7392
rect 35526 7324 35532 7336
rect 34572 7296 35532 7324
rect 34572 7284 34578 7296
rect 35526 7284 35532 7296
rect 35584 7284 35590 7336
rect 37369 7327 37427 7333
rect 37369 7293 37381 7327
rect 37415 7324 37427 7327
rect 37734 7324 37740 7336
rect 37415 7296 37740 7324
rect 37415 7293 37427 7296
rect 37369 7287 37427 7293
rect 37734 7284 37740 7296
rect 37792 7284 37798 7336
rect 38838 7324 38844 7336
rect 38799 7296 38844 7324
rect 38838 7284 38844 7296
rect 38896 7284 38902 7336
rect 38948 7324 38976 7364
rect 39025 7361 39037 7395
rect 39071 7392 39083 7395
rect 39206 7392 39212 7404
rect 39071 7364 39212 7392
rect 39071 7361 39083 7364
rect 39025 7355 39083 7361
rect 39206 7352 39212 7364
rect 39264 7352 39270 7404
rect 39316 7324 39344 7500
rect 39758 7460 39764 7472
rect 39719 7432 39764 7460
rect 39758 7420 39764 7432
rect 39816 7420 39822 7472
rect 41386 7432 45554 7460
rect 39666 7392 39672 7404
rect 39579 7364 39672 7392
rect 39666 7352 39672 7364
rect 39724 7392 39730 7404
rect 41386 7392 41414 7432
rect 39724 7364 41414 7392
rect 45526 7392 45554 7432
rect 50154 7420 50160 7472
rect 50212 7460 50218 7472
rect 50212 7432 57100 7460
rect 50212 7420 50218 7432
rect 53558 7392 53564 7404
rect 45526 7364 53564 7392
rect 39724 7352 39730 7364
rect 53558 7352 53564 7364
rect 53616 7352 53622 7404
rect 56137 7395 56195 7401
rect 56137 7361 56149 7395
rect 56183 7392 56195 7395
rect 56502 7392 56508 7404
rect 56183 7364 56508 7392
rect 56183 7361 56195 7364
rect 56137 7355 56195 7361
rect 56502 7352 56508 7364
rect 56560 7352 56566 7404
rect 57072 7401 57100 7432
rect 57238 7420 57244 7472
rect 57296 7460 57302 7472
rect 57333 7463 57391 7469
rect 57333 7460 57345 7463
rect 57296 7432 57345 7460
rect 57296 7420 57302 7432
rect 57333 7429 57345 7432
rect 57379 7460 57391 7463
rect 57422 7460 57428 7472
rect 57379 7432 57428 7460
rect 57379 7429 57391 7432
rect 57333 7423 57391 7429
rect 57422 7420 57428 7432
rect 57480 7420 57486 7472
rect 57606 7420 57612 7472
rect 57664 7460 57670 7472
rect 58253 7463 58311 7469
rect 58253 7460 58265 7463
rect 57664 7432 58265 7460
rect 57664 7420 57670 7432
rect 58253 7429 58265 7432
rect 58299 7429 58311 7463
rect 58253 7423 58311 7429
rect 57057 7395 57115 7401
rect 57057 7361 57069 7395
rect 57103 7361 57115 7395
rect 57057 7355 57115 7361
rect 57146 7352 57152 7404
rect 57204 7392 57210 7404
rect 58360 7401 58388 7500
rect 58069 7395 58127 7401
rect 58069 7392 58081 7395
rect 57204 7364 58081 7392
rect 57204 7352 57210 7364
rect 58069 7361 58081 7364
rect 58115 7361 58127 7395
rect 58069 7355 58127 7361
rect 58345 7395 58403 7401
rect 58345 7361 58357 7395
rect 58391 7361 58403 7395
rect 58345 7355 58403 7361
rect 38948 7296 39344 7324
rect 39942 7284 39948 7336
rect 40000 7324 40006 7336
rect 56226 7324 56232 7336
rect 40000 7296 56232 7324
rect 40000 7284 40006 7296
rect 56226 7284 56232 7296
rect 56284 7284 56290 7336
rect 56410 7324 56416 7336
rect 56371 7296 56416 7324
rect 56410 7284 56416 7296
rect 56468 7284 56474 7336
rect 33183 7228 34100 7256
rect 33183 7225 33195 7228
rect 33137 7219 33195 7225
rect 34698 7216 34704 7268
rect 34756 7256 34762 7268
rect 35158 7256 35164 7268
rect 34756 7228 35164 7256
rect 34756 7216 34762 7228
rect 35158 7216 35164 7228
rect 35216 7216 35222 7268
rect 39206 7216 39212 7268
rect 39264 7256 39270 7268
rect 55398 7256 55404 7268
rect 39264 7228 39309 7256
rect 47044 7228 55404 7256
rect 39264 7216 39270 7228
rect 33870 7188 33876 7200
rect 33060 7160 33876 7188
rect 33870 7148 33876 7160
rect 33928 7188 33934 7200
rect 34606 7188 34612 7200
rect 33928 7160 34612 7188
rect 33928 7148 33934 7160
rect 34606 7148 34612 7160
rect 34664 7148 34670 7200
rect 35250 7148 35256 7200
rect 35308 7188 35314 7200
rect 35526 7188 35532 7200
rect 35308 7160 35532 7188
rect 35308 7148 35314 7160
rect 35526 7148 35532 7160
rect 35584 7148 35590 7200
rect 37182 7148 37188 7200
rect 37240 7188 37246 7200
rect 37829 7191 37887 7197
rect 37829 7188 37841 7191
rect 37240 7160 37841 7188
rect 37240 7148 37246 7160
rect 37829 7157 37841 7160
rect 37875 7157 37887 7191
rect 38378 7188 38384 7200
rect 38339 7160 38384 7188
rect 37829 7151 37887 7157
rect 38378 7148 38384 7160
rect 38436 7188 38442 7200
rect 38654 7188 38660 7200
rect 38436 7160 38660 7188
rect 38436 7148 38442 7160
rect 38654 7148 38660 7160
rect 38712 7188 38718 7200
rect 38749 7191 38807 7197
rect 38749 7188 38761 7191
rect 38712 7160 38761 7188
rect 38712 7148 38718 7160
rect 38749 7157 38761 7160
rect 38795 7157 38807 7191
rect 38749 7151 38807 7157
rect 38838 7148 38844 7200
rect 38896 7188 38902 7200
rect 47044 7188 47072 7228
rect 55398 7216 55404 7228
rect 55456 7216 55462 7268
rect 38896 7160 47072 7188
rect 38896 7148 38902 7160
rect 47118 7148 47124 7200
rect 47176 7188 47182 7200
rect 56594 7188 56600 7200
rect 47176 7160 56600 7188
rect 47176 7148 47182 7160
rect 56594 7148 56600 7160
rect 56652 7148 56658 7200
rect 57514 7148 57520 7200
rect 57572 7188 57578 7200
rect 58069 7191 58127 7197
rect 58069 7188 58081 7191
rect 57572 7160 58081 7188
rect 57572 7148 57578 7160
rect 58069 7157 58081 7160
rect 58115 7157 58127 7191
rect 58069 7151 58127 7157
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 16850 6944 16856 6996
rect 16908 6984 16914 6996
rect 20530 6984 20536 6996
rect 16908 6956 20536 6984
rect 16908 6944 16914 6956
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 23566 6984 23572 6996
rect 23479 6956 23572 6984
rect 13633 6919 13691 6925
rect 13633 6885 13645 6919
rect 13679 6885 13691 6919
rect 13633 6879 13691 6885
rect 15197 6919 15255 6925
rect 15197 6885 15209 6919
rect 15243 6885 15255 6919
rect 15197 6879 15255 6885
rect 11054 6848 11060 6860
rect 11015 6820 11060 6848
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 11238 6848 11244 6860
rect 11199 6820 11244 6848
rect 11238 6808 11244 6820
rect 11296 6808 11302 6860
rect 11333 6851 11391 6857
rect 11333 6817 11345 6851
rect 11379 6848 11391 6851
rect 13538 6848 13544 6860
rect 11379 6820 13544 6848
rect 11379 6817 11391 6820
rect 11333 6811 11391 6817
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 13648 6848 13676 6879
rect 13814 6848 13820 6860
rect 13648 6820 13820 6848
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 13998 6808 14004 6860
rect 14056 6848 14062 6860
rect 15212 6848 15240 6879
rect 19242 6876 19248 6928
rect 19300 6916 19306 6928
rect 19300 6888 20392 6916
rect 19300 6876 19306 6888
rect 14056 6820 15240 6848
rect 14056 6808 14062 6820
rect 15286 6808 15292 6860
rect 15344 6848 15350 6860
rect 15381 6851 15439 6857
rect 15381 6848 15393 6851
rect 15344 6820 15393 6848
rect 15344 6808 15350 6820
rect 15381 6817 15393 6820
rect 15427 6817 15439 6851
rect 15381 6811 15439 6817
rect 18230 6808 18236 6860
rect 18288 6848 18294 6860
rect 20162 6848 20168 6860
rect 18288 6820 20168 6848
rect 18288 6808 18294 6820
rect 20162 6808 20168 6820
rect 20220 6808 20226 6860
rect 20364 6848 20392 6888
rect 20438 6876 20444 6928
rect 20496 6916 20502 6928
rect 21358 6916 21364 6928
rect 20496 6888 21364 6916
rect 20496 6876 20502 6888
rect 21358 6876 21364 6888
rect 21416 6876 21422 6928
rect 22370 6916 22376 6928
rect 22331 6888 22376 6916
rect 22370 6876 22376 6888
rect 22428 6876 22434 6928
rect 23492 6925 23520 6956
rect 23566 6944 23572 6956
rect 23624 6984 23630 6996
rect 26602 6984 26608 6996
rect 23624 6956 26608 6984
rect 23624 6944 23630 6956
rect 26602 6944 26608 6956
rect 26660 6944 26666 6996
rect 26786 6944 26792 6996
rect 26844 6984 26850 6996
rect 38378 6984 38384 6996
rect 26844 6956 38384 6984
rect 26844 6944 26850 6956
rect 38378 6944 38384 6956
rect 38436 6944 38442 6996
rect 38654 6944 38660 6996
rect 38712 6984 38718 6996
rect 47118 6984 47124 6996
rect 38712 6956 47124 6984
rect 38712 6944 38718 6956
rect 47118 6944 47124 6956
rect 47176 6944 47182 6996
rect 23477 6919 23535 6925
rect 22480 6888 23060 6916
rect 22480 6848 22508 6888
rect 20364 6820 22508 6848
rect 22830 6808 22836 6860
rect 22888 6848 22894 6860
rect 23032 6848 23060 6888
rect 23477 6885 23489 6919
rect 23523 6885 23535 6919
rect 23934 6916 23940 6928
rect 23477 6879 23535 6885
rect 23860 6888 23940 6916
rect 22888 6820 22968 6848
rect 23032 6820 23787 6848
rect 22888 6808 22894 6820
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 9398 6780 9404 6792
rect 1627 6752 2774 6780
rect 9359 6752 9404 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 1854 6712 1860 6724
rect 1815 6684 1860 6712
rect 1854 6672 1860 6684
rect 1912 6672 1918 6724
rect 2746 6712 2774 6752
rect 9398 6740 9404 6752
rect 9456 6740 9462 6792
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 9677 6783 9735 6789
rect 9548 6752 9593 6780
rect 9548 6740 9554 6752
rect 9677 6749 9689 6783
rect 9723 6780 9735 6783
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 9723 6752 11437 6780
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 11072 6724 11100 6752
rect 11425 6749 11437 6752
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 11514 6740 11520 6792
rect 11572 6780 11578 6792
rect 13262 6780 13268 6792
rect 11572 6752 11617 6780
rect 13223 6752 13268 6780
rect 11572 6740 11578 6752
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 22094 6780 22100 6792
rect 17696 6752 22100 6780
rect 9950 6712 9956 6724
rect 2746 6684 9956 6712
rect 9950 6672 9956 6684
rect 10008 6672 10014 6724
rect 10134 6712 10140 6724
rect 10095 6684 10140 6712
rect 10134 6672 10140 6684
rect 10192 6672 10198 6724
rect 11054 6672 11060 6724
rect 11112 6672 11118 6724
rect 13280 6712 13308 6740
rect 14921 6715 14979 6721
rect 14921 6712 14933 6715
rect 13280 6684 14933 6712
rect 14921 6681 14933 6684
rect 14967 6681 14979 6715
rect 14921 6675 14979 6681
rect 13725 6647 13783 6653
rect 13725 6613 13737 6647
rect 13771 6644 13783 6647
rect 17696 6644 17724 6752
rect 22094 6740 22100 6752
rect 22152 6740 22158 6792
rect 22940 6789 22968 6820
rect 22695 6783 22753 6789
rect 22695 6749 22707 6783
rect 22741 6780 22753 6783
rect 22925 6783 22983 6789
rect 22741 6752 22876 6780
rect 22741 6749 22753 6752
rect 22695 6743 22753 6749
rect 19429 6715 19487 6721
rect 19429 6681 19441 6715
rect 19475 6712 19487 6715
rect 20070 6712 20076 6724
rect 19475 6684 20076 6712
rect 19475 6681 19487 6684
rect 19429 6675 19487 6681
rect 20070 6672 20076 6684
rect 20128 6672 20134 6724
rect 22554 6712 22560 6724
rect 22515 6684 22560 6712
rect 22554 6672 22560 6684
rect 22612 6672 22618 6724
rect 13771 6616 17724 6644
rect 13771 6613 13783 6616
rect 13725 6607 13783 6613
rect 17770 6604 17776 6656
rect 17828 6644 17834 6656
rect 19978 6644 19984 6656
rect 17828 6616 19984 6644
rect 17828 6604 17834 6616
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 22370 6604 22376 6656
rect 22428 6644 22434 6656
rect 22741 6647 22799 6653
rect 22741 6644 22753 6647
rect 22428 6616 22753 6644
rect 22428 6604 22434 6616
rect 22741 6613 22753 6616
rect 22787 6613 22799 6647
rect 22848 6644 22876 6752
rect 22925 6749 22937 6783
rect 22971 6749 22983 6783
rect 22925 6743 22983 6749
rect 23014 6740 23020 6792
rect 23072 6780 23078 6792
rect 23759 6789 23787 6820
rect 23661 6783 23719 6789
rect 23661 6780 23673 6783
rect 23072 6752 23673 6780
rect 23072 6740 23078 6752
rect 23661 6749 23673 6752
rect 23707 6749 23719 6783
rect 23661 6743 23719 6749
rect 23752 6783 23810 6789
rect 23752 6749 23764 6783
rect 23798 6749 23810 6783
rect 23860 6780 23888 6888
rect 23934 6876 23940 6888
rect 23992 6876 23998 6928
rect 24026 6876 24032 6928
rect 24084 6916 24090 6928
rect 35894 6916 35900 6928
rect 24084 6888 24164 6916
rect 24084 6876 24090 6888
rect 23937 6783 23995 6789
rect 23937 6780 23949 6783
rect 23860 6752 23949 6780
rect 23752 6743 23810 6749
rect 23937 6749 23949 6752
rect 23983 6749 23995 6783
rect 23937 6743 23995 6749
rect 24024 6783 24082 6789
rect 24024 6749 24036 6783
rect 24070 6780 24082 6783
rect 24136 6780 24164 6888
rect 31036 6888 31616 6916
rect 24578 6848 24584 6860
rect 24539 6820 24584 6848
rect 24578 6808 24584 6820
rect 24636 6808 24642 6860
rect 27614 6808 27620 6860
rect 27672 6848 27678 6860
rect 28166 6848 28172 6860
rect 27672 6820 28172 6848
rect 27672 6808 27678 6820
rect 28166 6808 28172 6820
rect 28224 6848 28230 6860
rect 29178 6848 29184 6860
rect 28224 6820 28764 6848
rect 28224 6808 28230 6820
rect 25130 6780 25136 6792
rect 24070 6752 24164 6780
rect 25091 6752 25136 6780
rect 24070 6749 24082 6752
rect 24024 6743 24082 6749
rect 25130 6740 25136 6752
rect 25188 6740 25194 6792
rect 26421 6783 26479 6789
rect 26421 6749 26433 6783
rect 26467 6780 26479 6783
rect 28074 6780 28080 6792
rect 26467 6752 28080 6780
rect 26467 6749 26479 6752
rect 26421 6743 26479 6749
rect 28074 6740 28080 6752
rect 28132 6740 28138 6792
rect 28626 6780 28632 6792
rect 28587 6752 28632 6780
rect 28626 6740 28632 6752
rect 28684 6740 28690 6792
rect 28736 6789 28764 6820
rect 28828 6820 29184 6848
rect 28828 6789 28856 6820
rect 29178 6808 29184 6820
rect 29236 6808 29242 6860
rect 31036 6848 31064 6888
rect 31478 6848 31484 6860
rect 30576 6820 31064 6848
rect 31439 6820 31484 6848
rect 30576 6792 30604 6820
rect 31478 6808 31484 6820
rect 31536 6808 31542 6860
rect 31588 6848 31616 6888
rect 33060 6888 35900 6916
rect 31662 6848 31668 6860
rect 31575 6820 31668 6848
rect 31662 6808 31668 6820
rect 31720 6848 31726 6860
rect 32677 6851 32735 6857
rect 32677 6848 32689 6851
rect 31720 6820 32689 6848
rect 31720 6808 31726 6820
rect 32677 6817 32689 6820
rect 32723 6848 32735 6851
rect 33060 6848 33088 6888
rect 35894 6876 35900 6888
rect 35952 6916 35958 6928
rect 37366 6916 37372 6928
rect 35952 6888 37372 6916
rect 35952 6876 35958 6888
rect 37366 6876 37372 6888
rect 37424 6876 37430 6928
rect 37550 6876 37556 6928
rect 37608 6916 37614 6928
rect 39666 6916 39672 6928
rect 37608 6888 39672 6916
rect 37608 6876 37614 6888
rect 39666 6876 39672 6888
rect 39724 6876 39730 6928
rect 32723 6820 33088 6848
rect 34333 6851 34391 6857
rect 32723 6817 32735 6820
rect 32677 6811 32735 6817
rect 34333 6817 34345 6851
rect 34379 6848 34391 6851
rect 35434 6848 35440 6860
rect 34379 6820 35440 6848
rect 34379 6817 34391 6820
rect 34333 6811 34391 6817
rect 35434 6808 35440 6820
rect 35492 6808 35498 6860
rect 35989 6851 36047 6857
rect 35989 6817 36001 6851
rect 36035 6848 36047 6851
rect 36170 6848 36176 6860
rect 36035 6820 36176 6848
rect 36035 6817 36047 6820
rect 35989 6811 36047 6817
rect 36170 6808 36176 6820
rect 36228 6808 36234 6860
rect 37182 6848 37188 6860
rect 37143 6820 37188 6848
rect 37182 6808 37188 6820
rect 37240 6808 37246 6860
rect 37826 6848 37832 6860
rect 37787 6820 37832 6848
rect 37826 6808 37832 6820
rect 37884 6808 37890 6860
rect 38010 6808 38016 6860
rect 38068 6848 38074 6860
rect 39022 6848 39028 6860
rect 38068 6820 38516 6848
rect 38983 6820 39028 6848
rect 38068 6808 38074 6820
rect 28721 6783 28779 6789
rect 28721 6749 28733 6783
rect 28767 6749 28779 6783
rect 28721 6743 28779 6749
rect 28813 6783 28871 6789
rect 28813 6749 28825 6783
rect 28859 6749 28871 6783
rect 28813 6743 28871 6749
rect 28997 6783 29055 6789
rect 28997 6749 29009 6783
rect 29043 6780 29055 6783
rect 30374 6780 30380 6792
rect 29043 6752 30380 6780
rect 29043 6749 29055 6752
rect 28997 6743 29055 6749
rect 30374 6740 30380 6752
rect 30432 6780 30438 6792
rect 30558 6780 30564 6792
rect 30432 6752 30564 6780
rect 30432 6740 30438 6752
rect 30558 6740 30564 6752
rect 30616 6740 30622 6792
rect 31036 6780 31156 6782
rect 31202 6780 31208 6792
rect 31036 6754 31208 6780
rect 24670 6672 24676 6724
rect 24728 6712 24734 6724
rect 24765 6715 24823 6721
rect 24765 6712 24777 6715
rect 24728 6684 24777 6712
rect 24728 6672 24734 6684
rect 24765 6681 24777 6684
rect 24811 6681 24823 6715
rect 25590 6712 25596 6724
rect 24765 6675 24823 6681
rect 24872 6684 25596 6712
rect 24578 6644 24584 6656
rect 22848 6616 24584 6644
rect 22741 6607 22799 6613
rect 24578 6604 24584 6616
rect 24636 6604 24642 6656
rect 24872 6653 24900 6684
rect 25590 6672 25596 6684
rect 25648 6672 25654 6724
rect 26688 6715 26746 6721
rect 26688 6681 26700 6715
rect 26734 6712 26746 6715
rect 27154 6712 27160 6724
rect 26734 6684 27160 6712
rect 26734 6681 26746 6684
rect 26688 6675 26746 6681
rect 27154 6672 27160 6684
rect 27212 6672 27218 6724
rect 31036 6712 31064 6754
rect 31128 6752 31208 6754
rect 31202 6740 31208 6752
rect 31260 6740 31266 6792
rect 31298 6783 31356 6789
rect 31298 6758 31310 6783
rect 31344 6758 31356 6783
rect 31390 6783 31448 6789
rect 27540 6684 31064 6712
rect 31294 6706 31300 6758
rect 31352 6706 31358 6758
rect 31390 6749 31402 6783
rect 31436 6780 31448 6783
rect 32858 6780 32864 6792
rect 31436 6752 31524 6780
rect 32819 6752 32864 6780
rect 31436 6749 31448 6752
rect 31390 6743 31448 6749
rect 31496 6712 31524 6752
rect 32858 6740 32864 6752
rect 32916 6740 32922 6792
rect 35618 6780 35624 6792
rect 35579 6752 35624 6780
rect 35618 6740 35624 6752
rect 35676 6740 35682 6792
rect 38105 6783 38163 6789
rect 38105 6780 38117 6783
rect 36924 6752 38117 6780
rect 31570 6712 31576 6724
rect 31496 6684 31576 6712
rect 24857 6647 24915 6653
rect 24857 6613 24869 6647
rect 24903 6613 24915 6647
rect 24857 6607 24915 6613
rect 24946 6604 24952 6656
rect 25004 6644 25010 6656
rect 25004 6616 25049 6644
rect 25004 6604 25010 6616
rect 25130 6604 25136 6656
rect 25188 6644 25194 6656
rect 27540 6644 27568 6684
rect 31570 6672 31576 6684
rect 31628 6672 31634 6724
rect 33962 6712 33968 6724
rect 33923 6684 33968 6712
rect 33962 6672 33968 6684
rect 34020 6672 34026 6724
rect 34149 6715 34207 6721
rect 34149 6681 34161 6715
rect 34195 6681 34207 6715
rect 34149 6675 34207 6681
rect 25188 6616 27568 6644
rect 25188 6604 25194 6616
rect 27614 6604 27620 6656
rect 27672 6644 27678 6656
rect 27801 6647 27859 6653
rect 27801 6644 27813 6647
rect 27672 6616 27813 6644
rect 27672 6604 27678 6616
rect 27801 6613 27813 6616
rect 27847 6613 27859 6647
rect 27801 6607 27859 6613
rect 28353 6647 28411 6653
rect 28353 6613 28365 6647
rect 28399 6644 28411 6647
rect 28902 6644 28908 6656
rect 28399 6616 28908 6644
rect 28399 6613 28411 6616
rect 28353 6607 28411 6613
rect 28902 6604 28908 6616
rect 28960 6604 28966 6656
rect 31021 6647 31079 6653
rect 31021 6613 31033 6647
rect 31067 6644 31079 6647
rect 31754 6644 31760 6656
rect 31067 6616 31760 6644
rect 31067 6613 31079 6616
rect 31021 6607 31079 6613
rect 31754 6604 31760 6616
rect 31812 6604 31818 6656
rect 33042 6644 33048 6656
rect 33003 6616 33048 6644
rect 33042 6604 33048 6616
rect 33100 6604 33106 6656
rect 34164 6644 34192 6675
rect 34606 6672 34612 6724
rect 34664 6712 34670 6724
rect 35437 6715 35495 6721
rect 35437 6712 35449 6715
rect 34664 6684 35449 6712
rect 34664 6672 34670 6684
rect 35437 6681 35449 6684
rect 35483 6681 35495 6715
rect 35437 6675 35495 6681
rect 34698 6644 34704 6656
rect 34164 6616 34704 6644
rect 34698 6604 34704 6616
rect 34756 6604 34762 6656
rect 36538 6644 36544 6656
rect 36499 6616 36544 6644
rect 36538 6604 36544 6616
rect 36596 6604 36602 6656
rect 36814 6604 36820 6656
rect 36872 6644 36878 6656
rect 36924 6653 36952 6752
rect 38105 6749 38117 6752
rect 38151 6749 38163 6783
rect 38105 6743 38163 6749
rect 38197 6783 38255 6789
rect 38197 6749 38209 6783
rect 38243 6749 38255 6783
rect 38197 6743 38255 6749
rect 37642 6672 37648 6724
rect 37700 6712 37706 6724
rect 38212 6712 38240 6743
rect 38286 6740 38292 6792
rect 38344 6780 38350 6792
rect 38488 6789 38516 6820
rect 39022 6808 39028 6820
rect 39080 6808 39086 6860
rect 38473 6783 38531 6789
rect 38344 6752 38389 6780
rect 38344 6740 38350 6752
rect 38473 6749 38485 6783
rect 38519 6749 38531 6783
rect 38473 6743 38531 6749
rect 38746 6740 38752 6792
rect 38804 6780 38810 6792
rect 38933 6783 38991 6789
rect 38933 6780 38945 6783
rect 38804 6752 38945 6780
rect 38804 6740 38810 6752
rect 38933 6749 38945 6752
rect 38979 6749 38991 6783
rect 38933 6743 38991 6749
rect 39117 6783 39175 6789
rect 39117 6749 39129 6783
rect 39163 6749 39175 6783
rect 39117 6743 39175 6749
rect 37700 6684 38240 6712
rect 37700 6672 37706 6684
rect 36909 6647 36967 6653
rect 36909 6644 36921 6647
rect 36872 6616 36921 6644
rect 36872 6604 36878 6616
rect 36909 6613 36921 6616
rect 36955 6613 36967 6647
rect 36909 6607 36967 6613
rect 36998 6604 37004 6656
rect 37056 6644 37062 6656
rect 37056 6616 37101 6644
rect 37056 6604 37062 6616
rect 38470 6604 38476 6656
rect 38528 6644 38534 6656
rect 39132 6644 39160 6743
rect 56686 6740 56692 6792
rect 56744 6780 56750 6792
rect 56873 6783 56931 6789
rect 56873 6780 56885 6783
rect 56744 6752 56885 6780
rect 56744 6740 56750 6752
rect 56873 6749 56885 6752
rect 56919 6749 56931 6783
rect 56873 6743 56931 6749
rect 57140 6783 57198 6789
rect 57140 6749 57152 6783
rect 57186 6780 57198 6783
rect 57514 6780 57520 6792
rect 57186 6752 57520 6780
rect 57186 6749 57198 6752
rect 57140 6743 57198 6749
rect 57514 6740 57520 6752
rect 57572 6740 57578 6792
rect 38528 6616 39160 6644
rect 38528 6604 38534 6616
rect 57514 6604 57520 6656
rect 57572 6644 57578 6656
rect 58253 6647 58311 6653
rect 58253 6644 58265 6647
rect 57572 6616 58265 6644
rect 57572 6604 57578 6616
rect 58253 6613 58265 6616
rect 58299 6613 58311 6647
rect 58253 6607 58311 6613
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11514 6440 11520 6452
rect 11195 6412 11520 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 12161 6443 12219 6449
rect 12161 6409 12173 6443
rect 12207 6440 12219 6443
rect 12250 6440 12256 6452
rect 12207 6412 12256 6440
rect 12207 6409 12219 6412
rect 12161 6403 12219 6409
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 16301 6443 16359 6449
rect 16301 6409 16313 6443
rect 16347 6440 16359 6443
rect 17770 6440 17776 6452
rect 16347 6412 17776 6440
rect 16347 6409 16359 6412
rect 16301 6403 16359 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 19518 6440 19524 6452
rect 17920 6412 17965 6440
rect 18985 6412 19524 6440
rect 17920 6400 17926 6412
rect 11606 6372 11612 6384
rect 2746 6344 11612 6372
rect 1581 6307 1639 6313
rect 1581 6273 1593 6307
rect 1627 6304 1639 6307
rect 2746 6304 2774 6344
rect 11606 6332 11612 6344
rect 11664 6332 11670 6384
rect 13262 6332 13268 6384
rect 13320 6372 13326 6384
rect 13633 6375 13691 6381
rect 13633 6372 13645 6375
rect 13320 6344 13645 6372
rect 13320 6332 13326 6344
rect 13633 6341 13645 6344
rect 13679 6341 13691 6375
rect 18230 6372 18236 6384
rect 18191 6344 18236 6372
rect 13633 6335 13691 6341
rect 18230 6332 18236 6344
rect 18288 6332 18294 6384
rect 18506 6332 18512 6384
rect 18564 6332 18570 6384
rect 1627 6276 2774 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 16942 6304 16948 6316
rect 9548 6276 16948 6304
rect 9548 6264 9554 6276
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 18524 6304 18552 6332
rect 18985 6304 19013 6412
rect 19518 6400 19524 6412
rect 19576 6400 19582 6452
rect 20070 6400 20076 6452
rect 20128 6440 20134 6452
rect 20441 6443 20499 6449
rect 20441 6440 20453 6443
rect 20128 6412 20453 6440
rect 20128 6400 20134 6412
rect 20441 6409 20453 6412
rect 20487 6409 20499 6443
rect 20441 6403 20499 6409
rect 23845 6443 23903 6449
rect 23845 6409 23857 6443
rect 23891 6440 23903 6443
rect 23934 6440 23940 6452
rect 23891 6412 23940 6440
rect 23891 6409 23903 6412
rect 23845 6403 23903 6409
rect 23934 6400 23940 6412
rect 23992 6440 23998 6452
rect 24762 6440 24768 6452
rect 23992 6412 24768 6440
rect 23992 6400 23998 6412
rect 24762 6400 24768 6412
rect 24820 6400 24826 6452
rect 24946 6440 24952 6452
rect 24859 6412 24952 6440
rect 24946 6400 24952 6412
rect 25004 6440 25010 6452
rect 25314 6440 25320 6452
rect 25004 6412 25320 6440
rect 25004 6400 25010 6412
rect 25314 6400 25320 6412
rect 25372 6400 25378 6452
rect 25774 6440 25780 6452
rect 25735 6412 25780 6440
rect 25774 6400 25780 6412
rect 25832 6400 25838 6452
rect 26142 6400 26148 6452
rect 26200 6440 26206 6452
rect 26237 6443 26295 6449
rect 26237 6440 26249 6443
rect 26200 6412 26249 6440
rect 26200 6400 26206 6412
rect 26237 6409 26249 6412
rect 26283 6409 26295 6443
rect 27154 6440 27160 6452
rect 27115 6412 27160 6440
rect 26237 6403 26295 6409
rect 27154 6400 27160 6412
rect 27212 6400 27218 6452
rect 27525 6443 27583 6449
rect 27525 6409 27537 6443
rect 27571 6440 27583 6443
rect 28258 6440 28264 6452
rect 27571 6412 28264 6440
rect 27571 6409 27583 6412
rect 27525 6403 27583 6409
rect 28258 6400 28264 6412
rect 28316 6400 28322 6452
rect 28994 6440 29000 6452
rect 28368 6412 29000 6440
rect 19242 6332 19248 6384
rect 19300 6381 19306 6384
rect 19300 6375 19364 6381
rect 19300 6341 19318 6375
rect 19352 6341 19364 6375
rect 19300 6335 19364 6341
rect 19300 6332 19306 6335
rect 19978 6332 19984 6384
rect 20036 6372 20042 6384
rect 24029 6375 24087 6381
rect 24029 6372 24041 6375
rect 20036 6344 24041 6372
rect 20036 6332 20042 6344
rect 24029 6341 24041 6344
rect 24075 6341 24087 6375
rect 25038 6372 25044 6384
rect 24029 6335 24087 6341
rect 24780 6344 25044 6372
rect 19061 6307 19119 6313
rect 19061 6304 19073 6307
rect 17926 6276 18920 6304
rect 18985 6276 19073 6304
rect 1762 6236 1768 6248
rect 1723 6208 1768 6236
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6236 10747 6239
rect 11054 6236 11060 6248
rect 10735 6208 11060 6236
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 11054 6196 11060 6208
rect 11112 6236 11118 6248
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 11112 6208 11713 6236
rect 11112 6196 11118 6208
rect 11701 6205 11713 6208
rect 11747 6236 11759 6239
rect 12342 6236 12348 6248
rect 11747 6208 12348 6236
rect 11747 6205 11759 6208
rect 11701 6199 11759 6205
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 15562 6236 15568 6248
rect 13924 6208 15568 6236
rect 8846 6128 8852 6180
rect 8904 6168 8910 6180
rect 10965 6171 11023 6177
rect 10965 6168 10977 6171
rect 8904 6140 10977 6168
rect 8904 6128 8910 6140
rect 10965 6137 10977 6140
rect 11011 6137 11023 6171
rect 10965 6131 11023 6137
rect 11514 6128 11520 6180
rect 11572 6168 11578 6180
rect 11977 6171 12035 6177
rect 11977 6168 11989 6171
rect 11572 6140 11989 6168
rect 11572 6128 11578 6140
rect 11977 6137 11989 6140
rect 12023 6137 12035 6171
rect 11977 6131 12035 6137
rect 10134 6060 10140 6112
rect 10192 6100 10198 6112
rect 13924 6100 13952 6208
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 15654 6196 15660 6248
rect 15712 6236 15718 6248
rect 15841 6239 15899 6245
rect 15841 6236 15853 6239
rect 15712 6208 15853 6236
rect 15712 6196 15718 6208
rect 15841 6205 15853 6208
rect 15887 6236 15899 6239
rect 17926 6236 17954 6276
rect 18322 6236 18328 6248
rect 15887 6208 17954 6236
rect 18283 6208 18328 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 18509 6239 18567 6245
rect 18509 6205 18521 6239
rect 18555 6236 18567 6239
rect 18598 6236 18604 6248
rect 18555 6208 18604 6236
rect 18555 6205 18567 6208
rect 18509 6199 18567 6205
rect 18598 6196 18604 6208
rect 18656 6196 18662 6248
rect 14001 6171 14059 6177
rect 14001 6137 14013 6171
rect 14047 6168 14059 6171
rect 14550 6168 14556 6180
rect 14047 6140 14556 6168
rect 14047 6137 14059 6140
rect 14001 6131 14059 6137
rect 14550 6128 14556 6140
rect 14608 6128 14614 6180
rect 16114 6168 16120 6180
rect 16075 6140 16120 6168
rect 16114 6128 16120 6140
rect 16172 6128 16178 6180
rect 18892 6168 18920 6276
rect 19061 6273 19073 6276
rect 19107 6273 19119 6307
rect 19061 6267 19119 6273
rect 19150 6264 19156 6316
rect 19208 6304 19214 6316
rect 21634 6304 21640 6316
rect 19208 6276 21640 6304
rect 19208 6264 19214 6276
rect 21634 6264 21640 6276
rect 21692 6264 21698 6316
rect 22557 6307 22615 6313
rect 22557 6273 22569 6307
rect 22603 6304 22615 6307
rect 22922 6304 22928 6316
rect 22603 6276 22928 6304
rect 22603 6273 22615 6276
rect 22557 6267 22615 6273
rect 22922 6264 22928 6276
rect 22980 6264 22986 6316
rect 23658 6304 23664 6316
rect 23619 6276 23664 6304
rect 23658 6264 23664 6276
rect 23716 6264 23722 6316
rect 23799 6307 23857 6313
rect 23799 6273 23811 6307
rect 23845 6304 23857 6307
rect 24780 6304 24808 6344
rect 25038 6332 25044 6344
rect 25096 6332 25102 6384
rect 25590 6332 25596 6384
rect 25648 6372 25654 6384
rect 28368 6372 28396 6412
rect 28994 6400 29000 6412
rect 29052 6400 29058 6452
rect 30006 6440 30012 6452
rect 29967 6412 30012 6440
rect 30006 6400 30012 6412
rect 30064 6400 30070 6452
rect 31846 6400 31852 6452
rect 31904 6440 31910 6452
rect 57517 6443 57575 6449
rect 31904 6412 36676 6440
rect 31904 6400 31910 6412
rect 33042 6381 33048 6384
rect 25648 6344 28396 6372
rect 30852 6344 32996 6372
rect 25648 6332 25654 6344
rect 23845 6276 24808 6304
rect 23845 6273 23857 6276
rect 23799 6267 23857 6273
rect 24854 6264 24860 6316
rect 24912 6304 24918 6316
rect 25498 6304 25504 6316
rect 24912 6276 25504 6304
rect 24912 6264 24918 6276
rect 25498 6264 25504 6276
rect 25556 6264 25562 6316
rect 26050 6264 26056 6316
rect 26108 6304 26114 6316
rect 26145 6307 26203 6313
rect 26145 6304 26157 6307
rect 26108 6276 26157 6304
rect 26108 6264 26114 6276
rect 26145 6273 26157 6276
rect 26191 6273 26203 6307
rect 26145 6267 26203 6273
rect 27522 6264 27528 6316
rect 27580 6304 27586 6316
rect 27580 6276 27752 6304
rect 27580 6264 27586 6276
rect 22741 6239 22799 6245
rect 22741 6205 22753 6239
rect 22787 6205 22799 6239
rect 22741 6199 22799 6205
rect 19058 6168 19064 6180
rect 16224 6140 18092 6168
rect 18892 6140 19064 6168
rect 10192 6072 13952 6100
rect 14093 6103 14151 6109
rect 10192 6060 10198 6072
rect 14093 6069 14105 6103
rect 14139 6100 14151 6103
rect 16224 6100 16252 6140
rect 14139 6072 16252 6100
rect 18064 6100 18092 6140
rect 19058 6128 19064 6140
rect 19116 6128 19122 6180
rect 22554 6128 22560 6180
rect 22612 6168 22618 6180
rect 22756 6168 22784 6199
rect 22830 6196 22836 6248
rect 22888 6236 22894 6248
rect 25133 6239 25191 6245
rect 22888 6208 24992 6236
rect 22888 6196 22894 6208
rect 22612 6140 22784 6168
rect 23477 6171 23535 6177
rect 22612 6128 22618 6140
rect 23477 6137 23489 6171
rect 23523 6168 23535 6171
rect 23842 6168 23848 6180
rect 23523 6140 23848 6168
rect 23523 6137 23535 6140
rect 23477 6131 23535 6137
rect 23842 6128 23848 6140
rect 23900 6128 23906 6180
rect 24964 6168 24992 6208
rect 25133 6205 25145 6239
rect 25179 6236 25191 6239
rect 25682 6236 25688 6248
rect 25179 6208 25688 6236
rect 25179 6205 25191 6208
rect 25133 6199 25191 6205
rect 25682 6196 25688 6208
rect 25740 6236 25746 6248
rect 25958 6236 25964 6248
rect 25740 6208 25964 6236
rect 25740 6196 25746 6208
rect 25958 6196 25964 6208
rect 26016 6196 26022 6248
rect 26418 6236 26424 6248
rect 26379 6208 26424 6236
rect 26418 6196 26424 6208
rect 26476 6196 26482 6248
rect 27614 6236 27620 6248
rect 27527 6208 27620 6236
rect 27614 6196 27620 6208
rect 27672 6196 27678 6248
rect 27724 6245 27752 6276
rect 28074 6264 28080 6316
rect 28132 6304 28138 6316
rect 30852 6313 30880 6344
rect 28629 6307 28687 6313
rect 28629 6304 28641 6307
rect 28132 6276 28641 6304
rect 28132 6264 28138 6276
rect 28629 6273 28641 6276
rect 28675 6304 28687 6307
rect 30837 6307 30895 6313
rect 28675 6276 30420 6304
rect 28675 6273 28687 6276
rect 28629 6267 28687 6273
rect 27709 6239 27767 6245
rect 27709 6205 27721 6239
rect 27755 6205 27767 6239
rect 28902 6236 28908 6248
rect 28863 6208 28908 6236
rect 27709 6199 27767 6205
rect 28902 6196 28908 6208
rect 28960 6196 28966 6248
rect 30392 6236 30420 6276
rect 30837 6273 30849 6307
rect 30883 6273 30895 6307
rect 30837 6267 30895 6273
rect 31113 6307 31171 6313
rect 31113 6273 31125 6307
rect 31159 6304 31171 6307
rect 31202 6304 31208 6316
rect 31159 6276 31208 6304
rect 31159 6273 31171 6276
rect 31113 6267 31171 6273
rect 31202 6264 31208 6276
rect 31260 6304 31266 6316
rect 31938 6304 31944 6316
rect 31260 6276 31944 6304
rect 31260 6264 31266 6276
rect 31938 6264 31944 6276
rect 31996 6264 32002 6316
rect 32674 6264 32680 6316
rect 32732 6304 32738 6316
rect 32769 6307 32827 6313
rect 32769 6304 32781 6307
rect 32732 6276 32781 6304
rect 32732 6264 32738 6276
rect 32769 6273 32781 6276
rect 32815 6273 32827 6307
rect 32968 6304 32996 6344
rect 33036 6335 33048 6381
rect 33100 6372 33106 6384
rect 33100 6344 33136 6372
rect 33042 6332 33048 6335
rect 33100 6332 33106 6344
rect 35618 6332 35624 6384
rect 35676 6372 35682 6384
rect 35802 6372 35808 6384
rect 35676 6344 35808 6372
rect 35676 6332 35682 6344
rect 35802 6332 35808 6344
rect 35860 6332 35866 6384
rect 36648 6381 36676 6412
rect 57517 6409 57529 6443
rect 57563 6440 57575 6443
rect 57606 6440 57612 6452
rect 57563 6412 57612 6440
rect 57563 6409 57575 6412
rect 57517 6403 57575 6409
rect 57606 6400 57612 6412
rect 57664 6400 57670 6452
rect 36633 6375 36691 6381
rect 36633 6341 36645 6375
rect 36679 6341 36691 6375
rect 36633 6335 36691 6341
rect 34790 6304 34796 6316
rect 32968 6276 34796 6304
rect 32769 6267 32827 6273
rect 34790 6264 34796 6276
rect 34848 6264 34854 6316
rect 36265 6307 36323 6313
rect 36265 6273 36277 6307
rect 36311 6273 36323 6307
rect 36648 6304 36676 6335
rect 37366 6332 37372 6384
rect 37424 6372 37430 6384
rect 37737 6375 37795 6381
rect 37737 6372 37749 6375
rect 37424 6344 37749 6372
rect 37424 6332 37430 6344
rect 37737 6341 37749 6344
rect 37783 6341 37795 6375
rect 37737 6335 37795 6341
rect 37461 6307 37519 6313
rect 37461 6304 37473 6307
rect 36648 6276 37473 6304
rect 36265 6267 36323 6273
rect 37461 6273 37473 6276
rect 37507 6273 37519 6307
rect 37461 6267 37519 6273
rect 30926 6236 30932 6248
rect 30392 6208 30932 6236
rect 30926 6196 30932 6208
rect 30984 6236 30990 6248
rect 32692 6236 32720 6264
rect 30984 6208 32720 6236
rect 36280 6236 36308 6267
rect 57238 6264 57244 6316
rect 57296 6304 57302 6316
rect 57333 6307 57391 6313
rect 57333 6304 57345 6307
rect 57296 6276 57345 6304
rect 57296 6264 57302 6276
rect 57333 6273 57345 6276
rect 57379 6273 57391 6307
rect 57514 6304 57520 6316
rect 57475 6276 57520 6304
rect 57333 6267 57391 6273
rect 57514 6264 57520 6276
rect 57572 6264 57578 6316
rect 38562 6236 38568 6248
rect 36280 6208 38568 6236
rect 30984 6196 30990 6208
rect 38562 6196 38568 6208
rect 38620 6196 38626 6248
rect 27632 6168 27660 6196
rect 24964 6140 27660 6168
rect 30098 6128 30104 6180
rect 30156 6168 30162 6180
rect 31113 6171 31171 6177
rect 31113 6168 31125 6171
rect 30156 6140 31125 6168
rect 30156 6128 30162 6140
rect 31113 6137 31125 6140
rect 31159 6168 31171 6171
rect 31294 6168 31300 6180
rect 31159 6140 31300 6168
rect 31159 6137 31171 6140
rect 31113 6131 31171 6137
rect 31294 6128 31300 6140
rect 31352 6128 31358 6180
rect 33778 6128 33784 6180
rect 33836 6168 33842 6180
rect 37182 6168 37188 6180
rect 33836 6140 37188 6168
rect 33836 6128 33842 6140
rect 37182 6128 37188 6140
rect 37240 6128 37246 6180
rect 24026 6100 24032 6112
rect 18064 6072 24032 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 24026 6060 24032 6072
rect 24084 6060 24090 6112
rect 24486 6100 24492 6112
rect 24447 6072 24492 6100
rect 24486 6060 24492 6072
rect 24544 6060 24550 6112
rect 24578 6060 24584 6112
rect 24636 6100 24642 6112
rect 33134 6100 33140 6112
rect 24636 6072 33140 6100
rect 24636 6060 24642 6072
rect 33134 6060 33140 6072
rect 33192 6060 33198 6112
rect 33410 6060 33416 6112
rect 33468 6100 33474 6112
rect 34149 6103 34207 6109
rect 34149 6100 34161 6103
rect 33468 6072 34161 6100
rect 33468 6060 33474 6072
rect 34149 6069 34161 6072
rect 34195 6069 34207 6103
rect 34149 6063 34207 6069
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 11977 5899 12035 5905
rect 11977 5865 11989 5899
rect 12023 5896 12035 5899
rect 13078 5896 13084 5908
rect 12023 5868 13084 5896
rect 12023 5865 12035 5868
rect 11977 5859 12035 5865
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 13633 5899 13691 5905
rect 13633 5865 13645 5899
rect 13679 5896 13691 5899
rect 16114 5896 16120 5908
rect 13679 5868 16120 5896
rect 13679 5865 13691 5868
rect 13633 5859 13691 5865
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 22830 5896 22836 5908
rect 16224 5868 22836 5896
rect 12897 5831 12955 5837
rect 12897 5797 12909 5831
rect 12943 5828 12955 5831
rect 12986 5828 12992 5840
rect 12943 5800 12992 5828
rect 12943 5797 12955 5800
rect 12897 5791 12955 5797
rect 12986 5788 12992 5800
rect 13044 5788 13050 5840
rect 13538 5788 13544 5840
rect 13596 5828 13602 5840
rect 16224 5828 16252 5868
rect 22830 5856 22836 5868
rect 22888 5856 22894 5908
rect 26326 5856 26332 5908
rect 26384 5896 26390 5908
rect 31110 5896 31116 5908
rect 26384 5868 31116 5896
rect 26384 5856 26390 5868
rect 31110 5856 31116 5868
rect 31168 5856 31174 5908
rect 32858 5896 32864 5908
rect 32819 5868 32864 5896
rect 32858 5856 32864 5868
rect 32916 5856 32922 5908
rect 36814 5896 36820 5908
rect 33244 5868 36820 5896
rect 13596 5800 16252 5828
rect 18141 5831 18199 5837
rect 13596 5788 13602 5800
rect 18141 5797 18153 5831
rect 18187 5828 18199 5831
rect 18966 5828 18972 5840
rect 18187 5800 18972 5828
rect 18187 5797 18199 5800
rect 18141 5791 18199 5797
rect 18966 5788 18972 5800
rect 19024 5788 19030 5840
rect 23477 5831 23535 5837
rect 23477 5797 23489 5831
rect 23523 5828 23535 5831
rect 23566 5828 23572 5840
rect 23523 5800 23572 5828
rect 23523 5797 23535 5800
rect 23477 5791 23535 5797
rect 23566 5788 23572 5800
rect 23624 5788 23630 5840
rect 23658 5788 23664 5840
rect 23716 5828 23722 5840
rect 23716 5800 24716 5828
rect 23716 5788 23722 5800
rect 24688 5772 24716 5800
rect 28166 5788 28172 5840
rect 28224 5788 28230 5840
rect 28994 5788 29000 5840
rect 29052 5828 29058 5840
rect 33244 5828 33272 5868
rect 36814 5856 36820 5868
rect 36872 5896 36878 5908
rect 37829 5899 37887 5905
rect 37829 5896 37841 5899
rect 36872 5868 37841 5896
rect 36872 5856 36878 5868
rect 37829 5865 37841 5868
rect 37875 5865 37887 5899
rect 37829 5859 37887 5865
rect 34606 5828 34612 5840
rect 29052 5800 33272 5828
rect 33336 5800 34612 5828
rect 29052 5788 29058 5800
rect 18598 5720 18604 5772
rect 18656 5760 18662 5772
rect 18693 5763 18751 5769
rect 18693 5760 18705 5763
rect 18656 5732 18705 5760
rect 18656 5720 18662 5732
rect 18693 5729 18705 5732
rect 18739 5729 18751 5763
rect 19426 5760 19432 5772
rect 19387 5732 19432 5760
rect 18693 5723 18751 5729
rect 19426 5720 19432 5732
rect 19484 5720 19490 5772
rect 22002 5760 22008 5772
rect 21376 5732 22008 5760
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5692 17739 5695
rect 17770 5692 17776 5704
rect 17727 5664 17776 5692
rect 17727 5661 17739 5664
rect 17681 5655 17739 5661
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 21376 5692 21404 5732
rect 22002 5720 22008 5732
rect 22060 5720 22066 5772
rect 22462 5760 22468 5772
rect 22423 5732 22468 5760
rect 22462 5720 22468 5732
rect 22520 5720 22526 5772
rect 24670 5720 24676 5772
rect 24728 5760 24734 5772
rect 25590 5760 25596 5772
rect 24728 5732 25360 5760
rect 25551 5732 25596 5760
rect 24728 5720 24734 5732
rect 17972 5664 21404 5692
rect 21453 5695 21511 5701
rect 11698 5584 11704 5636
rect 11756 5624 11762 5636
rect 11885 5627 11943 5633
rect 11885 5624 11897 5627
rect 11756 5596 11897 5624
rect 11756 5584 11762 5596
rect 11885 5593 11897 5596
rect 11931 5593 11943 5627
rect 11885 5587 11943 5593
rect 12526 5584 12532 5636
rect 12584 5624 12590 5636
rect 12713 5627 12771 5633
rect 12713 5624 12725 5627
rect 12584 5596 12725 5624
rect 12584 5584 12590 5596
rect 12713 5593 12725 5596
rect 12759 5593 12771 5627
rect 12713 5587 12771 5593
rect 13354 5584 13360 5636
rect 13412 5624 13418 5636
rect 13541 5627 13599 5633
rect 13541 5624 13553 5627
rect 13412 5596 13553 5624
rect 13412 5584 13418 5596
rect 13541 5593 13553 5596
rect 13587 5593 13599 5627
rect 13541 5587 13599 5593
rect 14182 5584 14188 5636
rect 14240 5624 14246 5636
rect 14369 5627 14427 5633
rect 14369 5624 14381 5627
rect 14240 5596 14381 5624
rect 14240 5584 14246 5596
rect 14369 5593 14381 5596
rect 14415 5593 14427 5627
rect 14369 5587 14427 5593
rect 16574 5584 16580 5636
rect 16632 5624 16638 5636
rect 17972 5624 18000 5664
rect 21453 5661 21465 5695
rect 21499 5692 21511 5695
rect 22278 5692 22284 5704
rect 21499 5664 22284 5692
rect 21499 5661 21511 5664
rect 21453 5655 21511 5661
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 22646 5692 22652 5704
rect 22559 5664 22652 5692
rect 22646 5652 22652 5664
rect 22704 5692 22710 5704
rect 23799 5695 23857 5701
rect 22704 5664 23704 5692
rect 22704 5652 22710 5664
rect 23676 5636 23704 5664
rect 23799 5661 23811 5695
rect 23845 5661 23857 5695
rect 24026 5692 24032 5704
rect 23987 5664 24032 5692
rect 23799 5655 23857 5661
rect 16632 5596 18000 5624
rect 16632 5584 16638 5596
rect 18966 5584 18972 5636
rect 19024 5624 19030 5636
rect 19674 5627 19732 5633
rect 19674 5624 19686 5627
rect 19024 5596 19686 5624
rect 19024 5584 19030 5596
rect 19674 5593 19686 5596
rect 19720 5593 19732 5627
rect 19674 5587 19732 5593
rect 21358 5584 21364 5636
rect 21416 5624 21422 5636
rect 21729 5627 21787 5633
rect 21729 5624 21741 5627
rect 21416 5596 21741 5624
rect 21416 5584 21422 5596
rect 21729 5593 21741 5596
rect 21775 5593 21787 5627
rect 21729 5587 21787 5593
rect 21818 5584 21824 5636
rect 21876 5624 21882 5636
rect 22370 5624 22376 5636
rect 21876 5596 22376 5624
rect 21876 5584 21882 5596
rect 22370 5584 22376 5596
rect 22428 5624 22434 5636
rect 23014 5624 23020 5636
rect 22428 5596 22876 5624
rect 22975 5596 23020 5624
rect 22428 5584 22434 5596
rect 14458 5556 14464 5568
rect 14419 5528 14464 5556
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 17126 5516 17132 5568
rect 17184 5556 17190 5568
rect 18506 5556 18512 5568
rect 17184 5528 18512 5556
rect 17184 5516 17190 5528
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 18598 5516 18604 5568
rect 18656 5556 18662 5568
rect 18656 5528 18701 5556
rect 18656 5516 18662 5528
rect 18874 5516 18880 5568
rect 18932 5556 18938 5568
rect 20254 5556 20260 5568
rect 18932 5528 20260 5556
rect 18932 5516 18938 5528
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 20806 5556 20812 5568
rect 20767 5528 20812 5556
rect 20806 5516 20812 5528
rect 20864 5516 20870 5568
rect 22738 5556 22744 5568
rect 22699 5528 22744 5556
rect 22738 5516 22744 5528
rect 22796 5516 22802 5568
rect 22848 5565 22876 5596
rect 23014 5584 23020 5596
rect 23072 5584 23078 5636
rect 23658 5624 23664 5636
rect 23619 5596 23664 5624
rect 23658 5584 23664 5596
rect 23716 5584 23722 5636
rect 23814 5624 23842 5655
rect 24026 5652 24032 5664
rect 24084 5652 24090 5704
rect 24394 5624 24400 5636
rect 23814 5596 24400 5624
rect 24394 5584 24400 5596
rect 24452 5584 24458 5636
rect 24578 5624 24584 5636
rect 24539 5596 24584 5624
rect 24578 5584 24584 5596
rect 24636 5584 24642 5636
rect 24780 5633 24808 5732
rect 24903 5695 24961 5701
rect 24903 5661 24915 5695
rect 24949 5692 24961 5695
rect 25222 5692 25228 5704
rect 24949 5664 25228 5692
rect 24949 5661 24961 5664
rect 24903 5655 24961 5661
rect 25222 5652 25228 5664
rect 25280 5652 25286 5704
rect 25332 5692 25360 5732
rect 25590 5720 25596 5732
rect 25648 5720 25654 5772
rect 28184 5760 28212 5788
rect 28184 5732 28301 5760
rect 25774 5692 25780 5704
rect 25332 5664 25780 5692
rect 25774 5652 25780 5664
rect 25832 5652 25838 5704
rect 25958 5652 25964 5704
rect 26016 5692 26022 5704
rect 26145 5695 26203 5701
rect 26145 5692 26157 5695
rect 26016 5664 26157 5692
rect 26016 5652 26022 5664
rect 26145 5661 26157 5664
rect 26191 5661 26203 5695
rect 26145 5655 26203 5661
rect 27614 5652 27620 5704
rect 27672 5692 27678 5704
rect 28149 5695 28207 5701
rect 28273 5698 28301 5732
rect 28626 5720 28632 5772
rect 28684 5760 28690 5772
rect 33336 5760 33364 5800
rect 34606 5788 34612 5800
rect 34664 5788 34670 5840
rect 28684 5732 33364 5760
rect 33505 5763 33563 5769
rect 28684 5720 28690 5732
rect 33505 5729 33517 5763
rect 33551 5760 33563 5763
rect 33778 5760 33784 5772
rect 33551 5732 33784 5760
rect 33551 5729 33563 5732
rect 33505 5723 33563 5729
rect 33778 5720 33784 5732
rect 33836 5720 33842 5772
rect 34514 5720 34520 5772
rect 34572 5760 34578 5772
rect 35342 5760 35348 5772
rect 34572 5732 35348 5760
rect 34572 5720 34578 5732
rect 35342 5720 35348 5732
rect 35400 5760 35406 5772
rect 36449 5763 36507 5769
rect 36449 5760 36461 5763
rect 35400 5732 36461 5760
rect 35400 5720 35406 5732
rect 36449 5729 36461 5732
rect 36495 5729 36507 5763
rect 36449 5723 36507 5729
rect 28149 5692 28161 5695
rect 27672 5664 28161 5692
rect 27672 5652 27678 5664
rect 28149 5661 28161 5664
rect 28195 5661 28207 5695
rect 28149 5655 28207 5661
rect 28258 5692 28316 5698
rect 28258 5658 28270 5692
rect 28304 5658 28316 5692
rect 28258 5652 28316 5658
rect 28350 5652 28356 5704
rect 28408 5701 28414 5704
rect 28408 5692 28416 5701
rect 28537 5695 28595 5701
rect 28408 5664 28453 5692
rect 28408 5655 28416 5664
rect 28537 5661 28549 5695
rect 28583 5692 28595 5695
rect 30282 5692 30288 5704
rect 28583 5664 30288 5692
rect 28583 5661 28595 5664
rect 28537 5655 28595 5661
rect 28408 5652 28414 5655
rect 30282 5652 30288 5664
rect 30340 5652 30346 5704
rect 30466 5692 30472 5704
rect 30427 5664 30472 5692
rect 30466 5652 30472 5664
rect 30524 5652 30530 5704
rect 31662 5652 31668 5704
rect 31720 5692 31726 5704
rect 32122 5692 32128 5704
rect 31720 5664 32128 5692
rect 31720 5652 31726 5664
rect 32122 5652 32128 5664
rect 32180 5652 32186 5704
rect 33226 5692 33232 5704
rect 33187 5664 33232 5692
rect 33226 5652 33232 5664
rect 33284 5652 33290 5704
rect 33321 5695 33379 5701
rect 33321 5661 33333 5695
rect 33367 5692 33379 5695
rect 56965 5695 57023 5701
rect 33367 5664 45554 5692
rect 33367 5661 33379 5664
rect 33321 5655 33379 5661
rect 24765 5627 24823 5633
rect 24765 5593 24777 5627
rect 24811 5593 24823 5627
rect 24765 5587 24823 5593
rect 25130 5584 25136 5636
rect 25188 5624 25194 5636
rect 25188 5596 25233 5624
rect 25415 5596 26004 5624
rect 25188 5584 25194 5596
rect 22833 5559 22891 5565
rect 22833 5525 22845 5559
rect 22879 5556 22891 5559
rect 23845 5559 23903 5565
rect 23845 5556 23857 5559
rect 22879 5528 23857 5556
rect 22879 5525 22891 5528
rect 22833 5519 22891 5525
rect 23845 5525 23857 5528
rect 23891 5556 23903 5559
rect 23934 5556 23940 5568
rect 23891 5528 23940 5556
rect 23891 5525 23903 5528
rect 23845 5519 23903 5525
rect 23934 5516 23940 5528
rect 23992 5556 23998 5568
rect 24949 5559 25007 5565
rect 24949 5556 24961 5559
rect 23992 5528 24961 5556
rect 23992 5516 23998 5528
rect 24949 5525 24961 5528
rect 24995 5556 25007 5559
rect 25415 5556 25443 5596
rect 25866 5556 25872 5568
rect 24995 5528 25443 5556
rect 25827 5528 25872 5556
rect 24995 5525 25007 5528
rect 24949 5519 25007 5525
rect 25866 5516 25872 5528
rect 25924 5516 25930 5568
rect 25976 5565 26004 5596
rect 28902 5584 28908 5636
rect 28960 5624 28966 5636
rect 33336 5624 33364 5655
rect 28960 5596 33364 5624
rect 28960 5584 28966 5596
rect 33410 5584 33416 5636
rect 33468 5624 33474 5636
rect 33594 5624 33600 5636
rect 33468 5596 33600 5624
rect 33468 5584 33474 5596
rect 33594 5584 33600 5596
rect 33652 5584 33658 5636
rect 34977 5627 35035 5633
rect 34977 5593 34989 5627
rect 35023 5624 35035 5627
rect 35526 5624 35532 5636
rect 35023 5596 35532 5624
rect 35023 5593 35035 5596
rect 34977 5587 35035 5593
rect 35526 5584 35532 5596
rect 35584 5624 35590 5636
rect 35713 5627 35771 5633
rect 35713 5624 35725 5627
rect 35584 5596 35725 5624
rect 35584 5584 35590 5596
rect 35713 5593 35725 5596
rect 35759 5593 35771 5627
rect 35894 5624 35900 5636
rect 35855 5596 35900 5624
rect 35713 5587 35771 5593
rect 35894 5584 35900 5596
rect 35952 5584 35958 5636
rect 36722 5633 36728 5636
rect 36716 5587 36728 5633
rect 36780 5624 36786 5636
rect 36780 5596 36816 5624
rect 36722 5584 36728 5587
rect 36780 5584 36786 5596
rect 25961 5559 26019 5565
rect 25961 5525 25973 5559
rect 26007 5525 26019 5559
rect 25961 5519 26019 5525
rect 27893 5559 27951 5565
rect 27893 5525 27905 5559
rect 27939 5556 27951 5559
rect 28350 5556 28356 5568
rect 27939 5528 28356 5556
rect 27939 5525 27951 5528
rect 27893 5519 27951 5525
rect 28350 5516 28356 5528
rect 28408 5516 28414 5568
rect 28810 5516 28816 5568
rect 28868 5556 28874 5568
rect 28997 5559 29055 5565
rect 28997 5556 29009 5559
rect 28868 5528 29009 5556
rect 28868 5516 28874 5528
rect 28997 5525 29009 5528
rect 29043 5525 29055 5559
rect 30650 5556 30656 5568
rect 30611 5528 30656 5556
rect 28997 5519 29055 5525
rect 30650 5516 30656 5528
rect 30708 5516 30714 5568
rect 32674 5516 32680 5568
rect 32732 5556 32738 5568
rect 34514 5556 34520 5568
rect 32732 5528 34520 5556
rect 32732 5516 32738 5528
rect 34514 5516 34520 5528
rect 34572 5516 34578 5568
rect 34790 5516 34796 5568
rect 34848 5556 34854 5568
rect 35069 5559 35127 5565
rect 35069 5556 35081 5559
rect 34848 5528 35081 5556
rect 34848 5516 34854 5528
rect 35069 5525 35081 5528
rect 35115 5525 35127 5559
rect 45526 5556 45554 5664
rect 56965 5661 56977 5695
rect 57011 5692 57023 5695
rect 57514 5692 57520 5704
rect 57011 5664 57520 5692
rect 57011 5661 57023 5664
rect 56965 5655 57023 5661
rect 57514 5652 57520 5664
rect 57572 5652 57578 5704
rect 57974 5692 57980 5704
rect 57935 5664 57980 5692
rect 57974 5652 57980 5664
rect 58032 5652 58038 5704
rect 57238 5624 57244 5636
rect 57199 5596 57244 5624
rect 57238 5584 57244 5596
rect 57296 5584 57302 5636
rect 58069 5559 58127 5565
rect 58069 5556 58081 5559
rect 45526 5528 58081 5556
rect 35069 5519 35127 5525
rect 58069 5525 58081 5528
rect 58115 5525 58127 5559
rect 58069 5519 58127 5525
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 12342 5352 12348 5364
rect 12303 5324 12348 5352
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 18322 5312 18328 5364
rect 18380 5352 18386 5364
rect 18417 5355 18475 5361
rect 18417 5352 18429 5355
rect 18380 5324 18429 5352
rect 18380 5312 18386 5324
rect 18417 5321 18429 5324
rect 18463 5321 18475 5355
rect 18417 5315 18475 5321
rect 18877 5355 18935 5361
rect 18877 5321 18889 5355
rect 18923 5352 18935 5355
rect 28994 5352 29000 5364
rect 18923 5324 29000 5352
rect 18923 5321 18935 5324
rect 18877 5315 18935 5321
rect 11146 5284 11152 5296
rect 11107 5256 11152 5284
rect 11146 5244 11152 5256
rect 11204 5244 11210 5296
rect 13814 5284 13820 5296
rect 13775 5256 13820 5284
rect 13814 5244 13820 5256
rect 13872 5244 13878 5296
rect 18141 5287 18199 5293
rect 18141 5253 18153 5287
rect 18187 5284 18199 5287
rect 18892 5284 18920 5315
rect 28994 5312 29000 5324
rect 29052 5312 29058 5364
rect 29454 5352 29460 5364
rect 29415 5324 29460 5352
rect 29454 5312 29460 5324
rect 29512 5312 29518 5364
rect 30377 5355 30435 5361
rect 30377 5321 30389 5355
rect 30423 5352 30435 5355
rect 30466 5352 30472 5364
rect 30423 5324 30472 5352
rect 30423 5321 30435 5324
rect 30377 5315 30435 5321
rect 30466 5312 30472 5324
rect 30524 5312 30530 5364
rect 31938 5312 31944 5364
rect 31996 5352 32002 5364
rect 32677 5355 32735 5361
rect 32677 5352 32689 5355
rect 31996 5324 32689 5352
rect 31996 5312 32002 5324
rect 32677 5321 32689 5324
rect 32723 5352 32735 5355
rect 32766 5352 32772 5364
rect 32723 5324 32772 5352
rect 32723 5321 32735 5324
rect 32677 5315 32735 5321
rect 32766 5312 32772 5324
rect 32824 5352 32830 5364
rect 33689 5355 33747 5361
rect 33689 5352 33701 5355
rect 32824 5324 33701 5352
rect 32824 5312 32830 5324
rect 33689 5321 33701 5324
rect 33735 5321 33747 5355
rect 33689 5315 33747 5321
rect 34054 5312 34060 5364
rect 34112 5352 34118 5364
rect 34698 5352 34704 5364
rect 34112 5324 34704 5352
rect 34112 5312 34118 5324
rect 34698 5312 34704 5324
rect 34756 5312 34762 5364
rect 35437 5355 35495 5361
rect 35437 5321 35449 5355
rect 35483 5321 35495 5355
rect 36722 5352 36728 5364
rect 36683 5324 36728 5352
rect 35437 5315 35495 5321
rect 19889 5287 19947 5293
rect 19889 5284 19901 5287
rect 18187 5256 18920 5284
rect 18984 5256 19901 5284
rect 18187 5253 18199 5256
rect 18141 5247 18199 5253
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5216 1639 5219
rect 9858 5216 9864 5228
rect 1627 5188 9864 5216
rect 1627 5185 1639 5188
rect 1581 5179 1639 5185
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 10100 5188 10241 5216
rect 10100 5176 10106 5188
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10962 5216 10968 5228
rect 10923 5188 10968 5216
rect 10229 5179 10287 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5216 12219 5219
rect 13630 5216 13636 5228
rect 12207 5188 12434 5216
rect 13591 5188 13636 5216
rect 12207 5185 12219 5188
rect 12161 5179 12219 5185
rect 1762 5148 1768 5160
rect 1723 5120 1768 5148
rect 1762 5108 1768 5120
rect 1820 5108 1826 5160
rect 7926 5108 7932 5160
rect 7984 5148 7990 5160
rect 12406 5148 12434 5188
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 17736 5188 18797 5216
rect 17736 5176 17742 5188
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 18984 5216 19012 5256
rect 19889 5253 19901 5256
rect 19935 5253 19947 5287
rect 23106 5284 23112 5296
rect 19889 5247 19947 5253
rect 22480 5256 23112 5284
rect 18785 5179 18843 5185
rect 18892 5188 19012 5216
rect 19613 5219 19671 5225
rect 13262 5148 13268 5160
rect 7984 5120 10640 5148
rect 12406 5120 13268 5148
rect 7984 5108 7990 5120
rect 10410 5080 10416 5092
rect 10371 5052 10416 5080
rect 10410 5040 10416 5052
rect 10468 5040 10474 5092
rect 10612 5012 10640 5120
rect 13262 5108 13268 5120
rect 13320 5148 13326 5160
rect 14277 5151 14335 5157
rect 14277 5148 14289 5151
rect 13320 5120 14289 5148
rect 13320 5108 13326 5120
rect 14277 5117 14289 5120
rect 14323 5117 14335 5151
rect 14277 5111 14335 5117
rect 16114 5108 16120 5160
rect 16172 5148 16178 5160
rect 16172 5120 18460 5148
rect 16172 5108 16178 5120
rect 10686 5040 10692 5092
rect 10744 5080 10750 5092
rect 12802 5080 12808 5092
rect 10744 5052 12808 5080
rect 10744 5040 10750 5052
rect 12802 5040 12808 5052
rect 12860 5040 12866 5092
rect 14553 5083 14611 5089
rect 14553 5080 14565 5083
rect 13464 5052 14565 5080
rect 13464 5012 13492 5052
rect 14553 5049 14565 5052
rect 14599 5049 14611 5083
rect 14553 5043 14611 5049
rect 17773 5083 17831 5089
rect 17773 5049 17785 5083
rect 17819 5080 17831 5083
rect 18322 5080 18328 5092
rect 17819 5052 18328 5080
rect 17819 5049 17831 5052
rect 17773 5043 17831 5049
rect 18322 5040 18328 5052
rect 18380 5040 18386 5092
rect 18432 5080 18460 5120
rect 18506 5108 18512 5160
rect 18564 5148 18570 5160
rect 18892 5148 18920 5188
rect 19613 5185 19625 5219
rect 19659 5216 19671 5219
rect 20806 5216 20812 5228
rect 19659 5188 20812 5216
rect 19659 5185 19671 5188
rect 19613 5179 19671 5185
rect 20806 5176 20812 5188
rect 20864 5176 20870 5228
rect 20990 5216 20996 5228
rect 20951 5188 20996 5216
rect 20990 5176 20996 5188
rect 21048 5176 21054 5228
rect 22480 5225 22508 5256
rect 23106 5244 23112 5256
rect 23164 5244 23170 5296
rect 23652 5287 23710 5293
rect 23652 5253 23664 5287
rect 23698 5284 23710 5287
rect 25498 5284 25504 5296
rect 23698 5256 25504 5284
rect 23698 5253 23710 5256
rect 23652 5247 23710 5253
rect 25498 5244 25504 5256
rect 25556 5244 25562 5296
rect 25608 5256 25820 5284
rect 22465 5219 22523 5225
rect 22465 5185 22477 5219
rect 22511 5185 22523 5219
rect 23385 5219 23443 5225
rect 23385 5216 23397 5219
rect 22465 5179 22523 5185
rect 22572 5188 23397 5216
rect 19058 5148 19064 5160
rect 18564 5120 18920 5148
rect 19019 5120 19064 5148
rect 18564 5108 18570 5120
rect 19058 5108 19064 5120
rect 19116 5108 19122 5160
rect 21269 5151 21327 5157
rect 21269 5117 21281 5151
rect 21315 5148 21327 5151
rect 21634 5148 21640 5160
rect 21315 5120 21640 5148
rect 21315 5117 21327 5120
rect 21269 5111 21327 5117
rect 21634 5108 21640 5120
rect 21692 5108 21698 5160
rect 22002 5108 22008 5160
rect 22060 5148 22066 5160
rect 22572 5148 22600 5188
rect 23385 5185 23397 5188
rect 23431 5216 23443 5219
rect 23934 5216 23940 5228
rect 23431 5188 23940 5216
rect 23431 5185 23443 5188
rect 23385 5179 23443 5185
rect 23934 5176 23940 5188
rect 23992 5176 23998 5228
rect 24486 5176 24492 5228
rect 24544 5216 24550 5228
rect 25608 5216 25636 5256
rect 25792 5225 25820 5256
rect 25866 5244 25872 5296
rect 25924 5284 25930 5296
rect 25961 5287 26019 5293
rect 25961 5284 25973 5287
rect 25924 5256 25973 5284
rect 25924 5244 25930 5256
rect 25961 5253 25973 5256
rect 26007 5253 26019 5287
rect 35452 5284 35480 5315
rect 36722 5312 36728 5324
rect 36780 5312 36786 5364
rect 36814 5312 36820 5364
rect 36872 5352 36878 5364
rect 38381 5355 38439 5361
rect 38381 5352 38393 5355
rect 36872 5324 38393 5352
rect 36872 5312 36878 5324
rect 38381 5321 38393 5324
rect 38427 5321 38439 5355
rect 39850 5352 39856 5364
rect 39811 5324 39856 5352
rect 38381 5315 38439 5321
rect 39850 5312 39856 5324
rect 39908 5312 39914 5364
rect 40589 5355 40647 5361
rect 40589 5321 40601 5355
rect 40635 5352 40647 5355
rect 40954 5352 40960 5364
rect 40635 5324 40960 5352
rect 40635 5321 40647 5324
rect 40589 5315 40647 5321
rect 40954 5312 40960 5324
rect 41012 5312 41018 5364
rect 42150 5312 42156 5364
rect 42208 5352 42214 5364
rect 42797 5355 42855 5361
rect 42797 5352 42809 5355
rect 42208 5324 42809 5352
rect 42208 5312 42214 5324
rect 42797 5321 42809 5324
rect 42843 5321 42855 5355
rect 55582 5352 55588 5364
rect 42797 5315 42855 5321
rect 45526 5324 55588 5352
rect 35526 5284 35532 5296
rect 25961 5247 26019 5253
rect 29012 5256 35296 5284
rect 35439 5256 35532 5284
rect 24544 5188 25636 5216
rect 25777 5219 25835 5225
rect 24544 5176 24550 5188
rect 25777 5185 25789 5219
rect 25823 5185 25835 5219
rect 28074 5216 28080 5228
rect 28035 5188 28080 5216
rect 25777 5179 25835 5185
rect 28074 5176 28080 5188
rect 28132 5176 28138 5228
rect 28350 5216 28356 5228
rect 28311 5188 28356 5216
rect 28350 5176 28356 5188
rect 28408 5176 28414 5228
rect 22060 5120 22600 5148
rect 22741 5151 22799 5157
rect 22060 5108 22066 5120
rect 22741 5117 22753 5151
rect 22787 5148 22799 5151
rect 23290 5148 23296 5160
rect 22787 5120 23296 5148
rect 22787 5117 22799 5120
rect 22741 5111 22799 5117
rect 23290 5108 23296 5120
rect 23348 5108 23354 5160
rect 25593 5151 25651 5157
rect 25593 5117 25605 5151
rect 25639 5148 25651 5151
rect 26510 5148 26516 5160
rect 25639 5120 26516 5148
rect 25639 5117 25651 5120
rect 25593 5111 25651 5117
rect 26510 5108 26516 5120
rect 26568 5108 26574 5160
rect 26602 5108 26608 5160
rect 26660 5148 26666 5160
rect 29012 5148 29040 5256
rect 30558 5176 30564 5228
rect 30616 5216 30622 5228
rect 30745 5219 30803 5225
rect 30745 5216 30757 5219
rect 30616 5188 30757 5216
rect 30616 5176 30622 5188
rect 30745 5185 30757 5188
rect 30791 5216 30803 5219
rect 32398 5216 32404 5228
rect 30791 5188 32404 5216
rect 30791 5185 30803 5188
rect 30745 5179 30803 5185
rect 32398 5176 32404 5188
rect 32456 5176 32462 5228
rect 32769 5219 32827 5225
rect 32769 5185 32781 5219
rect 32815 5216 32827 5219
rect 33042 5216 33048 5228
rect 32815 5188 33048 5216
rect 32815 5185 32827 5188
rect 32769 5179 32827 5185
rect 33042 5176 33048 5188
rect 33100 5176 33106 5228
rect 33505 5219 33563 5225
rect 33505 5185 33517 5219
rect 33551 5216 33563 5219
rect 33686 5216 33692 5228
rect 33551 5188 33692 5216
rect 33551 5185 33563 5188
rect 33505 5179 33563 5185
rect 33686 5176 33692 5188
rect 33744 5176 33750 5228
rect 34606 5216 34612 5228
rect 34567 5188 34612 5216
rect 34606 5176 34612 5188
rect 34664 5176 34670 5228
rect 35268 5225 35296 5256
rect 35526 5244 35532 5256
rect 35584 5284 35590 5296
rect 35584 5256 37320 5284
rect 35584 5244 35590 5256
rect 35253 5219 35311 5225
rect 35253 5185 35265 5219
rect 35299 5185 35311 5219
rect 35253 5179 35311 5185
rect 35986 5176 35992 5228
rect 36044 5216 36050 5228
rect 36357 5219 36415 5225
rect 36357 5216 36369 5219
rect 36044 5188 36369 5216
rect 36044 5176 36050 5188
rect 36357 5185 36369 5188
rect 36403 5185 36415 5219
rect 36538 5216 36544 5228
rect 36499 5188 36544 5216
rect 36357 5179 36415 5185
rect 36538 5176 36544 5188
rect 36596 5176 36602 5228
rect 37292 5216 37320 5256
rect 37366 5244 37372 5296
rect 37424 5284 37430 5296
rect 38289 5287 38347 5293
rect 38289 5284 38301 5287
rect 37424 5256 38301 5284
rect 37424 5244 37430 5256
rect 38289 5253 38301 5256
rect 38335 5253 38347 5287
rect 43162 5284 43168 5296
rect 38289 5247 38347 5253
rect 42720 5256 43168 5284
rect 37553 5219 37611 5225
rect 37553 5216 37565 5219
rect 37292 5188 37565 5216
rect 37553 5185 37565 5188
rect 37599 5216 37611 5219
rect 38562 5216 38568 5228
rect 37599 5188 38568 5216
rect 37599 5185 37611 5188
rect 37553 5179 37611 5185
rect 38562 5176 38568 5188
rect 38620 5176 38626 5228
rect 38654 5176 38660 5228
rect 38712 5216 38718 5228
rect 39025 5219 39083 5225
rect 39025 5216 39037 5219
rect 38712 5188 39037 5216
rect 38712 5176 38718 5188
rect 39025 5185 39037 5188
rect 39071 5185 39083 5219
rect 39025 5179 39083 5185
rect 39114 5176 39120 5228
rect 39172 5216 39178 5228
rect 39669 5219 39727 5225
rect 39669 5216 39681 5219
rect 39172 5188 39681 5216
rect 39172 5176 39178 5188
rect 39669 5185 39681 5188
rect 39715 5185 39727 5219
rect 39669 5179 39727 5185
rect 40034 5176 40040 5228
rect 40092 5216 40098 5228
rect 42720 5225 42748 5256
rect 43162 5244 43168 5256
rect 43220 5284 43226 5296
rect 45526 5284 45554 5324
rect 55582 5312 55588 5324
rect 55640 5352 55646 5364
rect 56134 5352 56140 5364
rect 55640 5324 56140 5352
rect 55640 5312 55646 5324
rect 56134 5312 56140 5324
rect 56192 5352 56198 5364
rect 56192 5324 56916 5352
rect 56192 5312 56198 5324
rect 56888 5293 56916 5324
rect 43220 5256 45554 5284
rect 56873 5287 56931 5293
rect 43220 5244 43226 5256
rect 56873 5253 56885 5287
rect 56919 5253 56931 5287
rect 56873 5247 56931 5253
rect 40405 5219 40463 5225
rect 40405 5216 40417 5219
rect 40092 5188 40417 5216
rect 40092 5176 40098 5188
rect 40405 5185 40417 5188
rect 40451 5185 40463 5219
rect 40405 5179 40463 5185
rect 42705 5219 42763 5225
rect 42705 5185 42717 5219
rect 42751 5185 42763 5219
rect 43806 5216 43812 5228
rect 43767 5188 43812 5216
rect 42705 5179 42763 5185
rect 43806 5176 43812 5188
rect 43864 5176 43870 5228
rect 43990 5176 43996 5228
rect 44048 5216 44054 5228
rect 44637 5219 44695 5225
rect 44637 5216 44649 5219
rect 44048 5188 44649 5216
rect 44048 5176 44054 5188
rect 44637 5185 44649 5188
rect 44683 5185 44695 5219
rect 44637 5179 44695 5185
rect 56505 5219 56563 5225
rect 56505 5185 56517 5219
rect 56551 5216 56563 5219
rect 56594 5216 56600 5228
rect 56551 5188 56600 5216
rect 56551 5185 56563 5188
rect 56505 5179 56563 5185
rect 56594 5176 56600 5188
rect 56652 5176 56658 5228
rect 58066 5216 58072 5228
rect 58027 5188 58072 5216
rect 58066 5176 58072 5188
rect 58124 5176 58130 5228
rect 26660 5120 29040 5148
rect 26660 5108 26666 5120
rect 29546 5108 29552 5160
rect 29604 5148 29610 5160
rect 30837 5151 30895 5157
rect 30837 5148 30849 5151
rect 29604 5120 30849 5148
rect 29604 5108 29610 5120
rect 30837 5117 30849 5120
rect 30883 5117 30895 5151
rect 30837 5111 30895 5117
rect 31021 5151 31079 5157
rect 31021 5117 31033 5151
rect 31067 5148 31079 5151
rect 31110 5148 31116 5160
rect 31067 5120 31116 5148
rect 31067 5117 31079 5120
rect 31021 5111 31079 5117
rect 31110 5108 31116 5120
rect 31168 5148 31174 5160
rect 32674 5148 32680 5160
rect 31168 5120 32680 5148
rect 31168 5108 31174 5120
rect 32674 5108 32680 5120
rect 32732 5108 32738 5160
rect 32858 5108 32864 5160
rect 32916 5148 32922 5160
rect 32953 5151 33011 5157
rect 32953 5148 32965 5151
rect 32916 5120 32965 5148
rect 32916 5108 32922 5120
rect 32953 5117 32965 5120
rect 32999 5148 33011 5151
rect 33778 5148 33784 5160
rect 32999 5120 33784 5148
rect 32999 5117 33011 5120
rect 32953 5111 33011 5117
rect 33778 5108 33784 5120
rect 33836 5108 33842 5160
rect 36998 5148 37004 5160
rect 34716 5120 37004 5148
rect 25038 5080 25044 5092
rect 18432 5052 23428 5080
rect 14734 5012 14740 5024
rect 10612 4984 13492 5012
rect 14695 4984 14740 5012
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 17313 5015 17371 5021
rect 17313 4981 17325 5015
rect 17359 5012 17371 5015
rect 17954 5012 17960 5024
rect 17359 4984 17960 5012
rect 17359 4981 17371 4984
rect 17313 4975 17371 4981
rect 17954 4972 17960 4984
rect 18012 4972 18018 5024
rect 18046 4972 18052 5024
rect 18104 5012 18110 5024
rect 22922 5012 22928 5024
rect 18104 4984 22928 5012
rect 18104 4972 18110 4984
rect 22922 4972 22928 4984
rect 22980 4972 22986 5024
rect 23400 5012 23428 5052
rect 24688 5052 25044 5080
rect 24688 5012 24716 5052
rect 25038 5040 25044 5052
rect 25096 5040 25102 5092
rect 29086 5040 29092 5092
rect 29144 5080 29150 5092
rect 34716 5080 34744 5120
rect 36998 5108 37004 5120
rect 37056 5108 37062 5160
rect 37090 5108 37096 5160
rect 37148 5148 37154 5160
rect 39209 5151 39267 5157
rect 39209 5148 39221 5151
rect 37148 5120 39221 5148
rect 37148 5108 37154 5120
rect 39209 5117 39221 5120
rect 39255 5117 39267 5151
rect 39209 5111 39267 5117
rect 29144 5052 34744 5080
rect 34793 5083 34851 5089
rect 29144 5040 29150 5052
rect 34793 5049 34805 5083
rect 34839 5080 34851 5083
rect 37274 5080 37280 5092
rect 34839 5052 37280 5080
rect 34839 5049 34851 5052
rect 34793 5043 34851 5049
rect 37274 5040 37280 5052
rect 37332 5040 37338 5092
rect 37737 5083 37795 5089
rect 37737 5049 37749 5083
rect 37783 5080 37795 5083
rect 39298 5080 39304 5092
rect 37783 5052 39304 5080
rect 37783 5049 37795 5052
rect 37737 5043 37795 5049
rect 39298 5040 39304 5052
rect 39356 5040 39362 5092
rect 42058 5040 42064 5092
rect 42116 5080 42122 5092
rect 43993 5083 44051 5089
rect 43993 5080 44005 5083
rect 42116 5052 44005 5080
rect 42116 5040 42122 5052
rect 43993 5049 44005 5052
rect 44039 5049 44051 5083
rect 43993 5043 44051 5049
rect 23400 4984 24716 5012
rect 24762 4972 24768 5024
rect 24820 5012 24826 5024
rect 24820 4984 24865 5012
rect 24820 4972 24826 4984
rect 27246 4972 27252 5024
rect 27304 5012 27310 5024
rect 27433 5015 27491 5021
rect 27433 5012 27445 5015
rect 27304 4984 27445 5012
rect 27304 4972 27310 4984
rect 27433 4981 27445 4984
rect 27479 4981 27491 5015
rect 32306 5012 32312 5024
rect 32267 4984 32312 5012
rect 27433 4975 27491 4981
rect 32306 4972 32312 4984
rect 32364 4972 32370 5024
rect 44726 5012 44732 5024
rect 44687 4984 44732 5012
rect 44726 4972 44732 4984
rect 44784 4972 44790 5024
rect 58250 5012 58256 5024
rect 58211 4984 58256 5012
rect 58250 4972 58256 4984
rect 58308 4972 58314 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 9950 4768 9956 4820
rect 10008 4808 10014 4820
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 10008 4780 10609 4808
rect 10008 4768 10014 4780
rect 10597 4777 10609 4780
rect 10643 4777 10655 4811
rect 11238 4808 11244 4820
rect 10597 4771 10655 4777
rect 10796 4780 11244 4808
rect 6914 4700 6920 4752
rect 6972 4740 6978 4752
rect 9677 4743 9735 4749
rect 9677 4740 9689 4743
rect 6972 4712 9689 4740
rect 6972 4700 6978 4712
rect 9677 4709 9689 4712
rect 9723 4709 9735 4743
rect 9677 4703 9735 4709
rect 10686 4700 10692 4752
rect 10744 4700 10750 4752
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 10704 4672 10732 4700
rect 10796 4681 10824 4780
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 11606 4808 11612 4820
rect 11567 4780 11612 4808
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 11716 4780 11928 4808
rect 11716 4740 11744 4780
rect 10888 4712 11744 4740
rect 11900 4740 11928 4780
rect 11974 4768 11980 4820
rect 12032 4808 12038 4820
rect 12805 4811 12863 4817
rect 12805 4808 12817 4811
rect 12032 4780 12817 4808
rect 12032 4768 12038 4780
rect 12805 4777 12817 4780
rect 12851 4777 12863 4811
rect 12805 4771 12863 4777
rect 18141 4811 18199 4817
rect 18141 4777 18153 4811
rect 18187 4808 18199 4811
rect 18598 4808 18604 4820
rect 18187 4780 18604 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 20990 4808 20996 4820
rect 20951 4780 20996 4808
rect 20990 4768 20996 4780
rect 21048 4768 21054 4820
rect 22005 4811 22063 4817
rect 22005 4777 22017 4811
rect 22051 4808 22063 4811
rect 23014 4808 23020 4820
rect 22051 4780 23020 4808
rect 22051 4777 22063 4780
rect 22005 4771 22063 4777
rect 23014 4768 23020 4780
rect 23072 4768 23078 4820
rect 30558 4808 30564 4820
rect 24688 4780 30564 4808
rect 16114 4740 16120 4752
rect 11900 4712 16120 4740
rect 10888 4681 10916 4712
rect 16114 4700 16120 4712
rect 16172 4700 16178 4752
rect 16209 4743 16267 4749
rect 16209 4709 16221 4743
rect 16255 4740 16267 4743
rect 21821 4743 21879 4749
rect 21821 4740 21833 4743
rect 16255 4712 21833 4740
rect 16255 4709 16267 4712
rect 16209 4703 16267 4709
rect 21821 4709 21833 4712
rect 21867 4709 21879 4743
rect 21821 4703 21879 4709
rect 22278 4700 22284 4752
rect 22336 4740 22342 4752
rect 22465 4743 22523 4749
rect 22465 4740 22477 4743
rect 22336 4712 22477 4740
rect 22336 4700 22342 4712
rect 22465 4709 22477 4712
rect 22511 4709 22523 4743
rect 24688 4740 24716 4780
rect 30558 4768 30564 4780
rect 30616 4768 30622 4820
rect 33594 4768 33600 4820
rect 33652 4808 33658 4820
rect 40957 4811 41015 4817
rect 40957 4808 40969 4811
rect 33652 4780 40969 4808
rect 33652 4768 33658 4780
rect 40957 4777 40969 4780
rect 41003 4777 41015 4811
rect 41690 4808 41696 4820
rect 41651 4780 41696 4808
rect 40957 4771 41015 4777
rect 41690 4768 41696 4780
rect 41748 4768 41754 4820
rect 43622 4768 43628 4820
rect 43680 4808 43686 4820
rect 45373 4811 45431 4817
rect 45373 4808 45385 4811
rect 43680 4780 45385 4808
rect 43680 4768 43686 4780
rect 45373 4777 45385 4780
rect 45419 4777 45431 4811
rect 47578 4808 47584 4820
rect 47539 4780 47584 4808
rect 45373 4771 45431 4777
rect 47578 4768 47584 4780
rect 47636 4768 47642 4820
rect 55398 4768 55404 4820
rect 55456 4808 55462 4820
rect 58069 4811 58127 4817
rect 58069 4808 58081 4811
rect 55456 4780 58081 4808
rect 55456 4768 55462 4780
rect 58069 4777 58081 4780
rect 58115 4777 58127 4811
rect 58069 4771 58127 4777
rect 22465 4703 22523 4709
rect 22756 4712 24716 4740
rect 8619 4644 10732 4672
rect 10781 4675 10839 4681
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 10781 4641 10793 4675
rect 10827 4641 10839 4675
rect 10781 4635 10839 4641
rect 10873 4675 10931 4681
rect 10873 4641 10885 4675
rect 10919 4641 10931 4675
rect 10873 4635 10931 4641
rect 10965 4675 11023 4681
rect 10965 4641 10977 4675
rect 11011 4672 11023 4675
rect 11011 4644 11192 4672
rect 11011 4641 11023 4644
rect 10965 4635 11023 4641
rect 1581 4607 1639 4613
rect 1581 4573 1593 4607
rect 1627 4604 1639 4607
rect 8294 4604 8300 4616
rect 1627 4576 8300 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 9582 4604 9588 4616
rect 9447 4576 9588 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 9582 4564 9588 4576
rect 9640 4604 9646 4616
rect 10980 4604 11008 4635
rect 11164 4616 11192 4644
rect 11606 4632 11612 4684
rect 11664 4672 11670 4684
rect 11785 4675 11843 4681
rect 11785 4672 11797 4675
rect 11664 4644 11797 4672
rect 11664 4632 11670 4644
rect 11785 4641 11797 4644
rect 11831 4641 11843 4675
rect 11785 4635 11843 4641
rect 11885 4675 11943 4681
rect 11885 4641 11897 4675
rect 11931 4672 11943 4675
rect 18046 4672 18052 4684
rect 11931 4644 18052 4672
rect 11931 4641 11943 4644
rect 11885 4635 11943 4641
rect 18046 4632 18052 4644
rect 18104 4632 18110 4684
rect 18785 4675 18843 4681
rect 18432 4644 18736 4672
rect 9640 4576 11008 4604
rect 11057 4607 11115 4613
rect 9640 4564 9646 4576
rect 11057 4573 11069 4607
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 1854 4536 1860 4548
rect 1815 4508 1860 4536
rect 1854 4496 1860 4508
rect 1912 4496 1918 4548
rect 7282 4496 7288 4548
rect 7340 4536 7346 4548
rect 7469 4539 7527 4545
rect 7469 4536 7481 4539
rect 7340 4508 7481 4536
rect 7340 4496 7346 4508
rect 7469 4505 7481 4508
rect 7515 4505 7527 4539
rect 7469 4499 7527 4505
rect 8389 4539 8447 4545
rect 8389 4505 8401 4539
rect 8435 4536 8447 4539
rect 8570 4536 8576 4548
rect 8435 4508 8576 4536
rect 8435 4505 8447 4508
rect 8389 4499 8447 4505
rect 8570 4496 8576 4508
rect 8628 4496 8634 4548
rect 10318 4536 10324 4548
rect 9784 4508 10324 4536
rect 7558 4468 7564 4480
rect 7519 4440 7564 4468
rect 7558 4428 7564 4440
rect 7616 4428 7622 4480
rect 8754 4428 8760 4480
rect 8812 4468 8818 4480
rect 9784 4468 9812 4508
rect 10318 4496 10324 4508
rect 10376 4496 10382 4548
rect 11072 4536 11100 4567
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11974 4604 11980 4616
rect 11204 4576 11980 4604
rect 11204 4564 11210 4576
rect 11974 4564 11980 4576
rect 12032 4564 12038 4616
rect 12066 4564 12072 4616
rect 12124 4604 12130 4616
rect 12124 4576 12169 4604
rect 12124 4564 12130 4576
rect 12342 4564 12348 4616
rect 12400 4604 12406 4616
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12400 4576 12725 4604
rect 12400 4564 12406 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 17037 4607 17095 4613
rect 17037 4573 17049 4607
rect 17083 4604 17095 4607
rect 18432 4604 18460 4644
rect 17083 4576 18460 4604
rect 18708 4604 18736 4644
rect 18785 4641 18797 4675
rect 18831 4672 18843 4675
rect 19058 4672 19064 4684
rect 18831 4644 19064 4672
rect 18831 4641 18843 4644
rect 18785 4635 18843 4641
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 20165 4675 20223 4681
rect 20165 4641 20177 4675
rect 20211 4672 20223 4675
rect 20622 4672 20628 4684
rect 20211 4644 20628 4672
rect 20211 4641 20223 4644
rect 20165 4635 20223 4641
rect 20622 4632 20628 4644
rect 20680 4632 20686 4684
rect 22186 4672 22192 4684
rect 20824 4644 22192 4672
rect 19794 4604 19800 4616
rect 18708 4576 19800 4604
rect 17083 4573 17095 4576
rect 17037 4567 17095 4573
rect 19794 4564 19800 4576
rect 19852 4564 19858 4616
rect 19889 4607 19947 4613
rect 19889 4573 19901 4607
rect 19935 4604 19947 4607
rect 20824 4604 20852 4644
rect 22186 4632 22192 4644
rect 22244 4632 22250 4684
rect 19935 4576 20852 4604
rect 20901 4607 20959 4613
rect 19935 4573 19947 4576
rect 19889 4567 19947 4573
rect 20901 4573 20913 4607
rect 20947 4604 20959 4607
rect 21266 4604 21272 4616
rect 20947 4576 21272 4604
rect 20947 4573 20959 4576
rect 20901 4567 20959 4573
rect 21266 4564 21272 4576
rect 21324 4564 21330 4616
rect 22756 4604 22784 4712
rect 24762 4700 24768 4752
rect 24820 4740 24826 4752
rect 29086 4740 29092 4752
rect 24820 4712 29092 4740
rect 24820 4700 24826 4712
rect 29086 4700 29092 4712
rect 29144 4700 29150 4752
rect 39117 4743 39175 4749
rect 31956 4712 33640 4740
rect 22922 4672 22928 4684
rect 22883 4644 22928 4672
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 23109 4675 23167 4681
rect 23109 4641 23121 4675
rect 23155 4672 23167 4675
rect 25038 4672 25044 4684
rect 23155 4644 24808 4672
rect 24999 4644 25044 4672
rect 23155 4641 23167 4644
rect 23109 4635 23167 4641
rect 21376 4576 22784 4604
rect 12434 4536 12440 4548
rect 11072 4508 12440 4536
rect 12434 4496 12440 4508
rect 12492 4496 12498 4548
rect 14645 4539 14703 4545
rect 14645 4505 14657 4539
rect 14691 4536 14703 4539
rect 14918 4536 14924 4548
rect 14691 4508 14924 4536
rect 14691 4505 14703 4508
rect 14645 4499 14703 4505
rect 14918 4496 14924 4508
rect 14976 4496 14982 4548
rect 15838 4496 15844 4548
rect 15896 4536 15902 4548
rect 16025 4539 16083 4545
rect 16025 4536 16037 4539
rect 15896 4508 16037 4536
rect 15896 4496 15902 4508
rect 16025 4505 16037 4508
rect 16071 4505 16083 4539
rect 16025 4499 16083 4505
rect 16942 4496 16948 4548
rect 17000 4536 17006 4548
rect 17313 4539 17371 4545
rect 17313 4536 17325 4539
rect 17000 4508 17325 4536
rect 17000 4496 17006 4508
rect 17313 4505 17325 4508
rect 17359 4505 17371 4539
rect 17313 4499 17371 4505
rect 18601 4539 18659 4545
rect 18601 4505 18613 4539
rect 18647 4536 18659 4539
rect 21376 4536 21404 4576
rect 22830 4564 22836 4616
rect 22888 4604 22894 4616
rect 22888 4576 22933 4604
rect 22888 4564 22894 4576
rect 18647 4508 21404 4536
rect 21545 4539 21603 4545
rect 18647 4505 18659 4508
rect 18601 4499 18659 4505
rect 21545 4505 21557 4539
rect 21591 4536 21603 4539
rect 21726 4536 21732 4548
rect 21591 4508 21732 4536
rect 21591 4505 21603 4508
rect 21545 4499 21603 4505
rect 21726 4496 21732 4508
rect 21784 4496 21790 4548
rect 23124 4536 23152 4635
rect 22940 4508 23152 4536
rect 24780 4536 24808 4644
rect 25038 4632 25044 4644
rect 25096 4632 25102 4684
rect 25133 4675 25191 4681
rect 25133 4641 25145 4675
rect 25179 4672 25191 4675
rect 26418 4672 26424 4684
rect 25179 4644 26424 4672
rect 25179 4641 25191 4644
rect 25133 4635 25191 4641
rect 24946 4604 24952 4616
rect 24907 4576 24952 4604
rect 24946 4564 24952 4576
rect 25004 4564 25010 4616
rect 25148 4548 25176 4635
rect 26418 4632 26424 4644
rect 26476 4632 26482 4684
rect 26878 4632 26884 4684
rect 26936 4672 26942 4684
rect 31956 4672 31984 4712
rect 32122 4672 32128 4684
rect 26936 4644 30236 4672
rect 26936 4632 26942 4644
rect 26605 4607 26663 4613
rect 26605 4573 26617 4607
rect 26651 4604 26663 4607
rect 27430 4604 27436 4616
rect 26651 4576 27436 4604
rect 26651 4573 26663 4576
rect 26605 4567 26663 4573
rect 27430 4564 27436 4576
rect 27488 4564 27494 4616
rect 27614 4564 27620 4616
rect 27672 4604 27678 4616
rect 28902 4604 28908 4616
rect 27672 4576 28908 4604
rect 27672 4564 27678 4576
rect 28902 4564 28908 4576
rect 28960 4564 28966 4616
rect 28997 4607 29055 4613
rect 28997 4573 29009 4607
rect 29043 4604 29055 4607
rect 30098 4604 30104 4616
rect 29043 4576 30104 4604
rect 29043 4573 29055 4576
rect 28997 4567 29055 4573
rect 30098 4564 30104 4576
rect 30156 4564 30162 4616
rect 25130 4536 25136 4548
rect 24780 4508 25136 4536
rect 8812 4440 9812 4468
rect 9861 4471 9919 4477
rect 8812 4428 8818 4440
rect 9861 4437 9873 4471
rect 9907 4468 9919 4471
rect 10226 4468 10232 4480
rect 9907 4440 10232 4468
rect 9907 4437 9919 4440
rect 9861 4431 9919 4437
rect 10226 4428 10232 4440
rect 10284 4428 10290 4480
rect 11238 4428 11244 4480
rect 11296 4468 11302 4480
rect 12342 4468 12348 4480
rect 11296 4440 12348 4468
rect 11296 4428 11302 4440
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 14734 4468 14740 4480
rect 14695 4440 14740 4468
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 18506 4428 18512 4480
rect 18564 4468 18570 4480
rect 18564 4440 18609 4468
rect 18564 4428 18570 4440
rect 19334 4428 19340 4480
rect 19392 4468 19398 4480
rect 19521 4471 19579 4477
rect 19521 4468 19533 4471
rect 19392 4440 19533 4468
rect 19392 4428 19398 4440
rect 19521 4437 19533 4440
rect 19567 4437 19579 4471
rect 19978 4468 19984 4480
rect 19939 4440 19984 4468
rect 19521 4431 19579 4437
rect 19978 4428 19984 4440
rect 20036 4428 20042 4480
rect 20622 4428 20628 4480
rect 20680 4468 20686 4480
rect 22940 4468 22968 4508
rect 25130 4496 25136 4508
rect 25188 4496 25194 4548
rect 27709 4539 27767 4545
rect 27709 4505 27721 4539
rect 27755 4536 27767 4539
rect 28442 4536 28448 4548
rect 27755 4508 28448 4536
rect 27755 4505 27767 4508
rect 27709 4499 27767 4505
rect 28442 4496 28448 4508
rect 28500 4496 28506 4548
rect 28534 4496 28540 4548
rect 28592 4536 28598 4548
rect 30006 4536 30012 4548
rect 28592 4508 30012 4536
rect 28592 4496 28598 4508
rect 30006 4496 30012 4508
rect 30064 4496 30070 4548
rect 24578 4468 24584 4480
rect 20680 4440 22968 4468
rect 24539 4440 24584 4468
rect 20680 4428 20686 4440
rect 24578 4428 24584 4440
rect 24636 4428 24642 4480
rect 27065 4471 27123 4477
rect 27065 4437 27077 4471
rect 27111 4468 27123 4471
rect 28258 4468 28264 4480
rect 27111 4440 28264 4468
rect 27111 4437 27123 4440
rect 27065 4431 27123 4437
rect 28258 4428 28264 4440
rect 28316 4428 28322 4480
rect 28353 4471 28411 4477
rect 28353 4437 28365 4471
rect 28399 4468 28411 4471
rect 28994 4468 29000 4480
rect 28399 4440 29000 4468
rect 28399 4437 28411 4440
rect 28353 4431 28411 4437
rect 28994 4428 29000 4440
rect 29052 4428 29058 4480
rect 29086 4428 29092 4480
rect 29144 4468 29150 4480
rect 30208 4468 30236 4644
rect 31588 4644 31984 4672
rect 32083 4644 32128 4672
rect 30285 4607 30343 4613
rect 30285 4573 30297 4607
rect 30331 4604 30343 4607
rect 30926 4604 30932 4616
rect 30331 4576 30932 4604
rect 30331 4573 30343 4576
rect 30285 4567 30343 4573
rect 30926 4564 30932 4576
rect 30984 4564 30990 4616
rect 30552 4539 30610 4545
rect 30552 4505 30564 4539
rect 30598 4536 30610 4539
rect 30650 4536 30656 4548
rect 30598 4508 30656 4536
rect 30598 4505 30610 4508
rect 30552 4499 30610 4505
rect 30650 4496 30656 4508
rect 30708 4496 30714 4548
rect 31588 4468 31616 4644
rect 32122 4632 32128 4644
rect 32180 4632 32186 4684
rect 32306 4604 32312 4616
rect 32267 4576 32312 4604
rect 32306 4564 32312 4576
rect 32364 4564 32370 4616
rect 33612 4613 33640 4712
rect 39117 4709 39129 4743
rect 39163 4740 39175 4743
rect 39574 4740 39580 4752
rect 39163 4712 39580 4740
rect 39163 4709 39175 4712
rect 39117 4703 39175 4709
rect 39574 4700 39580 4712
rect 39632 4700 39638 4752
rect 43254 4740 43260 4752
rect 43215 4712 43260 4740
rect 43254 4700 43260 4712
rect 43312 4700 43318 4752
rect 44174 4740 44180 4752
rect 44135 4712 44180 4740
rect 44174 4700 44180 4712
rect 44232 4700 44238 4752
rect 45186 4700 45192 4752
rect 45244 4740 45250 4752
rect 48317 4743 48375 4749
rect 48317 4740 48329 4743
rect 45244 4712 48329 4740
rect 45244 4700 45250 4712
rect 48317 4709 48329 4712
rect 48363 4709 48375 4743
rect 48317 4703 48375 4709
rect 38381 4675 38439 4681
rect 38381 4672 38393 4675
rect 36096 4644 38393 4672
rect 33597 4607 33655 4613
rect 33597 4573 33609 4607
rect 33643 4604 33655 4607
rect 34422 4604 34428 4616
rect 33643 4576 34428 4604
rect 33643 4573 33655 4576
rect 33597 4567 33655 4573
rect 34422 4564 34428 4576
rect 34480 4564 34486 4616
rect 34790 4564 34796 4616
rect 34848 4604 34854 4616
rect 36096 4613 36124 4644
rect 38381 4641 38393 4644
rect 38427 4641 38439 4675
rect 39482 4672 39488 4684
rect 38381 4635 38439 4641
rect 38488 4644 39488 4672
rect 34885 4607 34943 4613
rect 34885 4604 34897 4607
rect 34848 4576 34897 4604
rect 34848 4564 34854 4576
rect 34885 4573 34897 4576
rect 34931 4573 34943 4607
rect 34885 4567 34943 4573
rect 36081 4607 36139 4613
rect 36081 4573 36093 4607
rect 36127 4573 36139 4607
rect 36081 4567 36139 4573
rect 36170 4564 36176 4616
rect 36228 4604 36234 4616
rect 37182 4604 37188 4616
rect 36228 4576 37188 4604
rect 36228 4564 36234 4576
rect 37182 4564 37188 4576
rect 37240 4564 37246 4616
rect 38197 4607 38255 4613
rect 38197 4573 38209 4607
rect 38243 4604 38255 4607
rect 38488 4604 38516 4644
rect 39482 4632 39488 4644
rect 39540 4632 39546 4684
rect 45462 4632 45468 4684
rect 45520 4672 45526 4684
rect 46842 4672 46848 4684
rect 45520 4644 46848 4672
rect 45520 4632 45526 4644
rect 46842 4632 46848 4644
rect 46900 4632 46906 4684
rect 56594 4632 56600 4684
rect 56652 4672 56658 4684
rect 57333 4675 57391 4681
rect 57333 4672 57345 4675
rect 56652 4644 57345 4672
rect 56652 4632 56658 4644
rect 57333 4641 57345 4644
rect 57379 4641 57391 4675
rect 57333 4635 57391 4641
rect 38562 4604 38568 4616
rect 38243 4576 38568 4604
rect 38243 4573 38255 4576
rect 38197 4567 38255 4573
rect 38562 4564 38568 4576
rect 38620 4564 38626 4616
rect 39206 4564 39212 4616
rect 39264 4604 39270 4616
rect 40865 4607 40923 4613
rect 40865 4604 40877 4607
rect 39264 4576 40877 4604
rect 39264 4564 39270 4576
rect 40865 4573 40877 4576
rect 40911 4573 40923 4607
rect 40865 4567 40923 4573
rect 45922 4564 45928 4616
rect 45980 4604 45986 4616
rect 45980 4576 46152 4604
rect 45980 4564 45986 4576
rect 32398 4536 32404 4548
rect 31680 4508 32404 4536
rect 31680 4477 31708 4508
rect 32398 4496 32404 4508
rect 32456 4496 32462 4548
rect 34606 4496 34612 4548
rect 34664 4536 34670 4548
rect 35161 4539 35219 4545
rect 35161 4536 35173 4539
rect 34664 4508 35173 4536
rect 34664 4496 34670 4508
rect 35161 4505 35173 4508
rect 35207 4505 35219 4539
rect 36357 4539 36415 4545
rect 36357 4536 36369 4539
rect 35161 4499 35219 4505
rect 36096 4508 36369 4536
rect 36096 4480 36124 4508
rect 36357 4505 36369 4508
rect 36403 4505 36415 4539
rect 36357 4499 36415 4505
rect 37090 4496 37096 4548
rect 37148 4536 37154 4548
rect 37461 4539 37519 4545
rect 37461 4536 37473 4539
rect 37148 4508 37473 4536
rect 37148 4496 37154 4508
rect 37461 4505 37473 4508
rect 37507 4505 37519 4539
rect 38930 4536 38936 4548
rect 38891 4508 38936 4536
rect 37461 4499 37519 4505
rect 38930 4496 38936 4508
rect 38988 4496 38994 4548
rect 40129 4539 40187 4545
rect 40129 4536 40141 4539
rect 39040 4508 40141 4536
rect 29144 4440 29189 4468
rect 30208 4440 31616 4468
rect 31665 4471 31723 4477
rect 29144 4428 29150 4440
rect 31665 4437 31677 4471
rect 31711 4437 31723 4471
rect 31665 4431 31723 4437
rect 32306 4428 32312 4480
rect 32364 4468 32370 4480
rect 32493 4471 32551 4477
rect 32493 4468 32505 4471
rect 32364 4440 32505 4468
rect 32364 4428 32370 4440
rect 32493 4437 32505 4440
rect 32539 4437 32551 4471
rect 32493 4431 32551 4437
rect 33689 4471 33747 4477
rect 33689 4437 33701 4471
rect 33735 4468 33747 4471
rect 35802 4468 35808 4480
rect 33735 4440 35808 4468
rect 33735 4437 33747 4440
rect 33689 4431 33747 4437
rect 35802 4428 35808 4440
rect 35860 4428 35866 4480
rect 36078 4428 36084 4480
rect 36136 4428 36142 4480
rect 38470 4428 38476 4480
rect 38528 4468 38534 4480
rect 39040 4468 39068 4508
rect 40129 4505 40141 4508
rect 40175 4505 40187 4539
rect 40129 4499 40187 4505
rect 41414 4496 41420 4548
rect 41472 4536 41478 4548
rect 41601 4539 41659 4545
rect 41601 4536 41613 4539
rect 41472 4508 41613 4536
rect 41472 4496 41478 4508
rect 41601 4505 41613 4508
rect 41647 4505 41659 4539
rect 41601 4499 41659 4505
rect 42058 4496 42064 4548
rect 42116 4536 42122 4548
rect 42337 4539 42395 4545
rect 42337 4536 42349 4539
rect 42116 4508 42349 4536
rect 42116 4496 42122 4508
rect 42337 4505 42349 4508
rect 42383 4505 42395 4539
rect 42337 4499 42395 4505
rect 42521 4539 42579 4545
rect 42521 4505 42533 4539
rect 42567 4536 42579 4539
rect 42886 4536 42892 4548
rect 42567 4508 42892 4536
rect 42567 4505 42579 4508
rect 42521 4499 42579 4505
rect 42886 4496 42892 4508
rect 42944 4496 42950 4548
rect 42978 4496 42984 4548
rect 43036 4536 43042 4548
rect 43073 4539 43131 4545
rect 43073 4536 43085 4539
rect 43036 4508 43085 4536
rect 43036 4496 43042 4508
rect 43073 4505 43085 4508
rect 43119 4505 43131 4539
rect 43073 4499 43131 4505
rect 43162 4496 43168 4548
rect 43220 4536 43226 4548
rect 43993 4539 44051 4545
rect 43993 4536 44005 4539
rect 43220 4508 44005 4536
rect 43220 4496 43226 4508
rect 43993 4505 44005 4508
rect 44039 4505 44051 4539
rect 43993 4499 44051 4505
rect 44358 4496 44364 4548
rect 44416 4536 44422 4548
rect 45281 4539 45339 4545
rect 45281 4536 45293 4539
rect 44416 4508 45293 4536
rect 44416 4496 44422 4508
rect 45281 4505 45293 4508
rect 45327 4505 45339 4539
rect 46017 4539 46075 4545
rect 46017 4536 46029 4539
rect 45281 4499 45339 4505
rect 45526 4508 46029 4536
rect 38528 4440 39068 4468
rect 38528 4428 38534 4440
rect 39114 4428 39120 4480
rect 39172 4468 39178 4480
rect 40221 4471 40279 4477
rect 40221 4468 40233 4471
rect 39172 4440 40233 4468
rect 39172 4428 39178 4440
rect 40221 4437 40233 4440
rect 40267 4437 40279 4471
rect 40221 4431 40279 4437
rect 45002 4428 45008 4480
rect 45060 4468 45066 4480
rect 45526 4468 45554 4508
rect 46017 4505 46029 4508
rect 46063 4505 46075 4539
rect 46124 4536 46152 4576
rect 46566 4564 46572 4616
rect 46624 4604 46630 4616
rect 47397 4607 47455 4613
rect 47397 4604 47409 4607
rect 46624 4576 47409 4604
rect 46624 4564 46630 4576
rect 47397 4573 47409 4576
rect 47443 4573 47455 4607
rect 47397 4567 47455 4573
rect 47486 4564 47492 4616
rect 47544 4604 47550 4616
rect 48133 4607 48191 4613
rect 48133 4604 48145 4607
rect 47544 4576 48145 4604
rect 47544 4564 47550 4576
rect 48133 4573 48145 4576
rect 48179 4573 48191 4607
rect 57974 4604 57980 4616
rect 57935 4576 57980 4604
rect 48133 4567 48191 4573
rect 57974 4564 57980 4576
rect 58032 4564 58038 4616
rect 58158 4604 58164 4616
rect 58119 4576 58164 4604
rect 58158 4564 58164 4576
rect 58216 4564 58222 4616
rect 46753 4539 46811 4545
rect 46753 4536 46765 4539
rect 46124 4508 46765 4536
rect 46017 4499 46075 4505
rect 46753 4505 46765 4508
rect 46799 4505 46811 4539
rect 56594 4536 56600 4548
rect 56555 4508 56600 4536
rect 46753 4499 46811 4505
rect 56594 4496 56600 4508
rect 56652 4496 56658 4548
rect 45060 4440 45554 4468
rect 45060 4428 45066 4440
rect 45738 4428 45744 4480
rect 45796 4468 45802 4480
rect 46109 4471 46167 4477
rect 46109 4468 46121 4471
rect 45796 4440 46121 4468
rect 45796 4428 45802 4440
rect 46109 4437 46121 4440
rect 46155 4437 46167 4471
rect 46109 4431 46167 4437
rect 46198 4428 46204 4480
rect 46256 4468 46262 4480
rect 46845 4471 46903 4477
rect 46845 4468 46857 4471
rect 46256 4440 46857 4468
rect 46256 4428 46262 4440
rect 46845 4437 46857 4440
rect 46891 4437 46903 4471
rect 46845 4431 46903 4437
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 7558 4224 7564 4276
rect 7616 4264 7622 4276
rect 18506 4264 18512 4276
rect 7616 4236 18512 4264
rect 7616 4224 7622 4236
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 18985 4236 19196 4264
rect 7285 4199 7343 4205
rect 7285 4165 7297 4199
rect 7331 4196 7343 4199
rect 7834 4196 7840 4208
rect 7331 4168 7840 4196
rect 7331 4165 7343 4168
rect 7285 4159 7343 4165
rect 7834 4156 7840 4168
rect 7892 4156 7898 4208
rect 8021 4199 8079 4205
rect 8021 4165 8033 4199
rect 8067 4196 8079 4199
rect 9490 4196 9496 4208
rect 8067 4168 9496 4196
rect 8067 4165 8079 4168
rect 8021 4159 8079 4165
rect 9490 4156 9496 4168
rect 9548 4156 9554 4208
rect 10870 4196 10876 4208
rect 10520 4168 10876 4196
rect 1581 4131 1639 4137
rect 1581 4097 1593 4131
rect 1627 4128 1639 4131
rect 8662 4128 8668 4140
rect 1627 4100 8668 4128
rect 1627 4097 1639 4100
rect 1581 4091 1639 4097
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 8754 4088 8760 4140
rect 8812 4128 8818 4140
rect 8941 4131 8999 4137
rect 8812 4100 8857 4128
rect 8812 4088 8818 4100
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 10520 4128 10548 4168
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 11330 4156 11336 4208
rect 11388 4196 11394 4208
rect 12529 4199 12587 4205
rect 12529 4196 12541 4199
rect 11388 4168 11744 4196
rect 11388 4156 11394 4168
rect 8987 4100 10548 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 11146 4128 11152 4140
rect 10744 4100 11152 4128
rect 10744 4088 10750 4100
rect 11146 4088 11152 4100
rect 11204 4088 11210 4140
rect 11716 4128 11744 4168
rect 12176 4168 12541 4196
rect 12176 4128 12204 4168
rect 12529 4165 12541 4168
rect 12575 4165 12587 4199
rect 12529 4159 12587 4165
rect 12618 4156 12624 4208
rect 12676 4196 12682 4208
rect 18985 4196 19013 4236
rect 12676 4168 19013 4196
rect 19168 4196 19196 4236
rect 19518 4224 19524 4276
rect 19576 4264 19582 4276
rect 19978 4264 19984 4276
rect 19576 4236 19984 4264
rect 19576 4224 19582 4236
rect 19978 4224 19984 4236
rect 20036 4264 20042 4276
rect 20530 4264 20536 4276
rect 20036 4236 20536 4264
rect 20036 4224 20042 4236
rect 20530 4224 20536 4236
rect 20588 4224 20594 4276
rect 22922 4224 22928 4276
rect 22980 4264 22986 4276
rect 23385 4267 23443 4273
rect 23385 4264 23397 4267
rect 22980 4236 23397 4264
rect 22980 4224 22986 4236
rect 23385 4233 23397 4236
rect 23431 4233 23443 4267
rect 23385 4227 23443 4233
rect 23492 4236 24716 4264
rect 23492 4196 23520 4236
rect 19168 4168 23520 4196
rect 24204 4199 24262 4205
rect 12676 4156 12682 4168
rect 24204 4165 24216 4199
rect 24250 4196 24262 4199
rect 24578 4196 24584 4208
rect 24250 4168 24584 4196
rect 24250 4165 24262 4168
rect 24204 4159 24262 4165
rect 24578 4156 24584 4168
rect 24636 4156 24642 4208
rect 24688 4196 24716 4236
rect 25038 4224 25044 4276
rect 25096 4264 25102 4276
rect 25317 4267 25375 4273
rect 25317 4264 25329 4267
rect 25096 4236 25329 4264
rect 25096 4224 25102 4236
rect 25317 4233 25329 4236
rect 25363 4233 25375 4267
rect 25317 4227 25375 4233
rect 27525 4267 27583 4273
rect 27525 4233 27537 4267
rect 27571 4264 27583 4267
rect 29546 4264 29552 4276
rect 27571 4236 29552 4264
rect 27571 4233 27583 4236
rect 27525 4227 27583 4233
rect 29546 4224 29552 4236
rect 29604 4224 29610 4276
rect 29641 4267 29699 4273
rect 29641 4233 29653 4267
rect 29687 4264 29699 4267
rect 30190 4264 30196 4276
rect 29687 4236 30196 4264
rect 29687 4233 29699 4236
rect 29641 4227 29699 4233
rect 30190 4224 30196 4236
rect 30248 4264 30254 4276
rect 33042 4264 33048 4276
rect 30248 4236 33048 4264
rect 30248 4224 30254 4236
rect 33042 4224 33048 4236
rect 33100 4264 33106 4276
rect 58250 4264 58256 4276
rect 33100 4236 58256 4264
rect 33100 4224 33106 4236
rect 58250 4224 58256 4236
rect 58308 4224 58314 4276
rect 28445 4199 28503 4205
rect 28445 4196 28457 4199
rect 24688 4168 28457 4196
rect 28445 4165 28457 4168
rect 28491 4196 28503 4199
rect 29086 4196 29092 4208
rect 28491 4168 29092 4196
rect 28491 4165 28503 4168
rect 28445 4159 28503 4165
rect 29086 4156 29092 4168
rect 29144 4196 29150 4208
rect 30098 4196 30104 4208
rect 29144 4168 30104 4196
rect 29144 4156 29150 4168
rect 30098 4156 30104 4168
rect 30156 4196 30162 4208
rect 30561 4199 30619 4205
rect 30561 4196 30573 4199
rect 30156 4168 30573 4196
rect 30156 4156 30162 4168
rect 30561 4165 30573 4168
rect 30607 4165 30619 4199
rect 30561 4159 30619 4165
rect 30668 4168 31708 4196
rect 12342 4128 12348 4140
rect 11716 4100 12204 4128
rect 12303 4100 12348 4128
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 13906 4128 13912 4140
rect 13311 4100 13912 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 13906 4088 13912 4100
rect 13964 4128 13970 4140
rect 14734 4128 14740 4140
rect 13964 4100 14740 4128
rect 13964 4088 13970 4100
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 15654 4128 15660 4140
rect 14976 4100 15660 4128
rect 14976 4088 14982 4100
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4128 15899 4131
rect 16850 4128 16856 4140
rect 15887 4100 16712 4128
rect 16811 4100 16856 4128
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 1762 4060 1768 4072
rect 1723 4032 1768 4060
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4060 7527 4063
rect 7650 4060 7656 4072
rect 7515 4032 7656 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 7650 4020 7656 4032
rect 7708 4020 7714 4072
rect 9401 4063 9459 4069
rect 9401 4029 9413 4063
rect 9447 4060 9459 4063
rect 9582 4060 9588 4072
rect 9447 4032 9588 4060
rect 9447 4029 9459 4032
rect 9401 4023 9459 4029
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 9858 4020 9864 4072
rect 9916 4060 9922 4072
rect 10321 4063 10379 4069
rect 10321 4060 10333 4063
rect 9916 4032 10333 4060
rect 9916 4020 9922 4032
rect 10321 4029 10333 4032
rect 10367 4029 10379 4063
rect 10502 4060 10508 4072
rect 10463 4032 10508 4060
rect 10321 4023 10379 4029
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 10597 4063 10655 4069
rect 10597 4029 10609 4063
rect 10643 4029 10655 4063
rect 10597 4023 10655 4029
rect 8205 3995 8263 4001
rect 8205 3961 8217 3995
rect 8251 3992 8263 3995
rect 9677 3995 9735 4001
rect 9677 3992 9689 3995
rect 8251 3964 9689 3992
rect 8251 3961 8263 3964
rect 8205 3955 8263 3961
rect 9677 3961 9689 3964
rect 9723 3961 9735 3995
rect 10612 3992 10640 4023
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 10836 4032 10881 4060
rect 10836 4020 10842 4032
rect 10962 4020 10968 4072
rect 11020 4060 11026 4072
rect 11422 4060 11428 4072
rect 11020 4032 11428 4060
rect 11020 4020 11026 4032
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 11606 4020 11612 4072
rect 11664 4060 11670 4072
rect 12713 4063 12771 4069
rect 12713 4060 12725 4063
rect 11664 4032 12725 4060
rect 11664 4020 11670 4032
rect 12713 4029 12725 4032
rect 12759 4060 12771 4063
rect 12802 4060 12808 4072
rect 12759 4032 12808 4060
rect 12759 4029 12771 4032
rect 12713 4023 12771 4029
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 14001 4063 14059 4069
rect 14001 4029 14013 4063
rect 14047 4060 14059 4063
rect 14090 4060 14096 4072
rect 14047 4032 14096 4060
rect 14047 4029 14059 4032
rect 14001 4023 14059 4029
rect 14090 4020 14096 4032
rect 14148 4020 14154 4072
rect 16117 4063 16175 4069
rect 16117 4029 16129 4063
rect 16163 4060 16175 4063
rect 16684 4060 16712 4100
rect 16850 4088 16856 4100
rect 16908 4088 16914 4140
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 17552 4100 17785 4128
rect 17552 4088 17558 4100
rect 17773 4097 17785 4100
rect 17819 4128 17831 4131
rect 17862 4128 17868 4140
rect 17819 4100 17868 4128
rect 17819 4097 17831 4100
rect 17773 4091 17831 4097
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 19058 4128 19064 4140
rect 19019 4100 19064 4128
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 19150 4088 19156 4140
rect 19208 4128 19214 4140
rect 20073 4131 20131 4137
rect 19208 4100 19253 4128
rect 19208 4088 19214 4100
rect 20073 4097 20085 4131
rect 20119 4128 20131 4131
rect 20438 4128 20444 4140
rect 20119 4100 20444 4128
rect 20119 4097 20131 4100
rect 20073 4091 20131 4097
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 20993 4131 21051 4137
rect 20993 4097 21005 4131
rect 21039 4128 21051 4131
rect 21082 4128 21088 4140
rect 21039 4100 21088 4128
rect 21039 4097 21051 4100
rect 20993 4091 21051 4097
rect 21082 4088 21088 4100
rect 21140 4088 21146 4140
rect 22002 4128 22008 4140
rect 21963 4100 22008 4128
rect 22002 4088 22008 4100
rect 22060 4088 22066 4140
rect 22278 4137 22284 4140
rect 22272 4091 22284 4137
rect 22336 4128 22342 4140
rect 23934 4128 23940 4140
rect 22336 4100 22372 4128
rect 23895 4100 23940 4128
rect 22278 4088 22284 4091
rect 22336 4088 22342 4100
rect 23934 4088 23940 4100
rect 23992 4088 23998 4140
rect 25777 4131 25835 4137
rect 25777 4097 25789 4131
rect 25823 4128 25835 4131
rect 25823 4100 26096 4128
rect 25823 4097 25835 4100
rect 25777 4091 25835 4097
rect 17129 4063 17187 4069
rect 16163 4032 16620 4060
rect 16684 4032 17080 4060
rect 16163 4029 16175 4032
rect 16117 4023 16175 4029
rect 13722 3992 13728 4004
rect 9677 3955 9735 3961
rect 9784 3964 10548 3992
rect 10612 3964 13728 3992
rect 9030 3884 9036 3936
rect 9088 3924 9094 3936
rect 9784 3924 9812 3964
rect 9088 3896 9812 3924
rect 9861 3927 9919 3933
rect 9088 3884 9094 3896
rect 9861 3893 9873 3927
rect 9907 3924 9919 3927
rect 10134 3924 10140 3936
rect 9907 3896 10140 3924
rect 9907 3893 9919 3896
rect 9861 3887 9919 3893
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10520 3924 10548 3964
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 13814 3952 13820 4004
rect 13872 3992 13878 4004
rect 14277 3995 14335 4001
rect 14277 3992 14289 3995
rect 13872 3964 14289 3992
rect 13872 3952 13878 3964
rect 14277 3961 14289 3964
rect 14323 3961 14335 3995
rect 14277 3955 14335 3961
rect 14366 3952 14372 4004
rect 14424 3992 14430 4004
rect 15197 3995 15255 4001
rect 15197 3992 15209 3995
rect 14424 3964 15209 3992
rect 14424 3952 14430 3964
rect 15197 3961 15209 3964
rect 15243 3961 15255 3995
rect 15197 3955 15255 3961
rect 15381 3995 15439 4001
rect 15381 3961 15393 3995
rect 15427 3992 15439 3995
rect 16390 3992 16396 4004
rect 15427 3964 16396 3992
rect 15427 3961 15439 3964
rect 15381 3955 15439 3961
rect 16390 3952 16396 3964
rect 16448 3952 16454 4004
rect 16592 3992 16620 4032
rect 16666 3992 16672 4004
rect 16592 3964 16672 3992
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 17052 3992 17080 4032
rect 17129 4029 17141 4063
rect 17175 4060 17187 4063
rect 17310 4060 17316 4072
rect 17175 4032 17316 4060
rect 17175 4029 17187 4032
rect 17129 4023 17187 4029
rect 17310 4020 17316 4032
rect 17368 4020 17374 4072
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4060 18107 4063
rect 18414 4060 18420 4072
rect 18095 4032 18420 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18414 4020 18420 4032
rect 18472 4020 18478 4072
rect 18690 4020 18696 4072
rect 18748 4020 18754 4072
rect 18877 4063 18935 4069
rect 18877 4029 18889 4063
rect 18923 4029 18935 4063
rect 18877 4023 18935 4029
rect 18969 4063 19027 4069
rect 18969 4029 18981 4063
rect 19015 4029 19027 4063
rect 20162 4060 20168 4072
rect 18969 4023 19027 4029
rect 19260 4032 20168 4060
rect 18708 3992 18736 4020
rect 17052 3964 18736 3992
rect 13078 3924 13084 3936
rect 10520 3896 13084 3924
rect 13078 3884 13084 3896
rect 13136 3884 13142 3936
rect 13262 3884 13268 3936
rect 13320 3924 13326 3936
rect 13449 3927 13507 3933
rect 13449 3924 13461 3927
rect 13320 3896 13461 3924
rect 13320 3884 13326 3896
rect 13449 3893 13461 3896
rect 13495 3924 13507 3927
rect 14090 3924 14096 3936
rect 13495 3896 14096 3924
rect 13495 3893 13507 3896
rect 13449 3887 13507 3893
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 14461 3927 14519 3933
rect 14461 3893 14473 3927
rect 14507 3924 14519 3927
rect 17402 3924 17408 3936
rect 14507 3896 17408 3924
rect 14507 3893 14519 3896
rect 14461 3887 14519 3893
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 18690 3924 18696 3936
rect 18651 3896 18696 3924
rect 18690 3884 18696 3896
rect 18748 3884 18754 3936
rect 18892 3924 18920 4023
rect 18984 3992 19012 4023
rect 19260 3992 19288 4032
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 20349 4063 20407 4069
rect 20349 4029 20361 4063
rect 20395 4060 20407 4063
rect 20622 4060 20628 4072
rect 20395 4032 20628 4060
rect 20395 4029 20407 4032
rect 20349 4023 20407 4029
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 21269 4063 21327 4069
rect 21269 4029 21281 4063
rect 21315 4029 21327 4063
rect 21269 4023 21327 4029
rect 18984 3964 19288 3992
rect 18966 3924 18972 3936
rect 18892 3896 18972 3924
rect 18966 3884 18972 3896
rect 19024 3884 19030 3936
rect 19702 3924 19708 3936
rect 19663 3896 19708 3924
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 21284 3924 21312 4023
rect 25498 4020 25504 4072
rect 25556 4060 25562 4072
rect 25961 4063 26019 4069
rect 25961 4060 25973 4063
rect 25556 4032 25973 4060
rect 25556 4020 25562 4032
rect 25961 4029 25973 4032
rect 26007 4029 26019 4063
rect 26068 4060 26096 4100
rect 26418 4088 26424 4140
rect 26476 4128 26482 4140
rect 26476 4100 27752 4128
rect 26476 4088 26482 4100
rect 26878 4060 26884 4072
rect 26068 4032 26884 4060
rect 25961 4023 26019 4029
rect 26878 4020 26884 4032
rect 26936 4020 26942 4072
rect 26970 4020 26976 4072
rect 27028 4060 27034 4072
rect 27724 4069 27752 4100
rect 28534 4088 28540 4140
rect 28592 4128 28598 4140
rect 28629 4131 28687 4137
rect 28629 4128 28641 4131
rect 28592 4100 28641 4128
rect 28592 4088 28598 4100
rect 28629 4097 28641 4100
rect 28675 4097 28687 4131
rect 28629 4091 28687 4097
rect 28718 4088 28724 4140
rect 28776 4128 28782 4140
rect 28776 4100 29868 4128
rect 28776 4088 28782 4100
rect 27617 4063 27675 4069
rect 27617 4060 27629 4063
rect 27028 4032 27629 4060
rect 27028 4020 27034 4032
rect 27617 4029 27629 4032
rect 27663 4029 27675 4063
rect 27617 4023 27675 4029
rect 27709 4063 27767 4069
rect 27709 4029 27721 4063
rect 27755 4029 27767 4063
rect 29730 4060 29736 4072
rect 29691 4032 29736 4060
rect 27709 4023 27767 4029
rect 29730 4020 29736 4032
rect 29788 4020 29794 4072
rect 29840 4069 29868 4100
rect 30006 4088 30012 4140
rect 30064 4128 30070 4140
rect 30668 4128 30696 4168
rect 30064 4100 30696 4128
rect 31573 4131 31631 4137
rect 30064 4088 30070 4100
rect 31573 4097 31585 4131
rect 31619 4097 31631 4131
rect 31573 4091 31631 4097
rect 29825 4063 29883 4069
rect 29825 4029 29837 4063
rect 29871 4029 29883 4063
rect 29825 4023 29883 4029
rect 24946 3952 24952 4004
rect 25004 3992 25010 4004
rect 31202 3992 31208 4004
rect 25004 3964 31208 3992
rect 25004 3952 25010 3964
rect 31202 3952 31208 3964
rect 31260 3952 31266 4004
rect 31588 3992 31616 4091
rect 31680 4060 31708 4168
rect 32030 4156 32036 4208
rect 32088 4196 32094 4208
rect 32401 4199 32459 4205
rect 32401 4196 32413 4199
rect 32088 4168 32413 4196
rect 32088 4156 32094 4168
rect 32401 4165 32413 4168
rect 32447 4165 32459 4199
rect 32401 4159 32459 4165
rect 33410 4156 33416 4208
rect 33468 4196 33474 4208
rect 33781 4199 33839 4205
rect 33468 4168 33732 4196
rect 33468 4156 33474 4168
rect 31754 4088 31760 4140
rect 31812 4128 31818 4140
rect 32950 4128 32956 4140
rect 31812 4100 32956 4128
rect 31812 4088 31818 4100
rect 32950 4088 32956 4100
rect 33008 4088 33014 4140
rect 33594 4128 33600 4140
rect 33555 4100 33600 4128
rect 33594 4088 33600 4100
rect 33652 4088 33658 4140
rect 33704 4128 33732 4168
rect 33781 4165 33793 4199
rect 33827 4196 33839 4199
rect 35069 4199 35127 4205
rect 35069 4196 35081 4199
rect 33827 4168 35081 4196
rect 33827 4165 33839 4168
rect 33781 4159 33839 4165
rect 35069 4165 35081 4168
rect 35115 4196 35127 4199
rect 36906 4196 36912 4208
rect 35115 4168 36912 4196
rect 35115 4165 35127 4168
rect 35069 4159 35127 4165
rect 36906 4156 36912 4168
rect 36964 4156 36970 4208
rect 37182 4156 37188 4208
rect 37240 4196 37246 4208
rect 38473 4199 38531 4205
rect 37240 4168 38424 4196
rect 37240 4156 37246 4168
rect 33865 4131 33923 4137
rect 33865 4128 33877 4131
rect 33704 4100 33877 4128
rect 33865 4097 33877 4100
rect 33911 4097 33923 4131
rect 33989 4131 34047 4137
rect 33989 4128 34001 4131
rect 33865 4091 33923 4097
rect 33980 4097 34001 4128
rect 34035 4097 34047 4131
rect 33980 4091 34047 4097
rect 34701 4131 34759 4137
rect 34701 4097 34713 4131
rect 34747 4128 34759 4131
rect 35618 4128 35624 4140
rect 34747 4100 35624 4128
rect 34747 4097 34759 4100
rect 34701 4091 34759 4097
rect 33980 4060 34008 4091
rect 35618 4088 35624 4100
rect 35676 4088 35682 4140
rect 35710 4088 35716 4140
rect 35768 4128 35774 4140
rect 35805 4131 35863 4137
rect 35805 4128 35817 4131
rect 35768 4100 35817 4128
rect 35768 4088 35774 4100
rect 35805 4097 35817 4100
rect 35851 4097 35863 4131
rect 35805 4091 35863 4097
rect 35989 4131 36047 4137
rect 35989 4097 36001 4131
rect 36035 4097 36047 4131
rect 35989 4091 36047 4097
rect 36173 4131 36231 4137
rect 36173 4097 36185 4131
rect 36219 4097 36231 4131
rect 36173 4091 36231 4097
rect 31680 4032 34008 4060
rect 34149 3995 34207 4001
rect 31588 3964 33364 3992
rect 23014 3924 23020 3936
rect 21284 3896 23020 3924
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 23198 3884 23204 3936
rect 23256 3924 23262 3936
rect 25406 3924 25412 3936
rect 23256 3896 25412 3924
rect 23256 3884 23262 3896
rect 25406 3884 25412 3896
rect 25464 3884 25470 3936
rect 27154 3924 27160 3936
rect 27115 3896 27160 3924
rect 27154 3884 27160 3896
rect 27212 3884 27218 3936
rect 28534 3884 28540 3936
rect 28592 3924 28598 3936
rect 28813 3927 28871 3933
rect 28813 3924 28825 3927
rect 28592 3896 28825 3924
rect 28592 3884 28598 3896
rect 28813 3893 28825 3896
rect 28859 3893 28871 3927
rect 29270 3924 29276 3936
rect 29231 3896 29276 3924
rect 28813 3887 28871 3893
rect 29270 3884 29276 3896
rect 29328 3884 29334 3936
rect 30282 3884 30288 3936
rect 30340 3924 30346 3936
rect 30653 3927 30711 3933
rect 30653 3924 30665 3927
rect 30340 3896 30665 3924
rect 30340 3884 30346 3896
rect 30653 3893 30665 3896
rect 30699 3893 30711 3927
rect 31662 3924 31668 3936
rect 31623 3896 31668 3924
rect 30653 3887 30711 3893
rect 31662 3884 31668 3896
rect 31720 3884 31726 3936
rect 32493 3927 32551 3933
rect 32493 3893 32505 3927
rect 32539 3924 32551 3927
rect 33226 3924 33232 3936
rect 32539 3896 33232 3924
rect 32539 3893 32551 3896
rect 32493 3887 32551 3893
rect 33226 3884 33232 3896
rect 33284 3884 33290 3936
rect 33336 3924 33364 3964
rect 34149 3961 34161 3995
rect 34195 3992 34207 3995
rect 36004 3992 36032 4091
rect 34195 3964 36032 3992
rect 36188 3992 36216 4091
rect 36262 4088 36268 4140
rect 36320 4128 36326 4140
rect 37461 4131 37519 4137
rect 36320 4100 36365 4128
rect 36320 4088 36326 4100
rect 37461 4097 37473 4131
rect 37507 4128 37519 4131
rect 37550 4128 37556 4140
rect 37507 4100 37556 4128
rect 37507 4097 37519 4100
rect 37461 4091 37519 4097
rect 37550 4088 37556 4100
rect 37608 4088 37614 4140
rect 38396 4128 38424 4168
rect 38473 4165 38485 4199
rect 38519 4196 38531 4199
rect 38562 4196 38568 4208
rect 38519 4168 38568 4196
rect 38519 4165 38531 4168
rect 38473 4159 38531 4165
rect 38562 4156 38568 4168
rect 38620 4156 38626 4208
rect 38746 4156 38752 4208
rect 38804 4196 38810 4208
rect 40681 4199 40739 4205
rect 40681 4196 40693 4199
rect 38804 4168 40693 4196
rect 38804 4156 38810 4168
rect 40681 4165 40693 4168
rect 40727 4165 40739 4199
rect 46198 4196 46204 4208
rect 40681 4159 40739 4165
rect 45572 4168 46204 4196
rect 39209 4131 39267 4137
rect 39209 4128 39221 4131
rect 38396 4100 39221 4128
rect 39209 4097 39221 4100
rect 39255 4097 39267 4131
rect 39942 4128 39948 4140
rect 39903 4100 39948 4128
rect 39209 4091 39267 4097
rect 36354 4020 36360 4072
rect 36412 4060 36418 4072
rect 37645 4063 37703 4069
rect 37645 4060 37657 4063
rect 36412 4032 37657 4060
rect 36412 4020 36418 4032
rect 37645 4029 37657 4032
rect 37691 4029 37703 4063
rect 37645 4023 37703 4029
rect 38194 4020 38200 4072
rect 38252 4060 38258 4072
rect 38654 4060 38660 4072
rect 38252 4032 38660 4060
rect 38252 4020 38258 4032
rect 38654 4020 38660 4032
rect 38712 4020 38718 4072
rect 38838 4020 38844 4072
rect 38896 4060 38902 4072
rect 39114 4060 39120 4072
rect 38896 4032 39120 4060
rect 38896 4020 38902 4032
rect 39114 4020 39120 4032
rect 39172 4020 39178 4072
rect 39224 4060 39252 4091
rect 39942 4088 39948 4100
rect 40000 4088 40006 4140
rect 41506 4088 41512 4140
rect 41564 4128 41570 4140
rect 41601 4131 41659 4137
rect 41601 4128 41613 4131
rect 41564 4100 41613 4128
rect 41564 4088 41570 4100
rect 41601 4097 41613 4100
rect 41647 4097 41659 4131
rect 41601 4091 41659 4097
rect 42518 4088 42524 4140
rect 42576 4128 42582 4140
rect 42613 4131 42671 4137
rect 42613 4128 42625 4131
rect 42576 4100 42625 4128
rect 42576 4088 42582 4100
rect 42613 4097 42625 4100
rect 42659 4097 42671 4131
rect 43254 4128 43260 4140
rect 43215 4100 43260 4128
rect 42613 4091 42671 4097
rect 43254 4088 43260 4100
rect 43312 4088 43318 4140
rect 43625 4131 43683 4137
rect 43625 4097 43637 4131
rect 43671 4097 43683 4131
rect 43625 4091 43683 4097
rect 43809 4131 43867 4137
rect 43809 4097 43821 4131
rect 43855 4128 43867 4131
rect 43898 4128 43904 4140
rect 43855 4100 43904 4128
rect 43855 4097 43867 4100
rect 43809 4091 43867 4097
rect 40126 4060 40132 4072
rect 39224 4032 40132 4060
rect 40126 4020 40132 4032
rect 40184 4020 40190 4072
rect 41782 4060 41788 4072
rect 41743 4032 41788 4060
rect 41782 4020 41788 4032
rect 41840 4020 41846 4072
rect 43349 4063 43407 4069
rect 43349 4029 43361 4063
rect 43395 4029 43407 4063
rect 43640 4060 43668 4091
rect 43898 4088 43904 4100
rect 43956 4128 43962 4140
rect 45281 4131 45339 4137
rect 45281 4128 45293 4131
rect 43956 4100 45293 4128
rect 43956 4088 43962 4100
rect 45281 4097 45293 4100
rect 45327 4097 45339 4131
rect 45281 4091 45339 4097
rect 45373 4131 45431 4137
rect 45373 4097 45385 4131
rect 45419 4128 45431 4131
rect 45572 4128 45600 4168
rect 46198 4156 46204 4168
rect 46256 4156 46262 4208
rect 46290 4156 46296 4208
rect 46348 4196 46354 4208
rect 46842 4196 46848 4208
rect 46348 4168 46704 4196
rect 46803 4168 46848 4196
rect 46348 4156 46354 4168
rect 45419 4100 45600 4128
rect 45419 4097 45431 4100
rect 45373 4091 45431 4097
rect 45646 4088 45652 4140
rect 45704 4128 45710 4140
rect 45925 4131 45983 4137
rect 45704 4100 45749 4128
rect 45704 4088 45710 4100
rect 45925 4097 45937 4131
rect 45971 4097 45983 4131
rect 45925 4091 45983 4097
rect 46109 4131 46167 4137
rect 46109 4097 46121 4131
rect 46155 4128 46167 4131
rect 46676 4128 46704 4168
rect 46842 4156 46848 4168
rect 46900 4156 46906 4208
rect 47026 4156 47032 4208
rect 47084 4196 47090 4208
rect 48593 4199 48651 4205
rect 48593 4196 48605 4199
rect 47084 4168 48605 4196
rect 47084 4156 47090 4168
rect 48593 4165 48605 4168
rect 48639 4165 48651 4199
rect 48593 4159 48651 4165
rect 47857 4131 47915 4137
rect 47857 4128 47869 4131
rect 46155 4100 46612 4128
rect 46676 4100 47869 4128
rect 46155 4097 46167 4100
rect 46109 4091 46167 4097
rect 45186 4060 45192 4072
rect 43640 4032 45192 4060
rect 43349 4023 43407 4029
rect 43070 3992 43076 4004
rect 36188 3964 43076 3992
rect 34195 3961 34207 3964
rect 34149 3955 34207 3961
rect 43070 3952 43076 3964
rect 43128 3952 43134 4004
rect 43364 3992 43392 4023
rect 45186 4020 45192 4032
rect 45244 4020 45250 4072
rect 45940 4060 45968 4091
rect 46198 4060 46204 4072
rect 45940 4032 46204 4060
rect 46198 4020 46204 4032
rect 46256 4020 46262 4072
rect 46382 3992 46388 4004
rect 43364 3964 46388 3992
rect 46382 3952 46388 3964
rect 46440 3952 46446 4004
rect 46584 3992 46612 4100
rect 47857 4097 47869 4100
rect 47903 4097 47915 4131
rect 55398 4128 55404 4140
rect 55359 4100 55404 4128
rect 47857 4091 47915 4097
rect 55398 4088 55404 4100
rect 55456 4088 55462 4140
rect 55582 4128 55588 4140
rect 55543 4100 55588 4128
rect 55582 4088 55588 4100
rect 55640 4088 55646 4140
rect 56301 4131 56359 4137
rect 56301 4128 56313 4131
rect 55876 4100 56313 4128
rect 47670 4020 47676 4072
rect 47728 4060 47734 4072
rect 48777 4063 48835 4069
rect 48777 4060 48789 4063
rect 47728 4032 48789 4060
rect 47728 4020 47734 4032
rect 48777 4029 48789 4032
rect 48823 4029 48835 4063
rect 48777 4023 48835 4029
rect 55493 4063 55551 4069
rect 55493 4029 55505 4063
rect 55539 4060 55551 4063
rect 55876 4060 55904 4100
rect 56301 4097 56313 4100
rect 56347 4097 56359 4131
rect 58066 4128 58072 4140
rect 58027 4100 58072 4128
rect 56301 4091 56359 4097
rect 58066 4088 58072 4100
rect 58124 4088 58130 4140
rect 55539 4032 55904 4060
rect 56045 4063 56103 4069
rect 55539 4029 55551 4032
rect 55493 4023 55551 4029
rect 56045 4029 56057 4063
rect 56091 4029 56103 4063
rect 56045 4023 56103 4029
rect 53926 3992 53932 4004
rect 46584 3964 53932 3992
rect 53926 3952 53932 3964
rect 53984 3952 53990 4004
rect 34330 3924 34336 3936
rect 33336 3896 34336 3924
rect 34330 3884 34336 3896
rect 34388 3884 34394 3936
rect 36262 3884 36268 3936
rect 36320 3924 36326 3936
rect 37182 3924 37188 3936
rect 36320 3896 37188 3924
rect 36320 3884 36326 3896
rect 37182 3884 37188 3896
rect 37240 3884 37246 3936
rect 37458 3884 37464 3936
rect 37516 3924 37522 3936
rect 38565 3927 38623 3933
rect 38565 3924 38577 3927
rect 37516 3896 38577 3924
rect 37516 3884 37522 3896
rect 38565 3893 38577 3896
rect 38611 3893 38623 3927
rect 38565 3887 38623 3893
rect 38654 3884 38660 3936
rect 38712 3924 38718 3936
rect 39301 3927 39359 3933
rect 39301 3924 39313 3927
rect 38712 3896 39313 3924
rect 38712 3884 38718 3896
rect 39301 3893 39313 3896
rect 39347 3893 39359 3927
rect 39301 3887 39359 3893
rect 40037 3927 40095 3933
rect 40037 3893 40049 3927
rect 40083 3924 40095 3927
rect 40218 3924 40224 3936
rect 40083 3896 40224 3924
rect 40083 3893 40095 3896
rect 40037 3887 40095 3893
rect 40218 3884 40224 3896
rect 40276 3884 40282 3936
rect 40678 3884 40684 3936
rect 40736 3924 40742 3936
rect 40773 3927 40831 3933
rect 40773 3924 40785 3927
rect 40736 3896 40785 3924
rect 40736 3884 40742 3896
rect 40773 3893 40785 3896
rect 40819 3893 40831 3927
rect 40773 3887 40831 3893
rect 42242 3884 42248 3936
rect 42300 3924 42306 3936
rect 44913 3927 44971 3933
rect 44913 3924 44925 3927
rect 42300 3896 44925 3924
rect 42300 3884 42306 3896
rect 44913 3893 44925 3896
rect 44959 3893 44971 3927
rect 44913 3887 44971 3893
rect 46658 3884 46664 3936
rect 46716 3924 46722 3936
rect 46937 3927 46995 3933
rect 46937 3924 46949 3927
rect 46716 3896 46949 3924
rect 46716 3884 46722 3896
rect 46937 3893 46949 3896
rect 46983 3893 46995 3927
rect 46937 3887 46995 3893
rect 47854 3884 47860 3936
rect 47912 3924 47918 3936
rect 47949 3927 48007 3933
rect 47949 3924 47961 3927
rect 47912 3896 47961 3924
rect 47912 3884 47918 3896
rect 47949 3893 47961 3896
rect 47995 3893 48007 3927
rect 56060 3924 56088 4023
rect 56686 3924 56692 3936
rect 56060 3896 56692 3924
rect 47949 3887 48007 3893
rect 56686 3884 56692 3896
rect 56744 3884 56750 3936
rect 57422 3924 57428 3936
rect 57383 3896 57428 3924
rect 57422 3884 57428 3896
rect 57480 3884 57486 3936
rect 58250 3924 58256 3936
rect 58211 3896 58256 3924
rect 58250 3884 58256 3896
rect 58308 3884 58314 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 7009 3723 7067 3729
rect 7009 3689 7021 3723
rect 7055 3720 7067 3723
rect 9398 3720 9404 3732
rect 7055 3692 9404 3720
rect 7055 3689 7067 3692
rect 7009 3683 7067 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 20070 3720 20076 3732
rect 12308 3692 20076 3720
rect 12308 3680 12314 3692
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 20162 3680 20168 3732
rect 20220 3720 20226 3732
rect 20809 3723 20867 3729
rect 20809 3720 20821 3723
rect 20220 3692 20821 3720
rect 20220 3680 20226 3692
rect 20809 3689 20821 3692
rect 20855 3689 20867 3723
rect 20809 3683 20867 3689
rect 22189 3723 22247 3729
rect 22189 3689 22201 3723
rect 22235 3720 22247 3723
rect 22462 3720 22468 3732
rect 22235 3692 22468 3720
rect 22235 3689 22247 3692
rect 22189 3683 22247 3689
rect 22462 3680 22468 3692
rect 22520 3680 22526 3732
rect 33502 3720 33508 3732
rect 23584 3692 33508 3720
rect 6273 3655 6331 3661
rect 6273 3621 6285 3655
rect 6319 3652 6331 3655
rect 7466 3652 7472 3664
rect 6319 3624 7472 3652
rect 6319 3621 6331 3624
rect 6273 3615 6331 3621
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 7837 3655 7895 3661
rect 7837 3621 7849 3655
rect 7883 3652 7895 3655
rect 7926 3652 7932 3664
rect 7883 3624 7932 3652
rect 7883 3621 7895 3624
rect 7837 3615 7895 3621
rect 7926 3612 7932 3624
rect 7984 3612 7990 3664
rect 8662 3612 8668 3664
rect 8720 3652 8726 3664
rect 9677 3655 9735 3661
rect 9677 3652 9689 3655
rect 8720 3624 9689 3652
rect 8720 3612 8726 3624
rect 9677 3621 9689 3624
rect 9723 3621 9735 3655
rect 9677 3615 9735 3621
rect 10502 3612 10508 3664
rect 10560 3652 10566 3664
rect 11425 3655 11483 3661
rect 11425 3652 11437 3655
rect 10560 3624 11437 3652
rect 10560 3612 10566 3624
rect 11425 3621 11437 3624
rect 11471 3621 11483 3655
rect 12342 3652 12348 3664
rect 12303 3624 12348 3652
rect 11425 3615 11483 3621
rect 12342 3612 12348 3624
rect 12400 3612 12406 3664
rect 12434 3612 12440 3664
rect 12492 3652 12498 3664
rect 12529 3655 12587 3661
rect 12529 3652 12541 3655
rect 12492 3624 12541 3652
rect 12492 3612 12498 3624
rect 12529 3621 12541 3624
rect 12575 3621 12587 3655
rect 12529 3615 12587 3621
rect 13633 3655 13691 3661
rect 13633 3621 13645 3655
rect 13679 3652 13691 3655
rect 14458 3652 14464 3664
rect 13679 3624 14464 3652
rect 13679 3621 13691 3624
rect 13633 3615 13691 3621
rect 14458 3612 14464 3624
rect 14516 3612 14522 3664
rect 15010 3652 15016 3664
rect 14971 3624 15016 3652
rect 15010 3612 15016 3624
rect 15068 3612 15074 3664
rect 17402 3612 17408 3664
rect 17460 3652 17466 3664
rect 18874 3652 18880 3664
rect 17460 3624 18880 3652
rect 17460 3612 17466 3624
rect 18874 3612 18880 3624
rect 18932 3612 18938 3664
rect 19058 3612 19064 3664
rect 19116 3652 19122 3664
rect 19116 3624 19334 3652
rect 19116 3612 19122 3624
rect 9398 3584 9404 3596
rect 2746 3556 9404 3584
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 2746 3516 2774 3556
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 9858 3584 9864 3596
rect 9819 3556 9864 3584
rect 9858 3544 9864 3556
rect 9916 3544 9922 3596
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 10134 3584 10140 3596
rect 10008 3556 10053 3584
rect 10095 3556 10140 3584
rect 10008 3544 10014 3556
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 13262 3584 13268 3596
rect 13223 3556 13268 3584
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 13722 3584 13728 3596
rect 13683 3556 13728 3584
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 14737 3587 14795 3593
rect 14737 3553 14749 3587
rect 14783 3584 14795 3587
rect 14918 3584 14924 3596
rect 14783 3556 14924 3584
rect 14783 3553 14795 3556
rect 14737 3547 14795 3553
rect 14918 3544 14924 3556
rect 14976 3544 14982 3596
rect 15933 3587 15991 3593
rect 15933 3553 15945 3587
rect 15979 3584 15991 3587
rect 17126 3584 17132 3596
rect 15979 3556 17132 3584
rect 15979 3553 15991 3556
rect 15933 3547 15991 3553
rect 17126 3544 17132 3556
rect 17184 3544 17190 3596
rect 18693 3587 18751 3593
rect 18693 3553 18705 3587
rect 18739 3584 18751 3587
rect 18966 3584 18972 3596
rect 18739 3556 18972 3584
rect 18739 3553 18751 3556
rect 18693 3547 18751 3553
rect 18966 3544 18972 3556
rect 19024 3544 19030 3596
rect 19306 3584 19334 3624
rect 20438 3612 20444 3664
rect 20496 3652 20502 3664
rect 22005 3655 22063 3661
rect 22005 3652 22017 3655
rect 20496 3624 22017 3652
rect 20496 3612 20502 3624
rect 22005 3621 22017 3624
rect 22051 3621 22063 3655
rect 22005 3615 22063 3621
rect 19426 3584 19432 3596
rect 19306 3556 19432 3584
rect 19426 3544 19432 3556
rect 19484 3544 19490 3596
rect 21726 3584 21732 3596
rect 21687 3556 21732 3584
rect 21726 3544 21732 3556
rect 21784 3584 21790 3596
rect 23017 3587 23075 3593
rect 23017 3584 23029 3587
rect 21784 3556 23029 3584
rect 21784 3544 21790 3556
rect 23017 3553 23029 3556
rect 23063 3553 23075 3587
rect 23017 3547 23075 3553
rect 1627 3488 2774 3516
rect 6917 3519 6975 3525
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 6917 3485 6929 3519
rect 6963 3516 6975 3519
rect 8294 3516 8300 3528
rect 6963 3488 8300 3516
rect 6963 3485 6975 3488
rect 6917 3479 6975 3485
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 9306 3516 9312 3528
rect 8435 3488 9312 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3516 10103 3519
rect 10686 3516 10692 3528
rect 10091 3488 10692 3516
rect 10091 3485 10103 3488
rect 10045 3479 10103 3485
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 11974 3476 11980 3528
rect 12032 3516 12038 3528
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 12032 3488 12081 3516
rect 12032 3476 12038 3488
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 15657 3519 15715 3525
rect 15657 3485 15669 3519
rect 15703 3516 15715 3519
rect 16206 3516 16212 3528
rect 15703 3488 16212 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 16574 3516 16580 3528
rect 16535 3488 16580 3516
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 17497 3519 17555 3525
rect 17497 3485 17509 3519
rect 17543 3516 17555 3519
rect 17586 3516 17592 3528
rect 17543 3488 17592 3516
rect 17543 3485 17555 3488
rect 17497 3479 17555 3485
rect 1854 3448 1860 3460
rect 1815 3420 1860 3448
rect 1854 3408 1860 3420
rect 1912 3408 1918 3460
rect 5902 3408 5908 3460
rect 5960 3448 5966 3460
rect 6089 3451 6147 3457
rect 6089 3448 6101 3451
rect 5960 3420 6101 3448
rect 5960 3408 5966 3420
rect 6089 3417 6101 3420
rect 6135 3417 6147 3451
rect 6089 3411 6147 3417
rect 7653 3451 7711 3457
rect 7653 3417 7665 3451
rect 7699 3448 7711 3451
rect 7699 3420 9628 3448
rect 7699 3417 7711 3420
rect 7653 3411 7711 3417
rect 8481 3383 8539 3389
rect 8481 3349 8493 3383
rect 8527 3380 8539 3383
rect 8846 3380 8852 3392
rect 8527 3352 8852 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 9600 3380 9628 3420
rect 11054 3408 11060 3460
rect 11112 3448 11118 3460
rect 11149 3451 11207 3457
rect 11149 3448 11161 3451
rect 11112 3420 11161 3448
rect 11112 3408 11118 3420
rect 11149 3417 11161 3420
rect 11195 3417 11207 3451
rect 16868 3448 16896 3479
rect 17586 3476 17592 3488
rect 17644 3476 17650 3528
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 18472 3488 18517 3516
rect 18472 3476 18478 3488
rect 19242 3476 19248 3528
rect 19300 3516 19306 3528
rect 19518 3516 19524 3528
rect 19300 3488 19524 3516
rect 19300 3476 19306 3488
rect 19518 3476 19524 3488
rect 19576 3476 19582 3528
rect 19702 3525 19708 3528
rect 19696 3516 19708 3525
rect 19663 3488 19708 3516
rect 19696 3479 19708 3488
rect 19702 3476 19708 3479
rect 19760 3476 19766 3528
rect 20070 3476 20076 3528
rect 20128 3516 20134 3528
rect 23584 3525 23612 3692
rect 33502 3680 33508 3692
rect 33560 3680 33566 3732
rect 34422 3680 34428 3732
rect 34480 3720 34486 3732
rect 34480 3692 35296 3720
rect 34480 3680 34486 3692
rect 24578 3652 24584 3664
rect 24539 3624 24584 3652
rect 24578 3612 24584 3624
rect 24636 3612 24642 3664
rect 26970 3612 26976 3664
rect 27028 3652 27034 3664
rect 27157 3655 27215 3661
rect 27157 3652 27169 3655
rect 27028 3624 27169 3652
rect 27028 3612 27034 3624
rect 27157 3621 27169 3624
rect 27203 3621 27215 3655
rect 29822 3652 29828 3664
rect 27157 3615 27215 3621
rect 27632 3624 29828 3652
rect 24854 3584 24860 3596
rect 23768 3556 24860 3584
rect 23569 3519 23627 3525
rect 20128 3488 23520 3516
rect 20128 3476 20134 3488
rect 17773 3451 17831 3457
rect 16868 3420 17724 3448
rect 11149 3411 11207 3417
rect 9766 3380 9772 3392
rect 9600 3352 9772 3380
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 11606 3380 11612 3392
rect 11567 3352 11612 3380
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 11882 3340 11888 3392
rect 11940 3380 11946 3392
rect 14458 3380 14464 3392
rect 11940 3352 14464 3380
rect 11940 3340 11946 3352
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 15197 3383 15255 3389
rect 15197 3349 15209 3383
rect 15243 3380 15255 3383
rect 17402 3380 17408 3392
rect 15243 3352 17408 3380
rect 15243 3349 15255 3352
rect 15197 3343 15255 3349
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 17696 3380 17724 3420
rect 17773 3417 17785 3451
rect 17819 3448 17831 3451
rect 18966 3448 18972 3460
rect 17819 3420 18972 3448
rect 17819 3417 17831 3420
rect 17773 3411 17831 3417
rect 18966 3408 18972 3420
rect 19024 3408 19030 3460
rect 19978 3448 19984 3460
rect 19058 3420 19984 3448
rect 19058 3380 19086 3420
rect 19978 3408 19984 3420
rect 20036 3408 20042 3460
rect 22741 3451 22799 3457
rect 22741 3417 22753 3451
rect 22787 3448 22799 3451
rect 23492 3448 23520 3488
rect 23569 3485 23581 3519
rect 23615 3485 23627 3519
rect 23569 3479 23627 3485
rect 23768 3448 23796 3556
rect 24854 3544 24860 3556
rect 24912 3584 24918 3596
rect 25041 3587 25099 3593
rect 25041 3584 25053 3587
rect 24912 3556 25053 3584
rect 24912 3544 24918 3556
rect 25041 3553 25053 3556
rect 25087 3553 25099 3587
rect 25041 3547 25099 3553
rect 25130 3544 25136 3596
rect 25188 3584 25194 3596
rect 25188 3556 25233 3584
rect 25188 3544 25194 3556
rect 26878 3544 26884 3596
rect 26936 3584 26942 3596
rect 27632 3584 27660 3624
rect 29822 3612 29828 3624
rect 29880 3612 29886 3664
rect 26936 3556 27660 3584
rect 27709 3587 27767 3593
rect 26936 3544 26942 3556
rect 27709 3553 27721 3587
rect 27755 3584 27767 3587
rect 29362 3584 29368 3596
rect 27755 3556 29368 3584
rect 27755 3553 27767 3556
rect 27709 3547 27767 3553
rect 29362 3544 29368 3556
rect 29420 3544 29426 3596
rect 30926 3544 30932 3596
rect 30984 3584 30990 3596
rect 32033 3587 32091 3593
rect 32033 3584 32045 3587
rect 30984 3556 32045 3584
rect 30984 3544 30990 3556
rect 32033 3553 32045 3556
rect 32079 3553 32091 3587
rect 32033 3547 32091 3553
rect 33502 3544 33508 3596
rect 33560 3584 33566 3596
rect 35069 3587 35127 3593
rect 35069 3584 35081 3587
rect 33560 3556 35081 3584
rect 33560 3544 33566 3556
rect 35069 3553 35081 3556
rect 35115 3553 35127 3587
rect 35069 3547 35127 3553
rect 23934 3476 23940 3528
rect 23992 3516 23998 3528
rect 25777 3519 25835 3525
rect 25777 3516 25789 3519
rect 23992 3488 25789 3516
rect 23992 3476 23998 3488
rect 25777 3485 25789 3488
rect 25823 3485 25835 3519
rect 25777 3479 25835 3485
rect 26044 3519 26102 3525
rect 26044 3485 26056 3519
rect 26090 3516 26102 3519
rect 27154 3516 27160 3528
rect 26090 3488 27160 3516
rect 26090 3485 26102 3488
rect 26044 3479 26102 3485
rect 27154 3476 27160 3488
rect 27212 3476 27218 3528
rect 28166 3476 28172 3528
rect 28224 3516 28230 3528
rect 28534 3516 28540 3528
rect 28224 3488 28540 3516
rect 28224 3476 28230 3488
rect 28534 3476 28540 3488
rect 28592 3476 28598 3528
rect 28675 3519 28733 3525
rect 28675 3485 28687 3519
rect 28721 3516 28733 3519
rect 29730 3516 29736 3528
rect 28721 3488 29736 3516
rect 28721 3485 28733 3488
rect 28675 3479 28733 3485
rect 29730 3476 29736 3488
rect 29788 3476 29794 3528
rect 30282 3516 30288 3528
rect 30243 3488 30288 3516
rect 30282 3476 30288 3488
rect 30340 3476 30346 3528
rect 31938 3516 31944 3528
rect 30668 3488 31944 3516
rect 22787 3420 23428 3448
rect 23492 3420 23796 3448
rect 23845 3451 23903 3457
rect 22787 3417 22799 3420
rect 22741 3411 22799 3417
rect 17696 3352 19086 3380
rect 19150 3340 19156 3392
rect 19208 3380 19214 3392
rect 20806 3380 20812 3392
rect 19208 3352 20812 3380
rect 19208 3340 19214 3352
rect 20806 3340 20812 3352
rect 20864 3340 20870 3392
rect 23400 3380 23428 3420
rect 23845 3417 23857 3451
rect 23891 3448 23903 3451
rect 24670 3448 24676 3460
rect 23891 3420 24676 3448
rect 23891 3417 23903 3420
rect 23845 3411 23903 3417
rect 24670 3408 24676 3420
rect 24728 3408 24734 3460
rect 28350 3448 28356 3460
rect 24872 3420 27752 3448
rect 28311 3420 28356 3448
rect 24872 3380 24900 3420
rect 23400 3352 24900 3380
rect 24949 3383 25007 3389
rect 24949 3349 24961 3383
rect 24995 3380 25007 3383
rect 27614 3380 27620 3392
rect 24995 3352 27620 3380
rect 24995 3349 25007 3352
rect 24949 3343 25007 3349
rect 27614 3340 27620 3352
rect 27672 3340 27678 3392
rect 27724 3380 27752 3420
rect 28350 3408 28356 3420
rect 28408 3408 28414 3460
rect 28902 3448 28908 3460
rect 28863 3420 28908 3448
rect 28902 3408 28908 3420
rect 28960 3408 28966 3460
rect 30190 3408 30196 3460
rect 30248 3448 30254 3460
rect 30561 3451 30619 3457
rect 30561 3448 30573 3451
rect 30248 3420 30573 3448
rect 30248 3408 30254 3420
rect 30561 3417 30573 3420
rect 30607 3417 30619 3451
rect 30561 3411 30619 3417
rect 28721 3383 28779 3389
rect 28721 3380 28733 3383
rect 27724 3352 28733 3380
rect 28721 3349 28733 3352
rect 28767 3380 28779 3383
rect 30668 3380 30696 3488
rect 31938 3476 31944 3488
rect 31996 3476 32002 3528
rect 32306 3525 32312 3528
rect 32300 3516 32312 3525
rect 32267 3488 32312 3516
rect 32300 3479 32312 3488
rect 32306 3476 32312 3479
rect 32364 3476 32370 3528
rect 32582 3476 32588 3528
rect 32640 3516 32646 3528
rect 34057 3519 34115 3525
rect 34057 3516 34069 3519
rect 32640 3488 34069 3516
rect 32640 3476 32646 3488
rect 34057 3485 34069 3488
rect 34103 3516 34115 3519
rect 34514 3516 34520 3528
rect 34103 3488 34520 3516
rect 34103 3485 34115 3488
rect 34057 3479 34115 3485
rect 34514 3476 34520 3488
rect 34572 3476 34578 3528
rect 34698 3476 34704 3528
rect 34756 3516 34762 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34756 3488 34897 3516
rect 34756 3476 34762 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 35268 3516 35296 3692
rect 37550 3680 37556 3732
rect 37608 3720 37614 3732
rect 40221 3723 40279 3729
rect 40221 3720 40233 3723
rect 37608 3692 40233 3720
rect 37608 3680 37614 3692
rect 40221 3689 40233 3692
rect 40267 3689 40279 3723
rect 40221 3683 40279 3689
rect 44177 3723 44235 3729
rect 44177 3689 44189 3723
rect 44223 3720 44235 3723
rect 44266 3720 44272 3732
rect 44223 3692 44272 3720
rect 44223 3689 44235 3692
rect 44177 3683 44235 3689
rect 44266 3680 44272 3692
rect 44324 3680 44330 3732
rect 44450 3680 44456 3732
rect 44508 3720 44514 3732
rect 46106 3720 46112 3732
rect 44508 3692 46112 3720
rect 44508 3680 44514 3692
rect 46106 3680 46112 3692
rect 46164 3680 46170 3732
rect 47578 3720 47584 3732
rect 46676 3692 47584 3720
rect 38657 3655 38715 3661
rect 38657 3621 38669 3655
rect 38703 3652 38715 3655
rect 39390 3652 39396 3664
rect 38703 3624 39396 3652
rect 38703 3621 38715 3624
rect 38657 3615 38715 3621
rect 39390 3612 39396 3624
rect 39448 3612 39454 3664
rect 39485 3655 39543 3661
rect 39485 3621 39497 3655
rect 39531 3652 39543 3655
rect 39666 3652 39672 3664
rect 39531 3624 39672 3652
rect 39531 3621 39543 3624
rect 39485 3615 39543 3621
rect 39666 3612 39672 3624
rect 39724 3612 39730 3664
rect 40402 3612 40408 3664
rect 40460 3652 40466 3664
rect 40460 3624 42564 3652
rect 40460 3612 40466 3624
rect 35986 3584 35992 3596
rect 35947 3556 35992 3584
rect 35986 3544 35992 3556
rect 36044 3544 36050 3596
rect 37642 3544 37648 3596
rect 37700 3584 37706 3596
rect 38930 3584 38936 3596
rect 37700 3556 38936 3584
rect 37700 3544 37706 3556
rect 38930 3544 38936 3556
rect 38988 3544 38994 3596
rect 39224 3556 40908 3584
rect 35805 3519 35863 3525
rect 35805 3516 35817 3519
rect 35268 3488 35817 3516
rect 34885 3479 34943 3485
rect 35805 3485 35817 3488
rect 35851 3485 35863 3519
rect 35805 3479 35863 3485
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 36725 3519 36783 3525
rect 36725 3516 36737 3519
rect 35952 3488 36737 3516
rect 35952 3476 35958 3488
rect 36725 3485 36737 3488
rect 36771 3485 36783 3519
rect 36725 3479 36783 3485
rect 36906 3476 36912 3528
rect 36964 3516 36970 3528
rect 38102 3516 38108 3528
rect 36964 3488 37964 3516
rect 38063 3488 38108 3516
rect 36964 3476 36970 3488
rect 31389 3451 31447 3457
rect 31389 3417 31401 3451
rect 31435 3448 31447 3451
rect 31435 3420 31754 3448
rect 31435 3417 31447 3420
rect 31389 3411 31447 3417
rect 31478 3380 31484 3392
rect 28767 3352 30696 3380
rect 31439 3352 31484 3380
rect 28767 3349 28779 3352
rect 28721 3343 28779 3349
rect 31478 3340 31484 3352
rect 31536 3340 31542 3392
rect 31726 3380 31754 3420
rect 32030 3408 32036 3460
rect 32088 3448 32094 3460
rect 33962 3448 33968 3460
rect 32088 3420 33968 3448
rect 32088 3408 32094 3420
rect 33962 3408 33968 3420
rect 34020 3408 34026 3460
rect 34241 3451 34299 3457
rect 34241 3417 34253 3451
rect 34287 3448 34299 3451
rect 34790 3448 34796 3460
rect 34287 3420 34796 3448
rect 34287 3417 34299 3420
rect 34241 3411 34299 3417
rect 34790 3408 34796 3420
rect 34848 3408 34854 3460
rect 37001 3451 37059 3457
rect 37001 3417 37013 3451
rect 37047 3417 37059 3451
rect 37936 3448 37964 3488
rect 38102 3476 38108 3488
rect 38160 3476 38166 3528
rect 38478 3519 38536 3525
rect 38478 3516 38490 3519
rect 38212 3488 38490 3516
rect 38212 3448 38240 3488
rect 38478 3485 38490 3488
rect 38524 3516 38536 3519
rect 39224 3516 39252 3556
rect 38524 3488 39252 3516
rect 39301 3519 39359 3525
rect 38524 3485 38536 3488
rect 38478 3479 38536 3485
rect 39301 3485 39313 3519
rect 39347 3516 39359 3519
rect 39482 3516 39488 3528
rect 39347 3488 39488 3516
rect 39347 3485 39359 3488
rect 39301 3479 39359 3485
rect 39482 3476 39488 3488
rect 39540 3476 39546 3528
rect 40126 3516 40132 3528
rect 40087 3488 40132 3516
rect 40126 3476 40132 3488
rect 40184 3476 40190 3528
rect 37936 3420 38240 3448
rect 38289 3451 38347 3457
rect 37001 3411 37059 3417
rect 38289 3417 38301 3451
rect 38335 3417 38347 3451
rect 38289 3411 38347 3417
rect 38381 3451 38439 3457
rect 38381 3417 38393 3451
rect 38427 3448 38439 3451
rect 38838 3448 38844 3460
rect 38427 3420 38844 3448
rect 38427 3417 38439 3420
rect 38381 3411 38439 3417
rect 32214 3380 32220 3392
rect 31726 3352 32220 3380
rect 32214 3340 32220 3352
rect 32272 3380 32278 3392
rect 33042 3380 33048 3392
rect 32272 3352 33048 3380
rect 32272 3340 32278 3352
rect 33042 3340 33048 3352
rect 33100 3340 33106 3392
rect 33410 3380 33416 3392
rect 33371 3352 33416 3380
rect 33410 3340 33416 3352
rect 33468 3380 33474 3392
rect 33686 3380 33692 3392
rect 33468 3352 33692 3380
rect 33468 3340 33474 3352
rect 33686 3340 33692 3352
rect 33744 3340 33750 3392
rect 34698 3340 34704 3392
rect 34756 3380 34762 3392
rect 37016 3380 37044 3411
rect 34756 3352 37044 3380
rect 34756 3340 34762 3352
rect 37182 3340 37188 3392
rect 37240 3380 37246 3392
rect 38304 3380 38332 3411
rect 38838 3408 38844 3420
rect 38896 3408 38902 3460
rect 40880 3448 40908 3556
rect 41046 3544 41052 3596
rect 41104 3584 41110 3596
rect 41141 3587 41199 3593
rect 41141 3584 41153 3587
rect 41104 3556 41153 3584
rect 41104 3544 41110 3556
rect 41141 3553 41153 3556
rect 41187 3553 41199 3587
rect 41874 3584 41880 3596
rect 41835 3556 41880 3584
rect 41141 3547 41199 3553
rect 41874 3544 41880 3556
rect 41932 3544 41938 3596
rect 40957 3519 41015 3525
rect 40957 3485 40969 3519
rect 41003 3516 41015 3519
rect 41782 3516 41788 3528
rect 41003 3488 41788 3516
rect 41003 3485 41015 3488
rect 40957 3479 41015 3485
rect 41782 3476 41788 3488
rect 41840 3476 41846 3528
rect 42536 3525 42564 3624
rect 42610 3544 42616 3596
rect 42668 3584 42674 3596
rect 43898 3584 43904 3596
rect 42668 3556 42713 3584
rect 42996 3556 43904 3584
rect 42668 3544 42674 3556
rect 42521 3519 42579 3525
rect 42521 3485 42533 3519
rect 42567 3485 42579 3519
rect 42886 3516 42892 3528
rect 42847 3488 42892 3516
rect 42521 3479 42579 3485
rect 42886 3476 42892 3488
rect 42944 3476 42950 3528
rect 42996 3525 43024 3556
rect 43898 3544 43904 3556
rect 43956 3584 43962 3596
rect 43956 3556 44041 3584
rect 43956 3544 43962 3556
rect 42981 3519 43039 3525
rect 42981 3485 42993 3519
rect 43027 3485 43039 3519
rect 42981 3479 43039 3485
rect 42996 3448 43024 3479
rect 43438 3476 43444 3528
rect 43496 3516 43502 3528
rect 43714 3525 43720 3528
rect 43533 3519 43591 3525
rect 43533 3516 43545 3519
rect 43496 3488 43545 3516
rect 43496 3476 43502 3488
rect 43533 3485 43545 3488
rect 43579 3485 43591 3519
rect 43533 3479 43591 3485
rect 43681 3519 43720 3525
rect 43681 3485 43693 3519
rect 43681 3479 43720 3485
rect 43714 3476 43720 3479
rect 43772 3476 43778 3528
rect 44013 3525 44041 3556
rect 44634 3544 44640 3596
rect 44692 3584 44698 3596
rect 45094 3584 45100 3596
rect 44692 3556 45100 3584
rect 44692 3544 44698 3556
rect 45094 3544 45100 3556
rect 45152 3544 45158 3596
rect 45554 3544 45560 3596
rect 45612 3544 45618 3596
rect 45830 3544 45836 3596
rect 45888 3584 45894 3596
rect 45888 3556 46152 3584
rect 45888 3544 45894 3556
rect 43998 3519 44056 3525
rect 43998 3485 44010 3519
rect 44044 3516 44056 3519
rect 44266 3516 44272 3528
rect 44044 3488 44272 3516
rect 44044 3485 44056 3488
rect 43998 3479 44056 3485
rect 44266 3476 44272 3488
rect 44324 3476 44330 3528
rect 45186 3516 45192 3528
rect 45147 3488 45192 3516
rect 45186 3476 45192 3488
rect 45244 3476 45250 3528
rect 45572 3516 45600 3544
rect 45649 3519 45707 3525
rect 45649 3516 45661 3519
rect 45480 3488 45661 3516
rect 40880 3420 43024 3448
rect 43346 3408 43352 3460
rect 43404 3448 43410 3460
rect 43809 3451 43867 3457
rect 43809 3448 43821 3451
rect 43404 3420 43821 3448
rect 43404 3408 43410 3420
rect 43809 3417 43821 3420
rect 43855 3417 43867 3451
rect 43809 3411 43867 3417
rect 43898 3408 43904 3460
rect 43956 3448 43962 3460
rect 44284 3448 44312 3476
rect 45480 3448 45508 3488
rect 45649 3485 45661 3488
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 45738 3476 45744 3528
rect 45796 3516 45802 3528
rect 46014 3516 46020 3528
rect 45796 3488 45841 3516
rect 45975 3488 46020 3516
rect 45796 3476 45802 3488
rect 46014 3476 46020 3488
rect 46072 3476 46078 3528
rect 43956 3420 44001 3448
rect 44284 3420 45508 3448
rect 46124 3448 46152 3556
rect 46198 3476 46204 3528
rect 46256 3516 46262 3528
rect 46293 3519 46351 3525
rect 46293 3516 46305 3519
rect 46256 3488 46305 3516
rect 46256 3476 46262 3488
rect 46293 3485 46305 3488
rect 46339 3485 46351 3519
rect 46293 3479 46351 3485
rect 46569 3519 46627 3525
rect 46569 3485 46581 3519
rect 46615 3516 46627 3519
rect 46676 3516 46704 3692
rect 47578 3680 47584 3692
rect 47636 3680 47642 3732
rect 48038 3720 48044 3732
rect 47999 3692 48044 3720
rect 48038 3680 48044 3692
rect 48096 3680 48102 3732
rect 49697 3723 49755 3729
rect 49697 3689 49709 3723
rect 49743 3720 49755 3723
rect 49878 3720 49884 3732
rect 49743 3692 49884 3720
rect 49743 3689 49755 3692
rect 49697 3683 49755 3689
rect 49878 3680 49884 3692
rect 49936 3680 49942 3732
rect 51258 3720 51264 3732
rect 51219 3692 51264 3720
rect 51258 3680 51264 3692
rect 51316 3680 51322 3732
rect 52730 3720 52736 3732
rect 52691 3692 52736 3720
rect 52730 3680 52736 3692
rect 52788 3680 52794 3732
rect 52914 3680 52920 3732
rect 52972 3720 52978 3732
rect 53469 3723 53527 3729
rect 53469 3720 53481 3723
rect 52972 3692 53481 3720
rect 52972 3680 52978 3692
rect 53469 3689 53481 3692
rect 53515 3689 53527 3723
rect 53469 3683 53527 3689
rect 53558 3680 53564 3732
rect 53616 3720 53622 3732
rect 58250 3720 58256 3732
rect 53616 3692 58256 3720
rect 53616 3680 53622 3692
rect 58250 3680 58256 3692
rect 58308 3680 58314 3732
rect 47118 3612 47124 3664
rect 47176 3652 47182 3664
rect 50617 3655 50675 3661
rect 50617 3652 50629 3655
rect 47176 3624 50629 3652
rect 47176 3612 47182 3624
rect 50617 3621 50629 3624
rect 50663 3621 50675 3655
rect 50617 3615 50675 3621
rect 50890 3612 50896 3664
rect 50948 3652 50954 3664
rect 52089 3655 52147 3661
rect 52089 3652 52101 3655
rect 50948 3624 52101 3652
rect 50948 3612 50954 3624
rect 52089 3621 52101 3624
rect 52135 3621 52147 3655
rect 52089 3615 52147 3621
rect 53190 3612 53196 3664
rect 53248 3652 53254 3664
rect 54297 3655 54355 3661
rect 54297 3652 54309 3655
rect 53248 3624 54309 3652
rect 53248 3612 53254 3624
rect 54297 3621 54309 3624
rect 54343 3621 54355 3655
rect 54297 3615 54355 3621
rect 46934 3544 46940 3596
rect 46992 3584 46998 3596
rect 46992 3556 49004 3584
rect 46992 3544 46998 3556
rect 46615 3488 46704 3516
rect 46615 3485 46627 3488
rect 46569 3479 46627 3485
rect 46842 3476 46848 3528
rect 46900 3516 46906 3528
rect 48869 3519 48927 3525
rect 48869 3516 48881 3519
rect 46900 3488 48881 3516
rect 46900 3476 46906 3488
rect 48869 3485 48881 3488
rect 48915 3485 48927 3519
rect 48869 3479 48927 3485
rect 47118 3448 47124 3460
rect 46124 3420 47124 3448
rect 43956 3408 43962 3420
rect 47118 3408 47124 3420
rect 47176 3408 47182 3460
rect 47213 3451 47271 3457
rect 47213 3417 47225 3451
rect 47259 3417 47271 3451
rect 47213 3411 47271 3417
rect 39114 3380 39120 3392
rect 37240 3352 39120 3380
rect 37240 3340 37246 3352
rect 39114 3340 39120 3352
rect 39172 3340 39178 3392
rect 44542 3340 44548 3392
rect 44600 3380 44606 3392
rect 47228 3380 47256 3411
rect 47394 3408 47400 3460
rect 47452 3448 47458 3460
rect 47949 3451 48007 3457
rect 47949 3448 47961 3451
rect 47452 3420 47961 3448
rect 47452 3408 47458 3420
rect 47949 3417 47961 3420
rect 47995 3417 48007 3451
rect 47949 3411 48007 3417
rect 48685 3451 48743 3457
rect 48685 3417 48697 3451
rect 48731 3448 48743 3451
rect 48976 3448 49004 3556
rect 50798 3544 50804 3596
rect 50856 3584 50862 3596
rect 50856 3556 55214 3584
rect 50856 3544 50862 3556
rect 50614 3476 50620 3528
rect 50672 3516 50678 3528
rect 51077 3519 51135 3525
rect 51077 3516 51089 3519
rect 50672 3488 51089 3516
rect 50672 3476 50678 3488
rect 51077 3485 51089 3488
rect 51123 3485 51135 3519
rect 51077 3479 51135 3485
rect 51718 3476 51724 3528
rect 51776 3516 51782 3528
rect 52549 3519 52607 3525
rect 52549 3516 52561 3519
rect 51776 3488 52561 3516
rect 51776 3476 51782 3488
rect 52549 3485 52561 3488
rect 52595 3485 52607 3519
rect 53285 3519 53343 3525
rect 53285 3516 53297 3519
rect 52549 3479 52607 3485
rect 52656 3488 53297 3516
rect 48731 3420 49004 3448
rect 48731 3417 48743 3420
rect 48685 3411 48743 3417
rect 49234 3408 49240 3460
rect 49292 3448 49298 3460
rect 49421 3451 49479 3457
rect 49421 3448 49433 3451
rect 49292 3420 49433 3448
rect 49292 3408 49298 3420
rect 49421 3417 49433 3420
rect 49467 3417 49479 3451
rect 49421 3411 49479 3417
rect 49510 3408 49516 3460
rect 49568 3448 49574 3460
rect 50433 3451 50491 3457
rect 50433 3448 50445 3451
rect 49568 3420 50445 3448
rect 49568 3408 49574 3420
rect 50433 3417 50445 3420
rect 50479 3417 50491 3451
rect 50433 3411 50491 3417
rect 50890 3408 50896 3460
rect 50948 3448 50954 3460
rect 51905 3451 51963 3457
rect 51905 3448 51917 3451
rect 50948 3420 51917 3448
rect 50948 3408 50954 3420
rect 51905 3417 51917 3420
rect 51951 3417 51963 3451
rect 51905 3411 51963 3417
rect 52270 3408 52276 3460
rect 52328 3448 52334 3460
rect 52656 3448 52684 3488
rect 53285 3485 53297 3488
rect 53331 3485 53343 3519
rect 55186 3516 55214 3556
rect 56686 3544 56692 3596
rect 56744 3584 56750 3596
rect 56873 3587 56931 3593
rect 56873 3584 56885 3587
rect 56744 3556 56885 3584
rect 56744 3544 56750 3556
rect 56873 3553 56885 3556
rect 56919 3553 56931 3587
rect 56873 3547 56931 3553
rect 56045 3519 56103 3525
rect 56045 3516 56057 3519
rect 55186 3488 56057 3516
rect 53285 3479 53343 3485
rect 56045 3485 56057 3488
rect 56091 3485 56103 3519
rect 56045 3479 56103 3485
rect 56229 3519 56287 3525
rect 56229 3485 56241 3519
rect 56275 3516 56287 3519
rect 57422 3516 57428 3528
rect 56275 3488 57428 3516
rect 56275 3485 56287 3488
rect 56229 3479 56287 3485
rect 57422 3476 57428 3488
rect 57480 3476 57486 3528
rect 52328 3420 52684 3448
rect 52328 3408 52334 3420
rect 53190 3408 53196 3460
rect 53248 3448 53254 3460
rect 54113 3451 54171 3457
rect 54113 3448 54125 3451
rect 53248 3420 54125 3448
rect 53248 3408 53254 3420
rect 54113 3417 54125 3420
rect 54159 3417 54171 3451
rect 54113 3411 54171 3417
rect 56413 3451 56471 3457
rect 56413 3417 56425 3451
rect 56459 3448 56471 3451
rect 57118 3451 57176 3457
rect 57118 3448 57130 3451
rect 56459 3420 57130 3448
rect 56459 3417 56471 3420
rect 56413 3411 56471 3417
rect 57118 3417 57130 3420
rect 57164 3417 57176 3451
rect 57118 3411 57176 3417
rect 44600 3352 47256 3380
rect 44600 3340 44606 3352
rect 47302 3340 47308 3392
rect 47360 3380 47366 3392
rect 47360 3352 47405 3380
rect 47360 3340 47366 3352
rect 47578 3340 47584 3392
rect 47636 3380 47642 3392
rect 54662 3380 54668 3392
rect 47636 3352 54668 3380
rect 47636 3340 47642 3352
rect 54662 3340 54668 3352
rect 54720 3340 54726 3392
rect 57238 3340 57244 3392
rect 57296 3380 57302 3392
rect 58253 3383 58311 3389
rect 58253 3380 58265 3383
rect 57296 3352 58265 3380
rect 57296 3340 57302 3352
rect 58253 3349 58265 3352
rect 58299 3349 58311 3383
rect 58253 3343 58311 3349
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 5905 3179 5963 3185
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 5994 3176 6000 3188
rect 5951 3148 6000 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 5994 3136 6000 3148
rect 6052 3136 6058 3188
rect 6914 3176 6920 3188
rect 6875 3148 6920 3176
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 8386 3176 8392 3188
rect 8347 3148 8392 3176
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 9122 3176 9128 3188
rect 9083 3148 9128 3176
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9674 3176 9680 3188
rect 9646 3136 9680 3176
rect 9732 3136 9738 3188
rect 11149 3179 11207 3185
rect 11149 3145 11161 3179
rect 11195 3176 11207 3179
rect 11974 3176 11980 3188
rect 11195 3148 11980 3176
rect 11195 3145 11207 3148
rect 11149 3139 11207 3145
rect 11974 3136 11980 3148
rect 12032 3136 12038 3188
rect 12713 3179 12771 3185
rect 12713 3145 12725 3179
rect 12759 3176 12771 3179
rect 15010 3176 15016 3188
rect 12759 3148 15016 3176
rect 12759 3145 12771 3148
rect 12713 3139 12771 3145
rect 15010 3136 15016 3148
rect 15068 3136 15074 3188
rect 18432 3148 22094 3176
rect 5813 3111 5871 3117
rect 5813 3077 5825 3111
rect 5859 3108 5871 3111
rect 8110 3108 8116 3120
rect 5859 3080 8116 3108
rect 5859 3077 5871 3080
rect 5813 3071 5871 3077
rect 8110 3068 8116 3080
rect 8168 3068 8174 3120
rect 9646 3108 9674 3136
rect 10686 3108 10692 3120
rect 8220 3080 9674 3108
rect 10060 3080 10692 3108
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 8220 3040 8248 3080
rect 7607 3012 8248 3040
rect 8297 3043 8355 3049
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 8846 3040 8852 3052
rect 8343 3012 8852 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 6840 2972 6868 3003
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 9030 3040 9036 3052
rect 8991 3012 9036 3040
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 9674 3040 9680 3052
rect 9324 3012 9680 3040
rect 9214 2972 9220 2984
rect 6840 2944 9220 2972
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 7745 2907 7803 2913
rect 7745 2873 7757 2907
rect 7791 2904 7803 2907
rect 9324 2904 9352 3012
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 10060 3049 10088 3080
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 11882 3108 11888 3120
rect 11843 3080 11888 3108
rect 11882 3068 11888 3080
rect 11940 3068 11946 3120
rect 12069 3111 12127 3117
rect 12069 3077 12081 3111
rect 12115 3108 12127 3111
rect 13357 3111 13415 3117
rect 12115 3080 13308 3108
rect 12115 3077 12127 3080
rect 12069 3071 12127 3077
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 12621 3043 12679 3049
rect 10192 3012 10237 3040
rect 10192 3000 10198 3012
rect 12621 3009 12633 3043
rect 12667 3009 12679 3043
rect 13280 3040 13308 3080
rect 13357 3077 13369 3111
rect 13403 3108 13415 3111
rect 15197 3111 15255 3117
rect 13403 3080 15148 3108
rect 13403 3077 13415 3080
rect 13357 3071 13415 3077
rect 13814 3040 13820 3052
rect 13280 3012 13820 3040
rect 12621 3003 12679 3009
rect 9398 2932 9404 2984
rect 9456 2972 9462 2984
rect 9858 2972 9864 2984
rect 9456 2944 9720 2972
rect 9771 2944 9864 2972
rect 9456 2932 9462 2944
rect 9692 2913 9720 2944
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 9953 2975 10011 2981
rect 9953 2941 9965 2975
rect 9999 2972 10011 2975
rect 12250 2972 12256 2984
rect 9999 2944 12256 2972
rect 9999 2941 10011 2944
rect 9953 2935 10011 2941
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 12636 2972 12664 3003
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 14001 3043 14059 3049
rect 14001 3009 14013 3043
rect 14047 3040 14059 3043
rect 14274 3040 14280 3052
rect 14047 3012 14280 3040
rect 14047 3009 14059 3012
rect 14001 3003 14059 3009
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 14826 3000 14832 3052
rect 14884 3040 14890 3052
rect 14921 3043 14979 3049
rect 14921 3040 14933 3043
rect 14884 3012 14933 3040
rect 14884 3000 14890 3012
rect 14921 3009 14933 3012
rect 14967 3009 14979 3043
rect 15120 3040 15148 3080
rect 15197 3077 15209 3111
rect 15243 3108 15255 3111
rect 17494 3108 17500 3120
rect 15243 3080 17500 3108
rect 15243 3077 15255 3080
rect 15197 3071 15255 3077
rect 17494 3068 17500 3080
rect 17552 3068 17558 3120
rect 18432 3117 18460 3148
rect 19334 3117 19340 3120
rect 18417 3111 18475 3117
rect 18417 3077 18429 3111
rect 18463 3077 18475 3111
rect 18417 3071 18475 3077
rect 19328 3071 19340 3117
rect 19392 3108 19398 3120
rect 19392 3080 19428 3108
rect 19334 3068 19340 3071
rect 19392 3068 19398 3080
rect 15562 3040 15568 3052
rect 15120 3012 15568 3040
rect 14921 3003 14979 3009
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3040 15899 3043
rect 16482 3040 16488 3052
rect 15887 3012 16488 3040
rect 15887 3009 15899 3012
rect 15841 3003 15899 3009
rect 16482 3000 16488 3012
rect 16540 3000 16546 3052
rect 17218 3040 17224 3052
rect 17179 3012 17224 3040
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 17420 3012 18092 3040
rect 14185 2975 14243 2981
rect 12636 2944 14136 2972
rect 7791 2876 9352 2904
rect 9677 2907 9735 2913
rect 7791 2873 7803 2876
rect 7745 2867 7803 2873
rect 9677 2873 9689 2907
rect 9723 2873 9735 2907
rect 9872 2904 9900 2932
rect 9872 2876 9996 2904
rect 9677 2867 9735 2873
rect 8846 2796 8852 2848
rect 8904 2836 8910 2848
rect 9858 2836 9864 2848
rect 8904 2808 9864 2836
rect 8904 2796 8910 2808
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 9968 2836 9996 2876
rect 10870 2864 10876 2916
rect 10928 2904 10934 2916
rect 10965 2907 11023 2913
rect 10965 2904 10977 2907
rect 10928 2876 10977 2904
rect 10928 2864 10934 2876
rect 10965 2873 10977 2876
rect 11011 2873 11023 2907
rect 13538 2904 13544 2916
rect 13499 2876 13544 2904
rect 10965 2867 11023 2873
rect 13538 2864 13544 2876
rect 13596 2864 13602 2916
rect 12618 2836 12624 2848
rect 9968 2808 12624 2836
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 14108 2836 14136 2944
rect 14185 2941 14197 2975
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 16117 2975 16175 2981
rect 16117 2941 16129 2975
rect 16163 2972 16175 2975
rect 17420 2972 17448 3012
rect 16163 2944 17448 2972
rect 17497 2975 17555 2981
rect 16163 2941 16175 2944
rect 16117 2935 16175 2941
rect 17497 2941 17509 2975
rect 17543 2941 17555 2975
rect 18064 2972 18092 3012
rect 18138 3000 18144 3052
rect 18196 3040 18202 3052
rect 19058 3040 19064 3052
rect 18196 3012 18241 3040
rect 19019 3012 19064 3040
rect 18196 3000 18202 3012
rect 19058 3000 19064 3012
rect 19116 3000 19122 3052
rect 20162 3040 20168 3052
rect 19168 3012 20168 3040
rect 19168 2972 19196 3012
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 20993 3043 21051 3049
rect 20993 3009 21005 3043
rect 21039 3040 21051 3043
rect 21174 3040 21180 3052
rect 21039 3012 21180 3040
rect 21039 3009 21051 3012
rect 20993 3003 21051 3009
rect 21174 3000 21180 3012
rect 21232 3000 21238 3052
rect 22066 3040 22094 3148
rect 22278 3136 22284 3188
rect 22336 3176 22342 3188
rect 33410 3176 33416 3188
rect 22336 3148 33416 3176
rect 22336 3136 22342 3148
rect 33410 3136 33416 3148
rect 33468 3136 33474 3188
rect 33778 3136 33784 3188
rect 33836 3176 33842 3188
rect 33836 3148 36308 3176
rect 33836 3136 33842 3148
rect 23198 3108 23204 3120
rect 22572 3080 23204 3108
rect 22186 3040 22192 3052
rect 22066 3012 22192 3040
rect 22186 3000 22192 3012
rect 22244 3000 22250 3052
rect 22572 3049 22600 3080
rect 23198 3068 23204 3080
rect 23256 3068 23262 3120
rect 23934 3108 23940 3120
rect 23492 3080 23940 3108
rect 23492 3049 23520 3080
rect 23934 3068 23940 3080
rect 23992 3068 23998 3120
rect 28804 3111 28862 3117
rect 26160 3080 28764 3108
rect 22557 3043 22615 3049
rect 22557 3009 22569 3043
rect 22603 3009 22615 3043
rect 23477 3043 23535 3049
rect 22557 3003 22615 3009
rect 22756 3012 22968 3040
rect 21082 2972 21088 2984
rect 18064 2944 19196 2972
rect 20180 2944 21088 2972
rect 17497 2935 17555 2941
rect 14200 2904 14228 2935
rect 16390 2904 16396 2916
rect 14200 2876 16396 2904
rect 16390 2864 16396 2876
rect 16448 2864 16454 2916
rect 15010 2836 15016 2848
rect 14108 2808 15016 2836
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 17512 2836 17540 2935
rect 20180 2836 20208 2944
rect 21082 2932 21088 2944
rect 21140 2932 21146 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 22756 2972 22784 3012
rect 21315 2944 22784 2972
rect 22833 2975 22891 2981
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 22833 2941 22845 2975
rect 22879 2941 22891 2975
rect 22940 2972 22968 3012
rect 23477 3009 23489 3043
rect 23523 3009 23535 3043
rect 23477 3003 23535 3009
rect 23566 3000 23572 3052
rect 23624 3000 23630 3052
rect 23744 3043 23802 3049
rect 23744 3009 23756 3043
rect 23790 3040 23802 3043
rect 24578 3040 24584 3052
rect 23790 3012 24584 3040
rect 23790 3009 23802 3012
rect 23744 3003 23802 3009
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 26160 3049 26188 3080
rect 26145 3043 26203 3049
rect 26145 3009 26157 3043
rect 26191 3009 26203 3043
rect 26145 3003 26203 3009
rect 27157 3043 27215 3049
rect 27157 3009 27169 3043
rect 27203 3040 27215 3043
rect 27203 3012 28028 3040
rect 27203 3009 27215 3012
rect 27157 3003 27215 3009
rect 23584 2972 23612 3000
rect 22940 2944 23612 2972
rect 22833 2935 22891 2941
rect 20254 2864 20260 2916
rect 20312 2904 20318 2916
rect 20312 2876 22094 2904
rect 20312 2864 20318 2876
rect 17512 2808 20208 2836
rect 20441 2839 20499 2845
rect 20441 2805 20453 2839
rect 20487 2836 20499 2839
rect 20714 2836 20720 2848
rect 20487 2808 20720 2836
rect 20487 2805 20499 2808
rect 20441 2799 20499 2805
rect 20714 2796 20720 2808
rect 20772 2796 20778 2848
rect 22066 2836 22094 2876
rect 22738 2836 22744 2848
rect 22066 2808 22744 2836
rect 22738 2796 22744 2808
rect 22796 2796 22802 2848
rect 22848 2836 22876 2935
rect 26050 2932 26056 2984
rect 26108 2972 26114 2984
rect 26329 2975 26387 2981
rect 26329 2972 26341 2975
rect 26108 2944 26341 2972
rect 26108 2932 26114 2944
rect 26329 2941 26341 2944
rect 26375 2941 26387 2975
rect 26329 2935 26387 2941
rect 26418 2932 26424 2984
rect 26476 2972 26482 2984
rect 27341 2975 27399 2981
rect 27341 2972 27353 2975
rect 26476 2944 27353 2972
rect 26476 2932 26482 2944
rect 27341 2941 27353 2944
rect 27387 2941 27399 2975
rect 27341 2935 27399 2941
rect 24854 2904 24860 2916
rect 24815 2876 24860 2904
rect 24854 2864 24860 2876
rect 24912 2864 24918 2916
rect 24946 2864 24952 2916
rect 25004 2904 25010 2916
rect 27706 2904 27712 2916
rect 25004 2876 27712 2904
rect 25004 2864 25010 2876
rect 27706 2864 27712 2876
rect 27764 2864 27770 2916
rect 28000 2904 28028 3012
rect 28074 3000 28080 3052
rect 28132 3040 28138 3052
rect 28537 3043 28595 3049
rect 28537 3040 28549 3043
rect 28132 3012 28549 3040
rect 28132 3000 28138 3012
rect 28537 3009 28549 3012
rect 28583 3009 28595 3043
rect 28736 3040 28764 3080
rect 28804 3077 28816 3111
rect 28850 3108 28862 3111
rect 29270 3108 29276 3120
rect 28850 3080 29276 3108
rect 28850 3077 28862 3080
rect 28804 3071 28862 3077
rect 29270 3068 29276 3080
rect 29328 3068 29334 3120
rect 30742 3068 30748 3120
rect 30800 3068 30806 3120
rect 32398 3068 32404 3120
rect 32456 3108 32462 3120
rect 36280 3117 36308 3148
rect 37918 3136 37924 3188
rect 37976 3176 37982 3188
rect 39942 3176 39948 3188
rect 37976 3148 39948 3176
rect 37976 3136 37982 3148
rect 39942 3136 39948 3148
rect 40000 3136 40006 3188
rect 42794 3176 42800 3188
rect 42755 3148 42800 3176
rect 42794 3136 42800 3148
rect 42852 3136 42858 3188
rect 43898 3136 43904 3188
rect 43956 3176 43962 3188
rect 46937 3179 46995 3185
rect 46937 3176 46949 3179
rect 43956 3148 46949 3176
rect 43956 3136 43962 3148
rect 46937 3145 46949 3148
rect 46983 3145 46995 3179
rect 47946 3176 47952 3188
rect 47907 3148 47952 3176
rect 46937 3139 46995 3145
rect 47946 3136 47952 3148
rect 48004 3136 48010 3188
rect 48682 3176 48688 3188
rect 48643 3148 48688 3176
rect 48682 3136 48688 3148
rect 48740 3136 48746 3188
rect 49786 3176 49792 3188
rect 49747 3148 49792 3176
rect 49786 3136 49792 3148
rect 49844 3136 49850 3188
rect 50525 3179 50583 3185
rect 50525 3145 50537 3179
rect 50571 3176 50583 3179
rect 50982 3176 50988 3188
rect 50571 3148 50988 3176
rect 50571 3145 50583 3148
rect 50525 3139 50583 3145
rect 50982 3136 50988 3148
rect 51040 3136 51046 3188
rect 51997 3179 52055 3185
rect 51997 3145 52009 3179
rect 52043 3176 52055 3179
rect 52178 3176 52184 3188
rect 52043 3148 52184 3176
rect 52043 3145 52055 3148
rect 51997 3139 52055 3145
rect 52178 3136 52184 3148
rect 52236 3136 52242 3188
rect 52454 3136 52460 3188
rect 52512 3176 52518 3188
rect 53837 3179 53895 3185
rect 53837 3176 53849 3179
rect 52512 3148 53849 3176
rect 52512 3136 52518 3148
rect 53837 3145 53849 3148
rect 53883 3145 53895 3179
rect 53837 3139 53895 3145
rect 53926 3136 53932 3188
rect 53984 3176 53990 3188
rect 55309 3179 55367 3185
rect 55309 3176 55321 3179
rect 53984 3148 55321 3176
rect 53984 3136 53990 3148
rect 55309 3145 55321 3148
rect 55355 3145 55367 3179
rect 58250 3176 58256 3188
rect 55309 3139 55367 3145
rect 57164 3148 58256 3176
rect 34425 3111 34483 3117
rect 34425 3108 34437 3111
rect 32456 3080 34437 3108
rect 32456 3068 32462 3080
rect 34425 3077 34437 3080
rect 34471 3077 34483 3111
rect 34425 3071 34483 3077
rect 36265 3111 36323 3117
rect 36265 3077 36277 3111
rect 36311 3077 36323 3111
rect 36265 3071 36323 3077
rect 39390 3068 39396 3120
rect 39448 3108 39454 3120
rect 39666 3108 39672 3120
rect 39448 3080 39672 3108
rect 39448 3068 39454 3080
rect 39666 3068 39672 3080
rect 39724 3068 39730 3120
rect 40681 3111 40739 3117
rect 40681 3077 40693 3111
rect 40727 3108 40739 3111
rect 40862 3108 40868 3120
rect 40727 3080 40868 3108
rect 40727 3077 40739 3080
rect 40681 3071 40739 3077
rect 40862 3068 40868 3080
rect 40920 3068 40926 3120
rect 41598 3108 41604 3120
rect 41559 3080 41604 3108
rect 41598 3068 41604 3080
rect 41656 3068 41662 3120
rect 45002 3068 45008 3120
rect 45060 3108 45066 3120
rect 45060 3080 47808 3108
rect 45060 3068 45066 3080
rect 30760 3040 30788 3068
rect 28736 3012 30788 3040
rect 30837 3043 30895 3049
rect 28537 3003 28595 3009
rect 30837 3009 30849 3043
rect 30883 3040 30895 3043
rect 31202 3040 31208 3052
rect 30883 3012 31208 3040
rect 30883 3009 30895 3012
rect 30837 3003 30895 3009
rect 31202 3000 31208 3012
rect 31260 3000 31266 3052
rect 31478 3000 31484 3052
rect 31536 3040 31542 3052
rect 32309 3043 32367 3049
rect 32309 3040 32321 3043
rect 31536 3012 32321 3040
rect 31536 3000 31542 3012
rect 32309 3009 32321 3012
rect 32355 3009 32367 3043
rect 33226 3040 33232 3052
rect 33187 3012 33232 3040
rect 32309 3003 32367 3009
rect 33226 3000 33232 3012
rect 33284 3000 33290 3052
rect 33336 3012 33548 3040
rect 30742 2932 30748 2984
rect 30800 2972 30806 2984
rect 31021 2975 31079 2981
rect 31021 2972 31033 2975
rect 30800 2944 31033 2972
rect 30800 2932 30806 2944
rect 31021 2941 31033 2944
rect 31067 2941 31079 2975
rect 31021 2935 31079 2941
rect 31570 2932 31576 2984
rect 31628 2972 31634 2984
rect 32493 2975 32551 2981
rect 32493 2972 32505 2975
rect 31628 2944 32505 2972
rect 31628 2932 31634 2944
rect 32493 2941 32505 2944
rect 32539 2941 32551 2975
rect 32493 2935 32551 2941
rect 32950 2932 32956 2984
rect 33008 2972 33014 2984
rect 33336 2972 33364 3012
rect 33008 2944 33364 2972
rect 33413 2975 33471 2981
rect 33008 2932 33014 2944
rect 33413 2941 33425 2975
rect 33459 2941 33471 2975
rect 33520 2972 33548 3012
rect 33962 3000 33968 3052
rect 34020 3040 34026 3052
rect 34149 3043 34207 3049
rect 34149 3040 34161 3043
rect 34020 3012 34161 3040
rect 34020 3000 34026 3012
rect 34149 3009 34161 3012
rect 34195 3009 34207 3043
rect 34149 3003 34207 3009
rect 34514 3000 34520 3052
rect 34572 3040 34578 3052
rect 35069 3043 35127 3049
rect 35069 3040 35081 3043
rect 34572 3012 35081 3040
rect 34572 3000 34578 3012
rect 35069 3009 35081 3012
rect 35115 3009 35127 3043
rect 35069 3003 35127 3009
rect 35802 3000 35808 3052
rect 35860 3040 35866 3052
rect 35989 3043 36047 3049
rect 35989 3040 36001 3043
rect 35860 3012 36001 3040
rect 35860 3000 35866 3012
rect 35989 3009 36001 3012
rect 36035 3009 36047 3043
rect 37458 3040 37464 3052
rect 37419 3012 37464 3040
rect 35989 3003 36047 3009
rect 37458 3000 37464 3012
rect 37516 3000 37522 3052
rect 38381 3043 38439 3049
rect 37568 3012 37780 3040
rect 35253 2975 35311 2981
rect 35253 2972 35265 2975
rect 33520 2944 35265 2972
rect 33413 2935 33471 2941
rect 35253 2941 35265 2944
rect 35299 2941 35311 2975
rect 35253 2935 35311 2941
rect 28000 2876 28580 2904
rect 24394 2836 24400 2848
rect 22848 2808 24400 2836
rect 24394 2796 24400 2808
rect 24452 2796 24458 2848
rect 25685 2839 25743 2845
rect 25685 2805 25697 2839
rect 25731 2836 25743 2839
rect 27982 2836 27988 2848
rect 25731 2808 27988 2836
rect 25731 2805 25743 2808
rect 25685 2799 25743 2805
rect 27982 2796 27988 2808
rect 28040 2796 28046 2848
rect 28552 2836 28580 2876
rect 29730 2864 29736 2916
rect 29788 2904 29794 2916
rect 29917 2907 29975 2913
rect 29917 2904 29929 2907
rect 29788 2876 29929 2904
rect 29788 2864 29794 2876
rect 29917 2873 29929 2876
rect 29963 2873 29975 2907
rect 29917 2867 29975 2873
rect 32122 2864 32128 2916
rect 32180 2904 32186 2916
rect 33428 2904 33456 2935
rect 35618 2932 35624 2984
rect 35676 2972 35682 2984
rect 37568 2972 37596 3012
rect 35676 2944 37596 2972
rect 37645 2975 37703 2981
rect 35676 2932 35682 2944
rect 37645 2941 37657 2975
rect 37691 2941 37703 2975
rect 37752 2972 37780 3012
rect 38381 3009 38393 3043
rect 38427 3040 38439 3043
rect 38654 3040 38660 3052
rect 38427 3012 38660 3040
rect 38427 3009 38439 3012
rect 38381 3003 38439 3009
rect 38654 3000 38660 3012
rect 38712 3000 38718 3052
rect 39298 3040 39304 3052
rect 39259 3012 39304 3040
rect 39298 3000 39304 3012
rect 39356 3000 39362 3052
rect 39574 3000 39580 3052
rect 39632 3040 39638 3052
rect 40313 3043 40371 3049
rect 40313 3040 40325 3043
rect 39632 3012 40325 3040
rect 39632 3000 39638 3012
rect 40313 3009 40325 3012
rect 40359 3009 40371 3043
rect 40313 3003 40371 3009
rect 40402 3000 40408 3052
rect 40460 3040 40466 3052
rect 41233 3043 41291 3049
rect 41233 3040 41245 3043
rect 40460 3012 41245 3040
rect 40460 3000 40466 3012
rect 41233 3009 41245 3012
rect 41279 3009 41291 3043
rect 41233 3003 41291 3009
rect 41322 3000 41328 3052
rect 41380 3040 41386 3052
rect 42705 3043 42763 3049
rect 42705 3040 42717 3043
rect 41380 3012 42717 3040
rect 41380 3000 41386 3012
rect 42705 3009 42717 3012
rect 42751 3009 42763 3043
rect 42705 3003 42763 3009
rect 44266 3000 44272 3052
rect 44324 3040 44330 3052
rect 44545 3043 44603 3049
rect 44545 3040 44557 3043
rect 44324 3012 44557 3040
rect 44324 3000 44330 3012
rect 44545 3009 44557 3012
rect 44591 3009 44603 3043
rect 44545 3003 44603 3009
rect 44637 3043 44695 3049
rect 44637 3009 44649 3043
rect 44683 3009 44695 3043
rect 44910 3040 44916 3052
rect 44871 3012 44916 3040
rect 44637 3003 44695 3009
rect 38565 2975 38623 2981
rect 38565 2972 38577 2975
rect 37752 2944 38577 2972
rect 37645 2935 37703 2941
rect 38565 2941 38577 2944
rect 38611 2941 38623 2975
rect 38565 2935 38623 2941
rect 39485 2975 39543 2981
rect 39485 2941 39497 2975
rect 39531 2941 39543 2975
rect 39485 2935 39543 2941
rect 32180 2876 33456 2904
rect 32180 2864 32186 2876
rect 35342 2864 35348 2916
rect 35400 2904 35406 2916
rect 37660 2904 37688 2935
rect 35400 2876 37688 2904
rect 35400 2864 35406 2876
rect 31754 2836 31760 2848
rect 28552 2808 31760 2836
rect 31754 2796 31760 2808
rect 31812 2796 31818 2848
rect 31846 2796 31852 2848
rect 31904 2836 31910 2848
rect 33410 2836 33416 2848
rect 31904 2808 33416 2836
rect 31904 2796 31910 2808
rect 33410 2796 33416 2808
rect 33468 2796 33474 2848
rect 33594 2796 33600 2848
rect 33652 2836 33658 2848
rect 35986 2836 35992 2848
rect 33652 2808 35992 2836
rect 33652 2796 33658 2808
rect 35986 2796 35992 2808
rect 36044 2796 36050 2848
rect 36538 2796 36544 2848
rect 36596 2836 36602 2848
rect 39500 2836 39528 2935
rect 42334 2932 42340 2984
rect 42392 2972 42398 2984
rect 44450 2972 44456 2984
rect 42392 2944 44456 2972
rect 42392 2932 42398 2944
rect 44450 2932 44456 2944
rect 44508 2932 44514 2984
rect 44652 2972 44680 3003
rect 44910 3000 44916 3012
rect 44968 3000 44974 3052
rect 45094 3000 45100 3052
rect 45152 3040 45158 3052
rect 45189 3043 45247 3049
rect 45189 3040 45201 3043
rect 45152 3012 45201 3040
rect 45152 3000 45158 3012
rect 45189 3009 45201 3012
rect 45235 3009 45247 3043
rect 45189 3003 45247 3009
rect 45465 3043 45523 3049
rect 45465 3009 45477 3043
rect 45511 3040 45523 3043
rect 45738 3040 45744 3052
rect 45511 3012 45744 3040
rect 45511 3009 45523 3012
rect 45465 3003 45523 3009
rect 45738 3000 45744 3012
rect 45796 3000 45802 3052
rect 46106 3040 46112 3052
rect 46067 3012 46112 3040
rect 46106 3000 46112 3012
rect 46164 3000 46170 3052
rect 47780 3049 47808 3080
rect 51534 3068 51540 3120
rect 51592 3108 51598 3120
rect 53009 3111 53067 3117
rect 53009 3108 53021 3111
rect 51592 3080 53021 3108
rect 51592 3068 51598 3080
rect 53009 3077 53021 3080
rect 53055 3077 53067 3111
rect 53009 3071 53067 3077
rect 53374 3068 53380 3120
rect 53432 3108 53438 3120
rect 55217 3111 55275 3117
rect 55217 3108 55229 3111
rect 53432 3080 55229 3108
rect 53432 3068 53438 3080
rect 55217 3077 55229 3080
rect 55263 3077 55275 3111
rect 56594 3108 56600 3120
rect 56555 3080 56600 3108
rect 55217 3071 55275 3077
rect 56594 3068 56600 3080
rect 56652 3068 56658 3120
rect 46845 3043 46903 3049
rect 46845 3009 46857 3043
rect 46891 3009 46903 3043
rect 46845 3003 46903 3009
rect 47765 3043 47823 3049
rect 47765 3009 47777 3043
rect 47811 3009 47823 3043
rect 47765 3003 47823 3009
rect 44652 2944 45554 2972
rect 44177 2907 44235 2913
rect 44177 2873 44189 2907
rect 44223 2904 44235 2907
rect 44818 2904 44824 2916
rect 44223 2876 44824 2904
rect 44223 2873 44235 2876
rect 44177 2867 44235 2873
rect 44818 2864 44824 2876
rect 44876 2864 44882 2916
rect 45526 2904 45554 2944
rect 45646 2932 45652 2984
rect 45704 2972 45710 2984
rect 46860 2972 46888 3003
rect 48406 3000 48412 3052
rect 48464 3040 48470 3052
rect 48593 3043 48651 3049
rect 48593 3040 48605 3043
rect 48464 3012 48605 3040
rect 48464 3000 48470 3012
rect 48593 3009 48605 3012
rect 48639 3009 48651 3043
rect 48593 3003 48651 3009
rect 48682 3000 48688 3052
rect 48740 3040 48746 3052
rect 49513 3043 49571 3049
rect 49513 3040 49525 3043
rect 48740 3012 49525 3040
rect 48740 3000 48746 3012
rect 49513 3009 49525 3012
rect 49559 3009 49571 3043
rect 50341 3043 50399 3049
rect 50341 3040 50353 3043
rect 49513 3003 49571 3009
rect 49620 3012 50353 3040
rect 45704 2944 46888 2972
rect 45704 2932 45710 2944
rect 48130 2932 48136 2984
rect 48188 2972 48194 2984
rect 49620 2972 49648 3012
rect 50341 3009 50353 3012
rect 50387 3009 50399 3043
rect 50341 3003 50399 3009
rect 51169 3043 51227 3049
rect 51169 3009 51181 3043
rect 51215 3009 51227 3043
rect 51169 3003 51227 3009
rect 51813 3043 51871 3049
rect 51813 3009 51825 3043
rect 51859 3009 51871 3043
rect 51813 3003 51871 3009
rect 48188 2944 49648 2972
rect 48188 2932 48194 2944
rect 49786 2932 49792 2984
rect 49844 2972 49850 2984
rect 51184 2972 51212 3003
rect 49844 2944 51212 2972
rect 49844 2932 49850 2944
rect 47302 2904 47308 2916
rect 45526 2876 47308 2904
rect 47302 2864 47308 2876
rect 47360 2864 47366 2916
rect 50062 2864 50068 2916
rect 50120 2904 50126 2916
rect 51828 2904 51856 3003
rect 51994 3000 52000 3052
rect 52052 3040 52058 3052
rect 53745 3043 53803 3049
rect 53745 3040 53757 3043
rect 52052 3012 53757 3040
rect 52052 3000 52058 3012
rect 53745 3009 53757 3012
rect 53791 3009 53803 3043
rect 53745 3003 53803 3009
rect 54481 3043 54539 3049
rect 54481 3009 54493 3043
rect 54527 3009 54539 3043
rect 54662 3040 54668 3052
rect 54623 3012 54668 3040
rect 54481 3003 54539 3009
rect 52546 2932 52552 2984
rect 52604 2972 52610 2984
rect 54496 2972 54524 3003
rect 54662 3000 54668 3012
rect 54720 3000 54726 3052
rect 56413 3043 56471 3049
rect 56413 3009 56425 3043
rect 56459 3040 56471 3043
rect 56502 3040 56508 3052
rect 56459 3012 56508 3040
rect 56459 3009 56471 3012
rect 56413 3003 56471 3009
rect 56502 3000 56508 3012
rect 56560 3000 56566 3052
rect 57164 3049 57192 3148
rect 58250 3136 58256 3148
rect 58308 3136 58314 3188
rect 58158 3108 58164 3120
rect 58119 3080 58164 3108
rect 58158 3068 58164 3080
rect 58216 3068 58222 3120
rect 57149 3043 57207 3049
rect 57149 3009 57161 3043
rect 57195 3009 57207 3043
rect 57149 3003 57207 3009
rect 57241 3043 57299 3049
rect 57241 3009 57253 3043
rect 57287 3040 57299 3043
rect 57974 3040 57980 3052
rect 57287 3012 57980 3040
rect 57287 3009 57299 3012
rect 57241 3003 57299 3009
rect 57974 3000 57980 3012
rect 58032 3000 58038 3052
rect 52604 2944 54524 2972
rect 52604 2932 52610 2944
rect 55306 2932 55312 2984
rect 55364 2972 55370 2984
rect 57425 2975 57483 2981
rect 57425 2972 57437 2975
rect 55364 2944 57437 2972
rect 55364 2932 55370 2944
rect 57425 2941 57437 2944
rect 57471 2941 57483 2975
rect 57425 2935 57483 2941
rect 50120 2876 51856 2904
rect 50120 2864 50126 2876
rect 36596 2808 39528 2836
rect 36596 2796 36602 2808
rect 40678 2796 40684 2848
rect 40736 2836 40742 2848
rect 41414 2836 41420 2848
rect 40736 2808 41420 2836
rect 40736 2796 40742 2808
rect 41414 2796 41420 2808
rect 41472 2796 41478 2848
rect 43438 2796 43444 2848
rect 43496 2836 43502 2848
rect 44910 2836 44916 2848
rect 43496 2808 44916 2836
rect 43496 2796 43502 2808
rect 44910 2796 44916 2808
rect 44968 2796 44974 2848
rect 45278 2796 45284 2848
rect 45336 2836 45342 2848
rect 46201 2839 46259 2845
rect 46201 2836 46213 2839
rect 45336 2808 46213 2836
rect 45336 2796 45342 2808
rect 46201 2805 46213 2808
rect 46247 2805 46259 2839
rect 46201 2799 46259 2805
rect 46382 2796 46388 2848
rect 46440 2836 46446 2848
rect 51261 2839 51319 2845
rect 51261 2836 51273 2839
rect 46440 2808 51273 2836
rect 46440 2796 46446 2808
rect 51261 2805 51273 2808
rect 51307 2805 51319 2839
rect 51261 2799 51319 2805
rect 51350 2796 51356 2848
rect 51408 2836 51414 2848
rect 53101 2839 53159 2845
rect 53101 2836 53113 2839
rect 51408 2808 53113 2836
rect 51408 2796 51414 2808
rect 53101 2805 53113 2808
rect 53147 2805 53159 2839
rect 53101 2799 53159 2805
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 10597 2635 10655 2641
rect 5951 2604 10548 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 10520 2576 10548 2604
rect 10597 2601 10609 2635
rect 10643 2632 10655 2635
rect 10778 2632 10784 2644
rect 10643 2604 10784 2632
rect 10643 2601 10655 2604
rect 10597 2595 10655 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 14734 2632 14740 2644
rect 12084 2604 14740 2632
rect 8478 2564 8484 2576
rect 6932 2536 8484 2564
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 1854 2428 1860 2440
rect 1815 2400 1860 2428
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 6822 2428 6828 2440
rect 5123 2400 6828 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 6932 2437 6960 2536
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 8573 2567 8631 2573
rect 8573 2533 8585 2567
rect 8619 2564 8631 2567
rect 8662 2564 8668 2576
rect 8619 2536 8668 2564
rect 8619 2533 8631 2536
rect 8573 2527 8631 2533
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 10410 2564 10416 2576
rect 10371 2536 10416 2564
rect 10410 2524 10416 2536
rect 10468 2524 10474 2576
rect 10502 2524 10508 2576
rect 10560 2524 10566 2576
rect 9582 2496 9588 2508
rect 7668 2468 9588 2496
rect 7668 2437 7696 2468
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 10137 2499 10195 2505
rect 10137 2465 10149 2499
rect 10183 2496 10195 2499
rect 10686 2496 10692 2508
rect 10183 2468 10692 2496
rect 10183 2465 10195 2468
rect 10137 2459 10195 2465
rect 10686 2456 10692 2468
rect 10744 2456 10750 2508
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 5813 2363 5871 2369
rect 5813 2329 5825 2363
rect 5859 2360 5871 2363
rect 8389 2363 8447 2369
rect 5859 2332 8156 2360
rect 5859 2329 5871 2332
rect 5813 2323 5871 2329
rect 5166 2292 5172 2304
rect 5127 2264 5172 2292
rect 5166 2252 5172 2264
rect 5224 2252 5230 2304
rect 7006 2292 7012 2304
rect 6967 2264 7012 2292
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 7742 2292 7748 2304
rect 7703 2264 7748 2292
rect 7742 2252 7748 2264
rect 7800 2252 7806 2304
rect 8128 2292 8156 2332
rect 8389 2329 8401 2363
rect 8435 2360 8447 2363
rect 9398 2360 9404 2372
rect 8435 2332 9404 2360
rect 8435 2329 8447 2332
rect 8389 2323 8447 2329
rect 9398 2320 9404 2332
rect 9456 2320 9462 2372
rect 8938 2292 8944 2304
rect 8128 2264 8944 2292
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 9508 2292 9536 2391
rect 9674 2360 9680 2372
rect 9635 2332 9680 2360
rect 9674 2320 9680 2332
rect 9732 2320 9738 2372
rect 12084 2369 12112 2604
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 17037 2635 17095 2641
rect 17037 2601 17049 2635
rect 17083 2632 17095 2635
rect 18874 2632 18880 2644
rect 17083 2604 18880 2632
rect 17083 2601 17095 2604
rect 17037 2595 17095 2601
rect 18874 2592 18880 2604
rect 18932 2592 18938 2644
rect 22097 2635 22155 2641
rect 22097 2632 22109 2635
rect 18984 2604 22109 2632
rect 12253 2567 12311 2573
rect 12253 2533 12265 2567
rect 12299 2564 12311 2567
rect 13170 2564 13176 2576
rect 12299 2536 13176 2564
rect 12299 2533 12311 2536
rect 12253 2527 12311 2533
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 13725 2567 13783 2573
rect 13725 2533 13737 2567
rect 13771 2564 13783 2567
rect 14366 2564 14372 2576
rect 13771 2536 14372 2564
rect 13771 2533 13783 2536
rect 13725 2527 13783 2533
rect 14366 2524 14372 2536
rect 14424 2524 14430 2576
rect 18984 2564 19012 2604
rect 22097 2601 22109 2604
rect 22143 2601 22155 2635
rect 22097 2595 22155 2601
rect 24765 2635 24823 2641
rect 24765 2601 24777 2635
rect 24811 2632 24823 2635
rect 24946 2632 24952 2644
rect 24811 2604 24952 2632
rect 24811 2601 24823 2604
rect 24765 2595 24823 2601
rect 24946 2592 24952 2604
rect 25004 2592 25010 2644
rect 27062 2632 27068 2644
rect 25148 2604 27068 2632
rect 24210 2564 24216 2576
rect 17512 2536 19012 2564
rect 22572 2536 24216 2564
rect 16022 2496 16028 2508
rect 13556 2468 16028 2496
rect 13556 2437 13584 2468
rect 16022 2456 16028 2468
rect 16080 2456 16086 2508
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2397 13599 2431
rect 13541 2391 13599 2397
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15746 2428 15752 2440
rect 14967 2400 15752 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 12069 2363 12127 2369
rect 12069 2329 12081 2363
rect 12115 2329 12127 2363
rect 12434 2360 12440 2372
rect 12069 2323 12127 2329
rect 12406 2320 12440 2360
rect 12492 2320 12498 2372
rect 12805 2363 12863 2369
rect 12805 2329 12817 2363
rect 12851 2360 12863 2363
rect 14366 2360 14372 2372
rect 12851 2332 14372 2360
rect 12851 2329 12863 2332
rect 12805 2323 12863 2329
rect 14366 2320 14372 2332
rect 14424 2320 14430 2372
rect 12406 2292 12434 2320
rect 9508 2264 12434 2292
rect 12897 2295 12955 2301
rect 12897 2261 12909 2295
rect 12943 2292 12955 2295
rect 13998 2292 14004 2304
rect 12943 2264 14004 2292
rect 12943 2261 12955 2264
rect 12897 2255 12955 2261
rect 13998 2252 14004 2264
rect 14056 2252 14062 2304
rect 14476 2292 14504 2391
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2428 15899 2431
rect 16298 2428 16304 2440
rect 15887 2400 16304 2428
rect 15887 2397 15899 2400
rect 15841 2391 15899 2397
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 17512 2437 17540 2536
rect 22370 2496 22376 2508
rect 18432 2468 22376 2496
rect 18432 2437 18460 2468
rect 22370 2456 22376 2468
rect 22428 2456 22434 2508
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 18417 2391 18475 2397
rect 19150 2388 19156 2440
rect 19208 2428 19214 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19208 2400 19625 2428
rect 19208 2388 19214 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 20070 2428 20076 2440
rect 20031 2400 20076 2428
rect 19613 2391 19671 2397
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 20990 2428 20996 2440
rect 20951 2400 20996 2428
rect 20990 2388 20996 2400
rect 21048 2388 21054 2440
rect 22005 2431 22063 2437
rect 21192 2400 21956 2428
rect 15194 2360 15200 2372
rect 15155 2332 15200 2360
rect 15194 2320 15200 2332
rect 15252 2320 15258 2372
rect 16114 2360 16120 2372
rect 16075 2332 16120 2360
rect 16114 2320 16120 2332
rect 16172 2320 16178 2372
rect 17773 2363 17831 2369
rect 17773 2329 17785 2363
rect 17819 2360 17831 2363
rect 18506 2360 18512 2372
rect 17819 2332 18512 2360
rect 17819 2329 17831 2332
rect 17773 2323 17831 2329
rect 18506 2320 18512 2332
rect 18564 2320 18570 2372
rect 18693 2363 18751 2369
rect 18693 2329 18705 2363
rect 18739 2360 18751 2363
rect 20254 2360 20260 2372
rect 18739 2332 20260 2360
rect 18739 2329 18751 2332
rect 18693 2323 18751 2329
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 20349 2363 20407 2369
rect 20349 2329 20361 2363
rect 20395 2360 20407 2363
rect 21192 2360 21220 2400
rect 20395 2332 21220 2360
rect 21269 2363 21327 2369
rect 20395 2329 20407 2332
rect 20349 2323 20407 2329
rect 21269 2329 21281 2363
rect 21315 2329 21327 2363
rect 21928 2360 21956 2400
rect 22005 2397 22017 2431
rect 22051 2428 22063 2431
rect 22572 2428 22600 2536
rect 24210 2524 24216 2536
rect 24268 2524 24274 2576
rect 22925 2499 22983 2505
rect 22925 2465 22937 2499
rect 22971 2496 22983 2499
rect 24946 2496 24952 2508
rect 22971 2468 24952 2496
rect 22971 2465 22983 2468
rect 22925 2459 22983 2465
rect 24946 2456 24952 2468
rect 25004 2456 25010 2508
rect 22051 2400 22600 2428
rect 22649 2431 22707 2437
rect 22051 2397 22063 2400
rect 22005 2391 22063 2397
rect 22649 2397 22661 2431
rect 22695 2428 22707 2431
rect 23382 2428 23388 2440
rect 22695 2400 23388 2428
rect 22695 2397 22707 2400
rect 22649 2391 22707 2397
rect 23382 2388 23388 2400
rect 23440 2388 23446 2440
rect 23569 2431 23627 2437
rect 23569 2397 23581 2431
rect 23615 2428 23627 2431
rect 25148 2428 25176 2604
rect 27062 2592 27068 2604
rect 27120 2592 27126 2644
rect 41138 2632 41144 2644
rect 41099 2604 41144 2632
rect 41138 2592 41144 2604
rect 41196 2592 41202 2644
rect 44177 2635 44235 2641
rect 44177 2601 44189 2635
rect 44223 2632 44235 2635
rect 44634 2632 44640 2644
rect 44223 2604 44640 2632
rect 44223 2601 44235 2604
rect 44177 2595 44235 2601
rect 44634 2592 44640 2604
rect 44692 2592 44698 2644
rect 45094 2592 45100 2644
rect 45152 2632 45158 2644
rect 45278 2632 45284 2644
rect 45152 2604 45284 2632
rect 45152 2592 45158 2604
rect 45278 2592 45284 2604
rect 45336 2592 45342 2644
rect 45370 2592 45376 2644
rect 45428 2632 45434 2644
rect 45741 2635 45799 2641
rect 45741 2632 45753 2635
rect 45428 2604 45753 2632
rect 45428 2592 45434 2604
rect 45741 2601 45753 2604
rect 45787 2601 45799 2635
rect 46474 2632 46480 2644
rect 46435 2604 46480 2632
rect 45741 2595 45799 2601
rect 46474 2592 46480 2604
rect 46532 2592 46538 2644
rect 49050 2592 49056 2644
rect 49108 2632 49114 2644
rect 50525 2635 50583 2641
rect 50525 2632 50537 2635
rect 49108 2604 50537 2632
rect 49108 2592 49114 2604
rect 50525 2601 50537 2604
rect 50571 2601 50583 2635
rect 51442 2632 51448 2644
rect 51403 2604 51448 2632
rect 50525 2595 50583 2601
rect 51442 2592 51448 2604
rect 51500 2592 51506 2644
rect 53098 2632 53104 2644
rect 53059 2604 53104 2632
rect 53098 2592 53104 2604
rect 53156 2592 53162 2644
rect 57974 2592 57980 2644
rect 58032 2632 58038 2644
rect 58253 2635 58311 2641
rect 58253 2632 58265 2635
rect 58032 2604 58265 2632
rect 58032 2592 58038 2604
rect 58253 2601 58265 2604
rect 58299 2601 58311 2635
rect 58253 2595 58311 2601
rect 27890 2564 27896 2576
rect 25240 2536 27896 2564
rect 25240 2437 25268 2536
rect 27890 2524 27896 2536
rect 27948 2524 27954 2576
rect 36814 2524 36820 2576
rect 36872 2564 36878 2576
rect 45296 2564 45324 2592
rect 46198 2564 46204 2576
rect 36872 2536 40264 2564
rect 45296 2536 46204 2564
rect 36872 2524 36878 2536
rect 28074 2496 28080 2508
rect 26160 2468 28080 2496
rect 26160 2437 26188 2468
rect 28074 2456 28080 2468
rect 28132 2456 28138 2508
rect 29178 2456 29184 2508
rect 29236 2496 29242 2508
rect 29236 2468 31156 2496
rect 29236 2456 29242 2468
rect 23615 2400 25176 2428
rect 25225 2431 25283 2437
rect 23615 2397 23627 2400
rect 23569 2391 23627 2397
rect 25225 2397 25237 2431
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2397 26203 2431
rect 26145 2391 26203 2397
rect 26234 2388 26240 2440
rect 26292 2428 26298 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 26292 2400 27169 2428
rect 26292 2388 26298 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 28166 2388 28172 2440
rect 28224 2428 28230 2440
rect 28721 2431 28779 2437
rect 28721 2428 28733 2431
rect 28224 2400 28733 2428
rect 28224 2388 28230 2400
rect 28721 2397 28733 2400
rect 28767 2397 28779 2431
rect 28721 2391 28779 2397
rect 30098 2388 30104 2440
rect 30156 2428 30162 2440
rect 31128 2437 31156 2468
rect 31202 2456 31208 2508
rect 31260 2496 31266 2508
rect 33410 2496 33416 2508
rect 31260 2468 32352 2496
rect 33371 2468 33416 2496
rect 31260 2456 31266 2468
rect 32324 2437 32352 2468
rect 33410 2456 33416 2468
rect 33468 2456 33474 2508
rect 35986 2496 35992 2508
rect 35947 2468 35992 2496
rect 35986 2456 35992 2468
rect 36044 2456 36050 2508
rect 40236 2505 40264 2536
rect 46198 2524 46204 2536
rect 46256 2524 46262 2576
rect 51350 2564 51356 2576
rect 48792 2536 51356 2564
rect 38565 2499 38623 2505
rect 38565 2496 38577 2499
rect 37292 2468 38577 2496
rect 30193 2431 30251 2437
rect 30193 2428 30205 2431
rect 30156 2400 30205 2428
rect 30156 2388 30162 2400
rect 30193 2397 30205 2400
rect 30239 2397 30251 2431
rect 30193 2391 30251 2397
rect 31113 2431 31171 2437
rect 31113 2397 31125 2431
rect 31159 2397 31171 2431
rect 31113 2391 31171 2397
rect 32309 2431 32367 2437
rect 32309 2397 32321 2431
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33042 2388 33048 2440
rect 33100 2428 33106 2440
rect 33229 2431 33287 2437
rect 33229 2428 33241 2431
rect 33100 2400 33241 2428
rect 33100 2388 33106 2400
rect 33229 2397 33241 2400
rect 33275 2397 33287 2431
rect 33229 2391 33287 2397
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35710 2388 35716 2440
rect 35768 2428 35774 2440
rect 35805 2431 35863 2437
rect 35805 2428 35817 2431
rect 35768 2400 35817 2428
rect 35768 2388 35774 2400
rect 35805 2397 35817 2400
rect 35851 2397 35863 2431
rect 37292 2428 37320 2468
rect 38565 2465 38577 2468
rect 38611 2465 38623 2499
rect 38565 2459 38623 2465
rect 40221 2499 40279 2505
rect 40221 2465 40233 2499
rect 40267 2465 40279 2499
rect 48792 2496 48820 2536
rect 51350 2524 51356 2536
rect 51408 2524 51414 2576
rect 48958 2496 48964 2508
rect 40221 2459 40279 2465
rect 43916 2468 48820 2496
rect 48919 2468 48964 2496
rect 35805 2391 35863 2397
rect 35912 2400 37320 2428
rect 37461 2431 37519 2437
rect 23474 2360 23480 2372
rect 21928 2332 23480 2360
rect 21269 2323 21327 2329
rect 18598 2292 18604 2304
rect 14476 2264 18604 2292
rect 18598 2252 18604 2264
rect 18656 2252 18662 2304
rect 21284 2292 21312 2323
rect 23474 2320 23480 2332
rect 23532 2320 23538 2372
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 25501 2363 25559 2369
rect 23891 2332 25268 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 25240 2304 25268 2332
rect 25501 2329 25513 2363
rect 25547 2360 25559 2363
rect 25774 2360 25780 2372
rect 25547 2332 25780 2360
rect 25547 2329 25559 2332
rect 25501 2323 25559 2329
rect 25774 2320 25780 2332
rect 25832 2320 25838 2372
rect 26421 2363 26479 2369
rect 26421 2329 26433 2363
rect 26467 2360 26479 2363
rect 26602 2360 26608 2372
rect 26467 2332 26608 2360
rect 26467 2329 26479 2332
rect 26421 2323 26479 2329
rect 26602 2320 26608 2332
rect 26660 2320 26666 2372
rect 26878 2320 26884 2372
rect 26936 2360 26942 2372
rect 27433 2363 27491 2369
rect 27433 2360 27445 2363
rect 26936 2332 27445 2360
rect 26936 2320 26942 2332
rect 27433 2329 27445 2332
rect 27479 2329 27491 2363
rect 27433 2323 27491 2329
rect 28997 2363 29055 2369
rect 28997 2329 29009 2363
rect 29043 2360 29055 2363
rect 29914 2360 29920 2372
rect 29043 2332 29920 2360
rect 29043 2329 29055 2332
rect 28997 2323 29055 2329
rect 29914 2320 29920 2332
rect 29972 2320 29978 2372
rect 30466 2360 30472 2372
rect 30427 2332 30472 2360
rect 30466 2320 30472 2332
rect 30524 2320 30530 2372
rect 31018 2320 31024 2372
rect 31076 2360 31082 2372
rect 31389 2363 31447 2369
rect 31389 2360 31401 2363
rect 31076 2332 31401 2360
rect 31076 2320 31082 2332
rect 31389 2329 31401 2332
rect 31435 2329 31447 2363
rect 31389 2323 31447 2329
rect 32585 2363 32643 2369
rect 32585 2329 32597 2363
rect 32631 2329 32643 2363
rect 32585 2323 32643 2329
rect 24118 2292 24124 2304
rect 21284 2264 24124 2292
rect 24118 2252 24124 2264
rect 24176 2252 24182 2304
rect 25222 2252 25228 2304
rect 25280 2252 25286 2304
rect 28077 2295 28135 2301
rect 28077 2261 28089 2295
rect 28123 2292 28135 2295
rect 29638 2292 29644 2304
rect 28123 2264 29644 2292
rect 28123 2261 28135 2264
rect 28077 2255 28135 2261
rect 29638 2252 29644 2264
rect 29696 2252 29702 2304
rect 31294 2252 31300 2304
rect 31352 2292 31358 2304
rect 32600 2292 32628 2323
rect 32674 2320 32680 2372
rect 32732 2360 32738 2372
rect 35161 2363 35219 2369
rect 35161 2360 35173 2363
rect 32732 2332 35173 2360
rect 32732 2320 32738 2332
rect 35161 2329 35173 2332
rect 35207 2329 35219 2363
rect 35161 2323 35219 2329
rect 35434 2320 35440 2372
rect 35492 2360 35498 2372
rect 35912 2360 35940 2400
rect 37461 2397 37473 2431
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 38381 2431 38439 2437
rect 38381 2397 38393 2431
rect 38427 2428 38439 2431
rect 39390 2428 39396 2440
rect 38427 2400 39396 2428
rect 38427 2397 38439 2400
rect 38381 2391 38439 2397
rect 35492 2332 35940 2360
rect 35492 2320 35498 2332
rect 37274 2320 37280 2372
rect 37332 2360 37338 2372
rect 37476 2360 37504 2391
rect 39390 2388 39396 2400
rect 39448 2388 39454 2440
rect 39482 2388 39488 2440
rect 39540 2428 39546 2440
rect 40037 2431 40095 2437
rect 40037 2428 40049 2431
rect 39540 2400 40049 2428
rect 39540 2388 39546 2400
rect 40037 2397 40049 2400
rect 40083 2397 40095 2431
rect 40037 2391 40095 2397
rect 40126 2388 40132 2440
rect 40184 2428 40190 2440
rect 41049 2431 41107 2437
rect 41049 2428 41061 2431
rect 40184 2400 41061 2428
rect 40184 2388 40190 2400
rect 41049 2397 41061 2400
rect 41095 2397 41107 2431
rect 41049 2391 41107 2397
rect 41138 2388 41144 2440
rect 41196 2428 41202 2440
rect 42613 2431 42671 2437
rect 42613 2428 42625 2431
rect 41196 2400 42625 2428
rect 41196 2388 41202 2400
rect 42613 2397 42625 2400
rect 42659 2397 42671 2431
rect 43530 2428 43536 2440
rect 43491 2400 43536 2428
rect 42613 2391 42671 2397
rect 43530 2388 43536 2400
rect 43588 2388 43594 2440
rect 43681 2431 43739 2437
rect 43681 2397 43693 2431
rect 43727 2428 43739 2431
rect 43916 2428 43944 2468
rect 48958 2456 48964 2468
rect 49016 2456 49022 2508
rect 54754 2496 54760 2508
rect 54715 2468 54760 2496
rect 54754 2456 54760 2468
rect 54812 2456 54818 2508
rect 43727 2400 43944 2428
rect 44039 2431 44097 2437
rect 43727 2397 43739 2400
rect 43681 2391 43739 2397
rect 44039 2397 44051 2431
rect 44085 2428 44097 2431
rect 44266 2428 44272 2440
rect 44085 2400 44272 2428
rect 44085 2397 44097 2400
rect 44039 2391 44097 2397
rect 44266 2388 44272 2400
rect 44324 2388 44330 2440
rect 45186 2428 45192 2440
rect 45147 2400 45192 2428
rect 45186 2388 45192 2400
rect 45244 2388 45250 2440
rect 45278 2388 45284 2440
rect 45336 2428 45342 2440
rect 45373 2431 45431 2437
rect 45373 2428 45385 2431
rect 45336 2400 45385 2428
rect 45336 2388 45342 2400
rect 45373 2397 45385 2400
rect 45419 2397 45431 2431
rect 45373 2391 45431 2397
rect 45554 2388 45560 2440
rect 45612 2437 45618 2440
rect 45612 2428 45620 2437
rect 46658 2428 46664 2440
rect 45612 2400 45657 2428
rect 46216 2400 46664 2428
rect 45612 2391 45620 2400
rect 45612 2388 45618 2391
rect 37332 2332 37504 2360
rect 37737 2363 37795 2369
rect 37332 2320 37338 2332
rect 37737 2329 37749 2363
rect 37783 2329 37795 2363
rect 37737 2323 37795 2329
rect 31352 2264 32628 2292
rect 31352 2252 31358 2264
rect 34330 2252 34336 2304
rect 34388 2292 34394 2304
rect 37752 2292 37780 2323
rect 40494 2320 40500 2372
rect 40552 2360 40558 2372
rect 42889 2363 42947 2369
rect 42889 2360 42901 2363
rect 40552 2332 42901 2360
rect 40552 2320 40558 2332
rect 42889 2329 42901 2332
rect 42935 2329 42947 2363
rect 42889 2323 42947 2329
rect 43346 2320 43352 2372
rect 43404 2360 43410 2372
rect 43809 2363 43867 2369
rect 43809 2360 43821 2363
rect 43404 2332 43821 2360
rect 43404 2320 43410 2332
rect 43809 2329 43821 2332
rect 43855 2329 43867 2363
rect 43809 2323 43867 2329
rect 43901 2363 43959 2369
rect 43901 2329 43913 2363
rect 43947 2360 43959 2363
rect 44726 2360 44732 2372
rect 43947 2332 44732 2360
rect 43947 2329 43959 2332
rect 43901 2323 43959 2329
rect 44726 2320 44732 2332
rect 44784 2320 44790 2372
rect 45465 2363 45523 2369
rect 45465 2329 45477 2363
rect 45511 2360 45523 2363
rect 46216 2360 46244 2400
rect 46658 2388 46664 2400
rect 46716 2388 46722 2440
rect 48038 2388 48044 2440
rect 48096 2428 48102 2440
rect 48685 2431 48743 2437
rect 48685 2428 48697 2431
rect 48096 2400 48697 2428
rect 48096 2388 48102 2400
rect 48685 2397 48697 2400
rect 48731 2397 48743 2431
rect 48685 2391 48743 2397
rect 51166 2388 51172 2440
rect 51224 2428 51230 2440
rect 52917 2431 52975 2437
rect 52917 2428 52929 2431
rect 51224 2400 52929 2428
rect 51224 2388 51230 2400
rect 52917 2397 52929 2400
rect 52963 2397 52975 2431
rect 52917 2391 52975 2397
rect 53650 2388 53656 2440
rect 53708 2428 53714 2440
rect 56321 2431 56379 2437
rect 56321 2428 56333 2431
rect 53708 2400 56333 2428
rect 53708 2388 53714 2400
rect 56321 2397 56333 2400
rect 56367 2397 56379 2431
rect 56321 2391 56379 2397
rect 57057 2431 57115 2437
rect 57057 2397 57069 2431
rect 57103 2428 57115 2431
rect 57238 2428 57244 2440
rect 57103 2400 57244 2428
rect 57103 2397 57115 2400
rect 57057 2391 57115 2397
rect 57238 2388 57244 2400
rect 57296 2388 57302 2440
rect 58158 2428 58164 2440
rect 58119 2400 58164 2428
rect 58158 2388 58164 2400
rect 58216 2388 58222 2440
rect 45511 2332 46244 2360
rect 46385 2363 46443 2369
rect 45511 2329 45523 2332
rect 45465 2323 45523 2329
rect 46385 2329 46397 2363
rect 46431 2329 46443 2363
rect 46385 2323 46443 2329
rect 34388 2264 37780 2292
rect 34388 2252 34394 2264
rect 42610 2252 42616 2304
rect 42668 2292 42674 2304
rect 46400 2292 46428 2323
rect 47578 2320 47584 2372
rect 47636 2360 47642 2372
rect 47857 2363 47915 2369
rect 47857 2360 47869 2363
rect 47636 2332 47869 2360
rect 47636 2320 47642 2332
rect 47857 2329 47869 2332
rect 47903 2329 47915 2363
rect 47857 2323 47915 2329
rect 48958 2320 48964 2372
rect 49016 2360 49022 2372
rect 50433 2363 50491 2369
rect 50433 2360 50445 2363
rect 49016 2332 50445 2360
rect 49016 2320 49022 2332
rect 50433 2329 50445 2332
rect 50479 2329 50491 2363
rect 51350 2360 51356 2372
rect 51311 2332 51356 2360
rect 50433 2323 50491 2329
rect 51350 2320 51356 2332
rect 51408 2320 51414 2372
rect 53926 2320 53932 2372
rect 53984 2360 53990 2372
rect 54021 2363 54079 2369
rect 54021 2360 54033 2363
rect 53984 2332 54033 2360
rect 53984 2320 53990 2332
rect 54021 2329 54033 2332
rect 54067 2329 54079 2363
rect 55585 2363 55643 2369
rect 55585 2360 55597 2363
rect 54021 2323 54079 2329
rect 55186 2332 55597 2360
rect 47946 2292 47952 2304
rect 42668 2264 46428 2292
rect 47907 2264 47952 2292
rect 42668 2252 42674 2264
rect 47946 2252 47952 2264
rect 48004 2252 48010 2304
rect 52822 2252 52828 2304
rect 52880 2292 52886 2304
rect 55186 2292 55214 2332
rect 55585 2329 55597 2332
rect 55631 2329 55643 2363
rect 57330 2360 57336 2372
rect 57291 2332 57336 2360
rect 55585 2323 55643 2329
rect 57330 2320 57336 2332
rect 57388 2320 57394 2372
rect 55674 2292 55680 2304
rect 52880 2264 55214 2292
rect 55635 2264 55680 2292
rect 52880 2252 52886 2264
rect 55674 2252 55680 2264
rect 55732 2252 55738 2304
rect 56410 2292 56416 2304
rect 56371 2264 56416 2292
rect 56410 2252 56416 2264
rect 56468 2252 56474 2304
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 9398 2048 9404 2100
rect 9456 2088 9462 2100
rect 12710 2088 12716 2100
rect 9456 2060 12716 2088
rect 9456 2048 9462 2060
rect 12710 2048 12716 2060
rect 12768 2048 12774 2100
rect 15194 2048 15200 2100
rect 15252 2088 15258 2100
rect 19702 2088 19708 2100
rect 15252 2060 19708 2088
rect 15252 2048 15258 2060
rect 19702 2048 19708 2060
rect 19760 2048 19766 2100
rect 20990 2048 20996 2100
rect 21048 2088 21054 2100
rect 24026 2088 24032 2100
rect 21048 2060 24032 2088
rect 21048 2048 21054 2060
rect 24026 2048 24032 2060
rect 24084 2048 24090 2100
rect 45186 2048 45192 2100
rect 45244 2088 45250 2100
rect 55674 2088 55680 2100
rect 45244 2060 55680 2088
rect 45244 2048 45250 2060
rect 55674 2048 55680 2060
rect 55732 2048 55738 2100
rect 1578 1980 1584 2032
rect 1636 2020 1642 2032
rect 1636 1992 22094 2020
rect 1636 1980 1642 1992
rect 7006 1912 7012 1964
rect 7064 1952 7070 1964
rect 11514 1952 11520 1964
rect 7064 1924 11520 1952
rect 7064 1912 7070 1924
rect 11514 1912 11520 1924
rect 11572 1912 11578 1964
rect 12802 1912 12808 1964
rect 12860 1952 12866 1964
rect 12860 1924 17816 1952
rect 12860 1912 12866 1924
rect 5166 1844 5172 1896
rect 5224 1884 5230 1896
rect 17678 1884 17684 1896
rect 5224 1856 17684 1884
rect 5224 1844 5230 1856
rect 17678 1844 17684 1856
rect 17736 1844 17742 1896
rect 17788 1884 17816 1924
rect 18506 1912 18512 1964
rect 18564 1952 18570 1964
rect 21910 1952 21916 1964
rect 18564 1924 21916 1952
rect 18564 1912 18570 1924
rect 21910 1912 21916 1924
rect 21968 1912 21974 1964
rect 22066 1952 22094 1992
rect 22370 1980 22376 2032
rect 22428 2020 22434 2032
rect 31662 2020 31668 2032
rect 22428 1992 31668 2020
rect 22428 1980 22434 1992
rect 31662 1980 31668 1992
rect 31720 1980 31726 2032
rect 38102 1980 38108 2032
rect 38160 2020 38166 2032
rect 56410 2020 56416 2032
rect 38160 1992 56416 2020
rect 38160 1980 38166 1992
rect 56410 1980 56416 1992
rect 56468 1980 56474 2032
rect 28350 1952 28356 1964
rect 22066 1924 28356 1952
rect 28350 1912 28356 1924
rect 28408 1912 28414 1964
rect 40494 1952 40500 1964
rect 35866 1924 40500 1952
rect 31202 1884 31208 1896
rect 17788 1856 31208 1884
rect 31202 1844 31208 1856
rect 31260 1844 31266 1896
rect 9674 1776 9680 1828
rect 9732 1816 9738 1828
rect 14550 1816 14556 1828
rect 9732 1788 14556 1816
rect 9732 1776 9738 1788
rect 14550 1776 14556 1788
rect 14608 1776 14614 1828
rect 20622 1776 20628 1828
rect 20680 1816 20686 1828
rect 35866 1816 35894 1924
rect 40494 1912 40500 1924
rect 40552 1912 40558 1964
rect 20680 1788 35894 1816
rect 20680 1776 20686 1788
rect 7742 1708 7748 1760
rect 7800 1748 7806 1760
rect 12618 1748 12624 1760
rect 7800 1720 12624 1748
rect 7800 1708 7806 1720
rect 12618 1708 12624 1720
rect 12676 1708 12682 1760
rect 16114 1708 16120 1760
rect 16172 1748 16178 1760
rect 20530 1748 20536 1760
rect 16172 1720 20536 1748
rect 16172 1708 16178 1720
rect 20530 1708 20536 1720
rect 20588 1708 20594 1760
rect 19242 1640 19248 1692
rect 19300 1680 19306 1692
rect 26234 1680 26240 1692
rect 19300 1652 26240 1680
rect 19300 1640 19306 1652
rect 26234 1640 26240 1652
rect 26292 1640 26298 1692
rect 9306 1504 9312 1556
rect 9364 1544 9370 1556
rect 10870 1544 10876 1556
rect 9364 1516 10876 1544
rect 9364 1504 9370 1516
rect 10870 1504 10876 1516
rect 10928 1504 10934 1556
rect 9858 1436 9864 1488
rect 9916 1476 9922 1488
rect 12250 1476 12256 1488
rect 9916 1448 12256 1476
rect 9916 1436 9922 1448
rect 12250 1436 12256 1448
rect 12308 1436 12314 1488
rect 33226 1436 33232 1488
rect 33284 1476 33290 1488
rect 33594 1476 33600 1488
rect 33284 1448 33600 1476
rect 33284 1436 33290 1448
rect 33594 1436 33600 1448
rect 33652 1436 33658 1488
rect 6822 1368 6828 1420
rect 6880 1408 6886 1420
rect 7558 1408 7564 1420
rect 6880 1380 7564 1408
rect 6880 1368 6886 1380
rect 7558 1368 7564 1380
rect 7616 1368 7622 1420
rect 8478 1368 8484 1420
rect 8536 1408 8542 1420
rect 11146 1408 11152 1420
rect 8536 1380 11152 1408
rect 8536 1368 8542 1380
rect 11146 1368 11152 1380
rect 11204 1368 11210 1420
rect 12434 1368 12440 1420
rect 12492 1408 12498 1420
rect 13906 1408 13912 1420
rect 12492 1380 13912 1408
rect 12492 1368 12498 1380
rect 13906 1368 13912 1380
rect 13964 1368 13970 1420
rect 14366 1368 14372 1420
rect 14424 1408 14430 1420
rect 15286 1408 15292 1420
rect 14424 1380 15292 1408
rect 14424 1368 14430 1380
rect 15286 1368 15292 1380
rect 15344 1368 15350 1420
rect 34054 1368 34060 1420
rect 34112 1408 34118 1420
rect 35894 1408 35900 1420
rect 34112 1380 35900 1408
rect 34112 1368 34118 1380
rect 35894 1368 35900 1380
rect 35952 1368 35958 1420
rect 50338 1368 50344 1420
rect 50396 1408 50402 1420
rect 51350 1408 51356 1420
rect 50396 1380 51356 1408
rect 50396 1368 50402 1380
rect 51350 1368 51356 1380
rect 51408 1368 51414 1420
rect 50706 1300 50712 1352
rect 50764 1340 50770 1352
rect 56502 1340 56508 1352
rect 50764 1312 56508 1340
rect 50764 1300 50770 1312
rect 56502 1300 56508 1312
rect 56560 1300 56566 1352
<< via1 >>
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 6184 61276 6236 61328
rect 17132 61276 17184 61328
rect 21732 61276 21784 61328
rect 2780 61208 2832 61260
rect 44456 61208 44508 61260
rect 56784 61208 56836 61260
rect 4620 61140 4672 61192
rect 5080 61183 5132 61192
rect 5080 61149 5089 61183
rect 5089 61149 5123 61183
rect 5123 61149 5132 61183
rect 5080 61140 5132 61149
rect 5816 61183 5868 61192
rect 5816 61149 5825 61183
rect 5825 61149 5859 61183
rect 5859 61149 5868 61183
rect 5816 61140 5868 61149
rect 6736 61183 6788 61192
rect 6736 61149 6745 61183
rect 6745 61149 6779 61183
rect 6779 61149 6788 61183
rect 6736 61140 6788 61149
rect 7564 61183 7616 61192
rect 7564 61149 7573 61183
rect 7573 61149 7607 61183
rect 7607 61149 7616 61183
rect 7564 61140 7616 61149
rect 7840 61183 7892 61192
rect 7840 61149 7849 61183
rect 7849 61149 7883 61183
rect 7883 61149 7892 61183
rect 7840 61140 7892 61149
rect 9680 61140 9732 61192
rect 10232 61183 10284 61192
rect 10232 61149 10241 61183
rect 10241 61149 10275 61183
rect 10275 61149 10284 61183
rect 10232 61140 10284 61149
rect 11152 61140 11204 61192
rect 12440 61183 12492 61192
rect 12440 61149 12449 61183
rect 12449 61149 12483 61183
rect 12483 61149 12492 61183
rect 12440 61140 12492 61149
rect 13268 61183 13320 61192
rect 13268 61149 13277 61183
rect 13277 61149 13311 61183
rect 13311 61149 13320 61183
rect 13268 61140 13320 61149
rect 14372 61183 14424 61192
rect 14372 61149 14381 61183
rect 14381 61149 14415 61183
rect 14415 61149 14424 61183
rect 14372 61140 14424 61149
rect 15384 61183 15436 61192
rect 15384 61149 15393 61183
rect 15393 61149 15427 61183
rect 15427 61149 15436 61183
rect 15384 61140 15436 61149
rect 16120 61183 16172 61192
rect 16120 61149 16129 61183
rect 16129 61149 16163 61183
rect 16163 61149 16172 61183
rect 16120 61140 16172 61149
rect 17224 61183 17276 61192
rect 17224 61149 17233 61183
rect 17233 61149 17267 61183
rect 17267 61149 17276 61183
rect 17224 61140 17276 61149
rect 17960 61183 18012 61192
rect 17960 61149 17969 61183
rect 17969 61149 18003 61183
rect 18003 61149 18012 61183
rect 17960 61140 18012 61149
rect 18696 61183 18748 61192
rect 18696 61149 18705 61183
rect 18705 61149 18739 61183
rect 18739 61149 18748 61183
rect 18696 61140 18748 61149
rect 19800 61183 19852 61192
rect 19800 61149 19809 61183
rect 19809 61149 19843 61183
rect 19843 61149 19852 61183
rect 19800 61140 19852 61149
rect 20720 61140 20772 61192
rect 21272 61183 21324 61192
rect 21272 61149 21281 61183
rect 21281 61149 21315 61183
rect 21315 61149 21324 61183
rect 21272 61140 21324 61149
rect 22376 61183 22428 61192
rect 22376 61149 22385 61183
rect 22385 61149 22419 61183
rect 22419 61149 22428 61183
rect 22376 61140 22428 61149
rect 23112 61183 23164 61192
rect 23112 61149 23121 61183
rect 23121 61149 23155 61183
rect 23155 61149 23164 61183
rect 23112 61140 23164 61149
rect 23848 61183 23900 61192
rect 23848 61149 23857 61183
rect 23857 61149 23891 61183
rect 23891 61149 23900 61183
rect 23848 61140 23900 61149
rect 25136 61140 25188 61192
rect 26056 61183 26108 61192
rect 26056 61149 26065 61183
rect 26065 61149 26099 61183
rect 26099 61149 26108 61183
rect 26056 61140 26108 61149
rect 27528 61183 27580 61192
rect 27528 61149 27537 61183
rect 27537 61149 27571 61183
rect 27571 61149 27580 61183
rect 27528 61140 27580 61149
rect 28356 61183 28408 61192
rect 28356 61149 28365 61183
rect 28365 61149 28399 61183
rect 28399 61149 28408 61183
rect 28356 61140 28408 61149
rect 29000 61140 29052 61192
rect 31024 61140 31076 61192
rect 31760 61140 31812 61192
rect 32496 61140 32548 61192
rect 33232 61140 33284 61192
rect 34704 61140 34756 61192
rect 35900 61183 35952 61192
rect 35900 61149 35909 61183
rect 35909 61149 35943 61183
rect 35943 61149 35952 61183
rect 35900 61140 35952 61149
rect 37280 61140 37332 61192
rect 37648 61140 37700 61192
rect 38384 61140 38436 61192
rect 40040 61140 40092 61192
rect 40960 61140 41012 61192
rect 42064 61140 42116 61192
rect 42800 61140 42852 61192
rect 44180 61140 44232 61192
rect 44548 61140 44600 61192
rect 45560 61140 45612 61192
rect 46112 61140 46164 61192
rect 47216 61140 47268 61192
rect 48320 61140 48372 61192
rect 48688 61140 48740 61192
rect 51080 61183 51132 61192
rect 51080 61149 51089 61183
rect 51089 61149 51123 61183
rect 51123 61149 51132 61183
rect 51080 61140 51132 61149
rect 52000 61183 52052 61192
rect 52000 61149 52009 61183
rect 52009 61149 52043 61183
rect 52043 61149 52052 61183
rect 52000 61140 52052 61149
rect 53196 61183 53248 61192
rect 53196 61149 53205 61183
rect 53205 61149 53239 61183
rect 53239 61149 53248 61183
rect 53196 61140 53248 61149
rect 54208 61183 54260 61192
rect 54208 61149 54217 61183
rect 54217 61149 54251 61183
rect 54251 61149 54260 61183
rect 54208 61140 54260 61149
rect 56140 61183 56192 61192
rect 56140 61149 56149 61183
rect 56149 61149 56183 61183
rect 56183 61149 56192 61183
rect 56140 61140 56192 61149
rect 57520 61140 57572 61192
rect 1676 61115 1728 61124
rect 1676 61081 1685 61115
rect 1685 61081 1719 61115
rect 1719 61081 1728 61115
rect 1676 61072 1728 61081
rect 4896 61072 4948 61124
rect 7656 61072 7708 61124
rect 13544 61115 13596 61124
rect 13544 61081 13553 61115
rect 13553 61081 13587 61115
rect 13587 61081 13596 61115
rect 13544 61072 13596 61081
rect 15660 61072 15712 61124
rect 16396 61072 16448 61124
rect 18144 61115 18196 61124
rect 18144 61081 18153 61115
rect 18153 61081 18187 61115
rect 18187 61081 18196 61115
rect 18144 61072 18196 61081
rect 20352 61072 20404 61124
rect 31668 61072 31720 61124
rect 37740 61115 37792 61124
rect 37740 61081 37749 61115
rect 37749 61081 37783 61115
rect 37783 61081 37792 61115
rect 37740 61072 37792 61081
rect 39488 61072 39540 61124
rect 46940 61115 46992 61124
rect 5172 61047 5224 61056
rect 5172 61013 5181 61047
rect 5181 61013 5215 61047
rect 5215 61013 5224 61047
rect 5172 61004 5224 61013
rect 5908 61047 5960 61056
rect 5908 61013 5917 61047
rect 5917 61013 5951 61047
rect 5951 61013 5960 61047
rect 5908 61004 5960 61013
rect 6920 61004 6972 61056
rect 10324 61047 10376 61056
rect 10324 61013 10333 61047
rect 10333 61013 10367 61047
rect 10367 61013 10376 61047
rect 10324 61004 10376 61013
rect 11980 61004 12032 61056
rect 12532 61047 12584 61056
rect 12532 61013 12541 61047
rect 12541 61013 12575 61047
rect 12575 61013 12584 61047
rect 12532 61004 12584 61013
rect 14464 61047 14516 61056
rect 14464 61013 14473 61047
rect 14473 61013 14507 61047
rect 14507 61013 14516 61047
rect 14464 61004 14516 61013
rect 16580 61004 16632 61056
rect 18512 61004 18564 61056
rect 20812 61004 20864 61056
rect 22284 61004 22336 61056
rect 22928 61004 22980 61056
rect 23940 61047 23992 61056
rect 23940 61013 23949 61047
rect 23949 61013 23983 61047
rect 23983 61013 23992 61047
rect 23940 61004 23992 61013
rect 25136 61004 25188 61056
rect 27620 61047 27672 61056
rect 27620 61013 27629 61047
rect 27629 61013 27663 61047
rect 27663 61013 27672 61047
rect 27620 61004 27672 61013
rect 28540 61047 28592 61056
rect 28540 61013 28549 61047
rect 28549 61013 28583 61047
rect 28583 61013 28592 61047
rect 28540 61004 28592 61013
rect 30012 61004 30064 61056
rect 31024 61004 31076 61056
rect 31944 61004 31996 61056
rect 33232 61047 33284 61056
rect 33232 61013 33241 61047
rect 33241 61013 33275 61047
rect 33275 61013 33284 61047
rect 33232 61004 33284 61013
rect 33324 61004 33376 61056
rect 35072 61047 35124 61056
rect 35072 61013 35081 61047
rect 35081 61013 35115 61047
rect 35115 61013 35124 61047
rect 35072 61004 35124 61013
rect 35992 61047 36044 61056
rect 35992 61013 36001 61047
rect 36001 61013 36035 61047
rect 36035 61013 36044 61047
rect 35992 61004 36044 61013
rect 37280 61004 37332 61056
rect 39764 61004 39816 61056
rect 40224 61047 40276 61056
rect 40224 61013 40233 61047
rect 40233 61013 40267 61047
rect 40267 61013 40276 61047
rect 40224 61004 40276 61013
rect 40960 61047 41012 61056
rect 40960 61013 40969 61047
rect 40969 61013 41003 61047
rect 41003 61013 41012 61047
rect 40960 61004 41012 61013
rect 41052 61004 41104 61056
rect 42064 61004 42116 61056
rect 42800 61047 42852 61056
rect 42800 61013 42809 61047
rect 42809 61013 42843 61047
rect 42843 61013 42852 61047
rect 42800 61004 42852 61013
rect 43720 61047 43772 61056
rect 43720 61013 43729 61047
rect 43729 61013 43763 61047
rect 43763 61013 43772 61047
rect 43720 61004 43772 61013
rect 44272 61004 44324 61056
rect 45376 61047 45428 61056
rect 45376 61013 45385 61047
rect 45385 61013 45419 61047
rect 45419 61013 45428 61047
rect 45376 61004 45428 61013
rect 46112 61047 46164 61056
rect 46112 61013 46121 61047
rect 46121 61013 46155 61047
rect 46155 61013 46164 61047
rect 46112 61004 46164 61013
rect 46940 61081 46949 61115
rect 46949 61081 46983 61115
rect 46983 61081 46992 61115
rect 46940 61072 46992 61081
rect 54392 61115 54444 61124
rect 54392 61081 54401 61115
rect 54401 61081 54435 61115
rect 54435 61081 54444 61115
rect 54392 61072 54444 61081
rect 56416 61115 56468 61124
rect 56416 61081 56425 61115
rect 56425 61081 56459 61115
rect 56459 61081 56468 61115
rect 56416 61072 56468 61081
rect 47952 61047 48004 61056
rect 47952 61013 47961 61047
rect 47961 61013 47995 61047
rect 47995 61013 48004 61047
rect 47952 61004 48004 61013
rect 48688 61047 48740 61056
rect 48688 61013 48697 61047
rect 48697 61013 48731 61047
rect 48731 61013 48740 61047
rect 48688 61004 48740 61013
rect 51172 61047 51224 61056
rect 51172 61013 51181 61047
rect 51181 61013 51215 61047
rect 51215 61013 51224 61047
rect 51172 61004 51224 61013
rect 52092 61047 52144 61056
rect 52092 61013 52101 61047
rect 52101 61013 52135 61047
rect 52135 61013 52144 61047
rect 52092 61004 52144 61013
rect 56876 61004 56928 61056
rect 58164 61004 58216 61056
rect 19574 60902 19626 60954
rect 19638 60902 19690 60954
rect 19702 60902 19754 60954
rect 19766 60902 19818 60954
rect 19830 60902 19882 60954
rect 50294 60902 50346 60954
rect 50358 60902 50410 60954
rect 50422 60902 50474 60954
rect 50486 60902 50538 60954
rect 50550 60902 50602 60954
rect 5908 60800 5960 60852
rect 23480 60800 23532 60852
rect 26884 60800 26936 60852
rect 40960 60800 41012 60852
rect 1676 60775 1728 60784
rect 1676 60741 1685 60775
rect 1685 60741 1719 60775
rect 1719 60741 1728 60775
rect 1676 60732 1728 60741
rect 3240 60775 3292 60784
rect 3240 60741 3249 60775
rect 3249 60741 3283 60775
rect 3283 60741 3292 60775
rect 3240 60732 3292 60741
rect 3976 60775 4028 60784
rect 3976 60741 3985 60775
rect 3985 60741 4019 60775
rect 4019 60741 4028 60775
rect 3976 60732 4028 60741
rect 8300 60732 8352 60784
rect 9128 60775 9180 60784
rect 9128 60741 9137 60775
rect 9137 60741 9171 60775
rect 9171 60741 9180 60775
rect 9128 60732 9180 60741
rect 12072 60775 12124 60784
rect 12072 60741 12081 60775
rect 12081 60741 12115 60775
rect 12115 60741 12124 60775
rect 12072 60732 12124 60741
rect 14832 60732 14884 60784
rect 19340 60732 19392 60784
rect 24584 60775 24636 60784
rect 24584 60741 24593 60775
rect 24593 60741 24627 60775
rect 24627 60741 24636 60775
rect 24584 60732 24636 60741
rect 33968 60732 34020 60784
rect 36360 60775 36412 60784
rect 36360 60741 36369 60775
rect 36369 60741 36403 60775
rect 36403 60741 36412 60775
rect 36360 60732 36412 60741
rect 46664 60775 46716 60784
rect 46664 60741 46673 60775
rect 46673 60741 46707 60775
rect 46707 60741 46716 60775
rect 46664 60732 46716 60741
rect 50160 60732 50212 60784
rect 52460 60732 52512 60784
rect 54760 60775 54812 60784
rect 54760 60741 54769 60775
rect 54769 60741 54803 60775
rect 54803 60741 54812 60775
rect 54760 60732 54812 60741
rect 55496 60775 55548 60784
rect 55496 60741 55505 60775
rect 55505 60741 55539 60775
rect 55539 60741 55548 60775
rect 55496 60732 55548 60741
rect 58256 60800 58308 60852
rect 57796 60732 57848 60784
rect 26608 60664 26660 60716
rect 29644 60707 29696 60716
rect 29644 60673 29653 60707
rect 29653 60673 29687 60707
rect 29687 60673 29696 60707
rect 29644 60664 29696 60673
rect 30288 60664 30340 60716
rect 41328 60664 41380 60716
rect 49516 60707 49568 60716
rect 49516 60673 49525 60707
rect 49525 60673 49559 60707
rect 49559 60673 49568 60707
rect 49516 60664 49568 60673
rect 56140 60707 56192 60716
rect 56140 60673 56149 60707
rect 56149 60673 56183 60707
rect 56183 60673 56192 60707
rect 56140 60664 56192 60673
rect 15108 60596 15160 60648
rect 56324 60639 56376 60648
rect 56324 60605 56333 60639
rect 56333 60605 56367 60639
rect 56367 60605 56376 60639
rect 56324 60596 56376 60605
rect 4804 60528 4856 60580
rect 8576 60571 8628 60580
rect 8576 60537 8585 60571
rect 8585 60537 8619 60571
rect 8619 60537 8628 60571
rect 8576 60528 8628 60537
rect 16028 60528 16080 60580
rect 20444 60528 20496 60580
rect 25320 60528 25372 60580
rect 1952 60503 2004 60512
rect 1952 60469 1961 60503
rect 1961 60469 1995 60503
rect 1995 60469 2004 60503
rect 1952 60460 2004 60469
rect 3332 60503 3384 60512
rect 3332 60469 3341 60503
rect 3341 60469 3375 60503
rect 3375 60469 3384 60503
rect 3332 60460 3384 60469
rect 12164 60503 12216 60512
rect 12164 60469 12173 60503
rect 12173 60469 12207 60503
rect 12207 60469 12216 60503
rect 12164 60460 12216 60469
rect 27344 60503 27396 60512
rect 27344 60469 27353 60503
rect 27353 60469 27387 60503
rect 27387 60469 27396 60503
rect 27344 60460 27396 60469
rect 29828 60503 29880 60512
rect 29828 60469 29837 60503
rect 29837 60469 29871 60503
rect 29871 60469 29880 60503
rect 29828 60460 29880 60469
rect 30564 60503 30616 60512
rect 30564 60469 30573 60503
rect 30573 60469 30607 60503
rect 30607 60469 30616 60503
rect 30564 60460 30616 60469
rect 34244 60503 34296 60512
rect 34244 60469 34253 60503
rect 34253 60469 34287 60503
rect 34287 60469 34296 60503
rect 34244 60460 34296 60469
rect 36452 60503 36504 60512
rect 36452 60469 36461 60503
rect 36461 60469 36495 60503
rect 36495 60469 36504 60503
rect 36452 60460 36504 60469
rect 41604 60503 41656 60512
rect 41604 60469 41613 60503
rect 41613 60469 41647 60503
rect 41647 60469 41656 60503
rect 41604 60460 41656 60469
rect 46756 60503 46808 60512
rect 46756 60469 46765 60503
rect 46765 60469 46799 60503
rect 46799 60469 46808 60503
rect 46756 60460 46808 60469
rect 49700 60503 49752 60512
rect 49700 60469 49709 60503
rect 49709 60469 49743 60503
rect 49743 60469 49752 60503
rect 49700 60460 49752 60469
rect 49792 60460 49844 60512
rect 53104 60503 53156 60512
rect 53104 60469 53113 60503
rect 53113 60469 53147 60503
rect 53147 60469 53156 60503
rect 53104 60460 53156 60469
rect 54852 60503 54904 60512
rect 54852 60469 54861 60503
rect 54861 60469 54895 60503
rect 54895 60469 54904 60503
rect 54852 60460 54904 60469
rect 55588 60503 55640 60512
rect 55588 60469 55597 60503
rect 55597 60469 55631 60503
rect 55631 60469 55640 60503
rect 55588 60460 55640 60469
rect 57060 60460 57112 60512
rect 58256 60503 58308 60512
rect 58256 60469 58265 60503
rect 58265 60469 58299 60503
rect 58299 60469 58308 60503
rect 58256 60460 58308 60469
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 12164 60256 12216 60308
rect 21824 60256 21876 60308
rect 28264 60256 28316 60308
rect 41604 60256 41656 60308
rect 49608 60256 49660 60308
rect 58256 60256 58308 60308
rect 54484 60188 54536 60240
rect 1584 60052 1636 60104
rect 2504 60095 2556 60104
rect 2504 60061 2513 60095
rect 2513 60061 2547 60095
rect 2547 60061 2556 60095
rect 2504 60052 2556 60061
rect 56232 60095 56284 60104
rect 56232 60061 56241 60095
rect 56241 60061 56275 60095
rect 56275 60061 56284 60095
rect 56232 60052 56284 60061
rect 2044 59984 2096 60036
rect 56048 59984 56100 60036
rect 57980 60027 58032 60036
rect 57980 59993 57989 60027
rect 57989 59993 58023 60027
rect 58023 59993 58032 60027
rect 57980 59984 58032 59993
rect 58992 59984 59044 60036
rect 2412 59916 2464 59968
rect 54760 59916 54812 59968
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 848 59644 900 59696
rect 1584 59619 1636 59628
rect 1584 59585 1593 59619
rect 1593 59585 1627 59619
rect 1627 59585 1636 59619
rect 1584 59576 1636 59585
rect 58716 59644 58768 59696
rect 57888 59576 57940 59628
rect 57244 59551 57296 59560
rect 57244 59517 57253 59551
rect 57253 59517 57287 59551
rect 57287 59517 57296 59551
rect 57244 59508 57296 59517
rect 2596 59483 2648 59492
rect 2596 59449 2605 59483
rect 2605 59449 2639 59483
rect 2639 59449 2648 59483
rect 2596 59440 2648 59449
rect 2688 59372 2740 59424
rect 31668 59372 31720 59424
rect 33692 59372 33744 59424
rect 59176 59372 59228 59424
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 1952 59032 2004 59084
rect 1584 59007 1636 59016
rect 1584 58973 1593 59007
rect 1593 58973 1627 59007
rect 1627 58973 1636 59007
rect 1584 58964 1636 58973
rect 40132 58964 40184 59016
rect 44088 59007 44140 59016
rect 44088 58973 44097 59007
rect 44097 58973 44131 59007
rect 44131 58973 44140 59007
rect 53104 59032 53156 59084
rect 44088 58964 44140 58973
rect 57336 58964 57388 59016
rect 56508 58896 56560 58948
rect 1768 58871 1820 58880
rect 1768 58837 1777 58871
rect 1777 58837 1811 58871
rect 1811 58837 1820 58871
rect 1768 58828 1820 58837
rect 44824 58828 44876 58880
rect 57336 58871 57388 58880
rect 57336 58837 57345 58871
rect 57345 58837 57379 58871
rect 57379 58837 57388 58871
rect 57336 58828 57388 58837
rect 58072 58871 58124 58880
rect 58072 58837 58081 58871
rect 58081 58837 58115 58871
rect 58115 58837 58124 58871
rect 58072 58828 58124 58837
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 1676 58531 1728 58540
rect 1676 58497 1685 58531
rect 1685 58497 1719 58531
rect 1719 58497 1728 58531
rect 1676 58488 1728 58497
rect 23112 58624 23164 58676
rect 15108 58599 15160 58608
rect 15108 58565 15117 58599
rect 15117 58565 15151 58599
rect 15151 58565 15160 58599
rect 15108 58556 15160 58565
rect 16672 58556 16724 58608
rect 17224 58599 17276 58608
rect 17224 58565 17233 58599
rect 17233 58565 17267 58599
rect 17267 58565 17276 58599
rect 58164 58624 58216 58676
rect 17224 58556 17276 58565
rect 16764 58488 16816 58540
rect 17408 58531 17460 58540
rect 17408 58497 17411 58531
rect 17411 58497 17460 58531
rect 16856 58420 16908 58472
rect 17408 58488 17460 58497
rect 21916 58488 21968 58540
rect 15384 58327 15436 58336
rect 15384 58293 15393 58327
rect 15393 58293 15427 58327
rect 15427 58293 15436 58327
rect 15384 58284 15436 58293
rect 16580 58352 16632 58404
rect 17224 58420 17276 58472
rect 39672 58531 39724 58540
rect 39672 58497 39681 58531
rect 39681 58497 39715 58531
rect 39715 58497 39724 58531
rect 39672 58488 39724 58497
rect 39764 58531 39816 58540
rect 39764 58497 39773 58531
rect 39773 58497 39807 58531
rect 39807 58497 39816 58531
rect 39764 58488 39816 58497
rect 43996 58488 44048 58540
rect 58164 58531 58216 58540
rect 58164 58497 58173 58531
rect 58173 58497 58207 58531
rect 58207 58497 58216 58531
rect 58164 58488 58216 58497
rect 57336 58420 57388 58472
rect 43904 58352 43956 58404
rect 17500 58327 17552 58336
rect 17500 58293 17509 58327
rect 17509 58293 17543 58327
rect 17543 58293 17552 58327
rect 17500 58284 17552 58293
rect 40040 58327 40092 58336
rect 40040 58293 40049 58327
rect 40049 58293 40083 58327
rect 40083 58293 40092 58327
rect 40040 58284 40092 58293
rect 55220 58284 55272 58336
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 16672 58080 16724 58132
rect 17132 58080 17184 58132
rect 1584 57919 1636 57928
rect 1584 57885 1593 57919
rect 1593 57885 1627 57919
rect 1627 57885 1636 57919
rect 1584 57876 1636 57885
rect 21272 57919 21324 57928
rect 21272 57885 21281 57919
rect 21281 57885 21315 57919
rect 21315 57885 21324 57919
rect 21272 57876 21324 57885
rect 21364 57919 21416 57928
rect 21364 57885 21373 57919
rect 21373 57885 21407 57919
rect 21407 57885 21416 57919
rect 21640 57919 21692 57928
rect 21364 57876 21416 57885
rect 21640 57885 21649 57919
rect 21649 57885 21683 57919
rect 21683 57885 21692 57919
rect 21640 57876 21692 57885
rect 22008 57876 22060 57928
rect 18144 57808 18196 57860
rect 1952 57740 2004 57792
rect 20904 57783 20956 57792
rect 20904 57749 20913 57783
rect 20913 57749 20947 57783
rect 20947 57749 20956 57783
rect 20904 57740 20956 57749
rect 21824 57808 21876 57860
rect 22468 57876 22520 57928
rect 23020 57919 23072 57928
rect 23020 57885 23029 57919
rect 23029 57885 23063 57919
rect 23063 57885 23072 57919
rect 23020 57876 23072 57885
rect 23204 57919 23256 57928
rect 23204 57885 23218 57919
rect 23218 57885 23252 57919
rect 23252 57885 23256 57919
rect 23204 57876 23256 57885
rect 23480 57876 23532 57928
rect 30748 57876 30800 57928
rect 31852 57919 31904 57928
rect 24768 57851 24820 57860
rect 23388 57783 23440 57792
rect 23388 57749 23397 57783
rect 23397 57749 23431 57783
rect 23431 57749 23440 57783
rect 23388 57740 23440 57749
rect 24768 57817 24777 57851
rect 24777 57817 24811 57851
rect 24811 57817 24820 57851
rect 24768 57808 24820 57817
rect 24860 57851 24912 57860
rect 24860 57817 24869 57851
rect 24869 57817 24903 57851
rect 24903 57817 24912 57851
rect 31852 57885 31861 57919
rect 31861 57885 31895 57919
rect 31895 57885 31904 57919
rect 31852 57876 31904 57885
rect 31944 57919 31996 57928
rect 31944 57885 31953 57919
rect 31953 57885 31987 57919
rect 31987 57885 31996 57919
rect 32220 57919 32272 57928
rect 31944 57876 31996 57885
rect 32220 57885 32229 57919
rect 32229 57885 32263 57919
rect 32263 57885 32272 57919
rect 32220 57876 32272 57885
rect 32496 57919 32548 57928
rect 32496 57885 32505 57919
rect 32505 57885 32539 57919
rect 32539 57885 32548 57919
rect 32496 57876 32548 57885
rect 32680 57919 32732 57928
rect 32680 57885 32689 57919
rect 32689 57885 32723 57919
rect 32723 57885 32732 57919
rect 32680 57876 32732 57885
rect 43904 57987 43956 57996
rect 37280 57876 37332 57928
rect 38660 57919 38712 57928
rect 38660 57885 38669 57919
rect 38669 57885 38703 57919
rect 38703 57885 38712 57919
rect 38660 57876 38712 57885
rect 38476 57851 38528 57860
rect 24860 57808 24912 57817
rect 25412 57740 25464 57792
rect 25504 57740 25556 57792
rect 31484 57783 31536 57792
rect 31484 57749 31493 57783
rect 31493 57749 31527 57783
rect 31527 57749 31536 57783
rect 31484 57740 31536 57749
rect 38476 57817 38485 57851
rect 38485 57817 38519 57851
rect 38519 57817 38528 57851
rect 38476 57808 38528 57817
rect 40224 57876 40276 57928
rect 43904 57953 43913 57987
rect 43913 57953 43947 57987
rect 43947 57953 43956 57987
rect 43904 57944 43956 57953
rect 43996 57944 44048 57996
rect 43812 57876 43864 57928
rect 44088 57919 44140 57928
rect 44088 57885 44097 57919
rect 44097 57885 44131 57919
rect 44131 57885 44140 57919
rect 44088 57876 44140 57885
rect 38936 57851 38988 57860
rect 38936 57817 38945 57851
rect 38945 57817 38979 57851
rect 38979 57817 38988 57851
rect 38936 57808 38988 57817
rect 39672 57808 39724 57860
rect 50068 57876 50120 57928
rect 49792 57808 49844 57860
rect 38844 57783 38896 57792
rect 38844 57749 38853 57783
rect 38853 57749 38887 57783
rect 38887 57749 38896 57783
rect 38844 57740 38896 57749
rect 44088 57740 44140 57792
rect 54576 57919 54628 57928
rect 54576 57885 54579 57919
rect 54579 57885 54628 57919
rect 54576 57876 54628 57885
rect 55220 57876 55272 57928
rect 54024 57808 54076 57860
rect 54760 57808 54812 57860
rect 58164 57851 58216 57860
rect 58164 57817 58173 57851
rect 58173 57817 58207 57851
rect 58207 57817 58216 57851
rect 58164 57808 58216 57817
rect 58256 57783 58308 57792
rect 58256 57749 58265 57783
rect 58265 57749 58299 57783
rect 58299 57749 58308 57783
rect 58256 57740 58308 57749
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 21640 57536 21692 57588
rect 20444 57511 20496 57520
rect 20444 57477 20453 57511
rect 20453 57477 20487 57511
rect 20487 57477 20496 57511
rect 20444 57468 20496 57477
rect 21364 57468 21416 57520
rect 25504 57536 25556 57588
rect 21824 57468 21876 57520
rect 23388 57468 23440 57520
rect 20168 57443 20220 57452
rect 20168 57409 20177 57443
rect 20177 57409 20211 57443
rect 20211 57409 20220 57443
rect 20168 57400 20220 57409
rect 20628 57400 20680 57452
rect 21272 57400 21324 57452
rect 22192 57400 22244 57452
rect 22468 57400 22520 57452
rect 34520 57536 34572 57588
rect 38660 57579 38712 57588
rect 32220 57468 32272 57520
rect 23204 57332 23256 57384
rect 29920 57400 29972 57452
rect 30748 57443 30800 57452
rect 30748 57409 30757 57443
rect 30757 57409 30791 57443
rect 30791 57409 30800 57443
rect 30748 57400 30800 57409
rect 31024 57443 31076 57452
rect 31024 57409 31033 57443
rect 31033 57409 31067 57443
rect 31067 57409 31076 57443
rect 31024 57400 31076 57409
rect 31116 57443 31168 57452
rect 31116 57409 31125 57443
rect 31125 57409 31159 57443
rect 31159 57409 31168 57443
rect 31392 57443 31444 57452
rect 31116 57400 31168 57409
rect 31392 57409 31401 57443
rect 31401 57409 31435 57443
rect 31435 57409 31444 57443
rect 31392 57400 31444 57409
rect 31576 57443 31628 57452
rect 31576 57409 31585 57443
rect 31585 57409 31619 57443
rect 31619 57409 31628 57443
rect 31576 57400 31628 57409
rect 37740 57468 37792 57520
rect 38660 57545 38669 57579
rect 38669 57545 38703 57579
rect 38703 57545 38712 57579
rect 38660 57536 38712 57545
rect 38844 57536 38896 57588
rect 49608 57536 49660 57588
rect 51080 57468 51132 57520
rect 25780 57332 25832 57384
rect 36084 57443 36136 57452
rect 36084 57409 36093 57443
rect 36093 57409 36127 57443
rect 36127 57409 36136 57443
rect 36360 57443 36412 57452
rect 36084 57400 36136 57409
rect 36360 57409 36369 57443
rect 36369 57409 36403 57443
rect 36403 57409 36412 57443
rect 36360 57400 36412 57409
rect 36636 57443 36688 57452
rect 36636 57409 36645 57443
rect 36645 57409 36679 57443
rect 36679 57409 36688 57443
rect 36636 57400 36688 57409
rect 38108 57443 38160 57452
rect 38108 57409 38117 57443
rect 38117 57409 38151 57443
rect 38151 57409 38160 57443
rect 38108 57400 38160 57409
rect 38200 57400 38252 57452
rect 38568 57400 38620 57452
rect 40132 57400 40184 57452
rect 54576 57536 54628 57588
rect 54024 57400 54076 57452
rect 54852 57443 54904 57452
rect 54852 57409 54861 57443
rect 54861 57409 54895 57443
rect 54895 57409 54904 57443
rect 54852 57400 54904 57409
rect 58164 57443 58216 57452
rect 58164 57409 58173 57443
rect 58173 57409 58207 57443
rect 58207 57409 58216 57443
rect 58164 57400 58216 57409
rect 53932 57375 53984 57384
rect 21548 57264 21600 57316
rect 20628 57196 20680 57248
rect 21916 57196 21968 57248
rect 23020 57196 23072 57248
rect 23112 57196 23164 57248
rect 25596 57196 25648 57248
rect 38016 57264 38068 57316
rect 53932 57341 53941 57375
rect 53941 57341 53975 57375
rect 53975 57341 53984 57375
rect 53932 57332 53984 57341
rect 40592 57264 40644 57316
rect 45376 57264 45428 57316
rect 51080 57264 51132 57316
rect 30380 57239 30432 57248
rect 30380 57205 30389 57239
rect 30389 57205 30423 57239
rect 30423 57205 30432 57239
rect 30380 57196 30432 57205
rect 31392 57196 31444 57248
rect 32496 57196 32548 57248
rect 35348 57239 35400 57248
rect 35348 57205 35357 57239
rect 35357 57205 35391 57239
rect 35391 57205 35400 57239
rect 35348 57196 35400 57205
rect 36360 57196 36412 57248
rect 54024 57196 54076 57248
rect 55588 57196 55640 57248
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 1768 56992 1820 57044
rect 31576 56992 31628 57044
rect 34520 56992 34572 57044
rect 34980 56992 35032 57044
rect 36084 56992 36136 57044
rect 36636 56992 36688 57044
rect 58256 56992 58308 57044
rect 22100 56924 22152 56976
rect 24860 56924 24912 56976
rect 40592 56924 40644 56976
rect 43812 56924 43864 56976
rect 2688 56856 2740 56908
rect 32680 56856 32732 56908
rect 1676 56831 1728 56840
rect 1676 56797 1685 56831
rect 1685 56797 1719 56831
rect 1719 56797 1728 56831
rect 1676 56788 1728 56797
rect 21640 56831 21692 56840
rect 21640 56797 21649 56831
rect 21649 56797 21683 56831
rect 21683 56797 21692 56831
rect 21640 56788 21692 56797
rect 21732 56831 21784 56840
rect 21732 56797 21742 56831
rect 21742 56797 21776 56831
rect 21776 56797 21784 56831
rect 21732 56788 21784 56797
rect 21916 56831 21968 56840
rect 21916 56797 21925 56831
rect 21925 56797 21959 56831
rect 21959 56797 21968 56831
rect 21916 56788 21968 56797
rect 22192 56788 22244 56840
rect 29920 56788 29972 56840
rect 38568 56788 38620 56840
rect 15752 56720 15804 56772
rect 17132 56720 17184 56772
rect 20628 56720 20680 56772
rect 21364 56720 21416 56772
rect 21824 56720 21876 56772
rect 41052 56788 41104 56840
rect 43996 56788 44048 56840
rect 44456 56831 44508 56840
rect 44456 56797 44465 56831
rect 44465 56797 44499 56831
rect 44499 56797 44508 56831
rect 44456 56788 44508 56797
rect 54024 56831 54076 56840
rect 54024 56797 54033 56831
rect 54033 56797 54067 56831
rect 54067 56797 54076 56831
rect 54024 56788 54076 56797
rect 54392 56831 54444 56840
rect 54392 56797 54401 56831
rect 54401 56797 54435 56831
rect 54435 56797 54444 56831
rect 54392 56788 54444 56797
rect 54576 56831 54628 56840
rect 54576 56797 54585 56831
rect 54585 56797 54619 56831
rect 54619 56797 54628 56831
rect 54576 56788 54628 56797
rect 58164 56763 58216 56772
rect 58164 56729 58173 56763
rect 58173 56729 58207 56763
rect 58207 56729 58216 56763
rect 58164 56720 58216 56729
rect 43996 56652 44048 56704
rect 53472 56695 53524 56704
rect 53472 56661 53481 56695
rect 53481 56661 53515 56695
rect 53515 56661 53524 56695
rect 53472 56652 53524 56661
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 8576 56448 8628 56500
rect 15660 56423 15712 56432
rect 15660 56389 15669 56423
rect 15669 56389 15703 56423
rect 15703 56389 15712 56423
rect 15660 56380 15712 56389
rect 29552 56448 29604 56500
rect 1676 56355 1728 56364
rect 1676 56321 1685 56355
rect 1685 56321 1719 56355
rect 1719 56321 1728 56355
rect 1676 56312 1728 56321
rect 9036 56312 9088 56364
rect 15568 56355 15620 56364
rect 15568 56321 15577 56355
rect 15577 56321 15611 56355
rect 15611 56321 15620 56355
rect 15568 56312 15620 56321
rect 15752 56355 15804 56364
rect 15752 56321 15761 56355
rect 15761 56321 15795 56355
rect 15795 56321 15804 56355
rect 15752 56312 15804 56321
rect 29460 56355 29512 56364
rect 29460 56321 29469 56355
rect 29469 56321 29503 56355
rect 29503 56321 29512 56355
rect 29460 56312 29512 56321
rect 29644 56355 29696 56364
rect 29644 56321 29653 56355
rect 29653 56321 29687 56355
rect 29687 56321 29696 56355
rect 29644 56312 29696 56321
rect 29920 56355 29972 56364
rect 29920 56321 29923 56355
rect 29923 56321 29972 56355
rect 20996 56244 21048 56296
rect 22008 56244 22060 56296
rect 29920 56312 29972 56321
rect 33600 56355 33652 56364
rect 33600 56321 33609 56355
rect 33609 56321 33643 56355
rect 33643 56321 33652 56355
rect 33600 56312 33652 56321
rect 33784 56423 33836 56432
rect 33784 56389 33793 56423
rect 33793 56389 33827 56423
rect 33827 56389 33836 56423
rect 33784 56380 33836 56389
rect 33968 56355 34020 56364
rect 33968 56321 33977 56355
rect 33977 56321 34011 56355
rect 34011 56321 34020 56355
rect 33968 56312 34020 56321
rect 48688 56448 48740 56500
rect 34980 56287 35032 56296
rect 29552 56176 29604 56228
rect 34980 56253 34989 56287
rect 34989 56253 35023 56287
rect 35023 56253 35032 56287
rect 34980 56244 35032 56253
rect 33968 56176 34020 56228
rect 1768 56151 1820 56160
rect 1768 56117 1777 56151
rect 1777 56117 1811 56151
rect 1811 56117 1820 56151
rect 1768 56108 1820 56117
rect 28356 56108 28408 56160
rect 29644 56108 29696 56160
rect 30472 56108 30524 56160
rect 35532 56108 35584 56160
rect 50068 56108 50120 56160
rect 58348 56151 58400 56160
rect 58348 56117 58357 56151
rect 58357 56117 58391 56151
rect 58391 56117 58400 56151
rect 58348 56108 58400 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 1768 55904 1820 55956
rect 29460 55904 29512 55956
rect 29644 55904 29696 55956
rect 31392 55904 31444 55956
rect 43996 55904 44048 55956
rect 44916 55904 44968 55956
rect 33600 55836 33652 55888
rect 39396 55836 39448 55888
rect 1676 55675 1728 55684
rect 1676 55641 1685 55675
rect 1685 55641 1719 55675
rect 1719 55641 1728 55675
rect 1676 55632 1728 55641
rect 43444 55564 43496 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 9128 55360 9180 55412
rect 43536 55360 43588 55412
rect 1584 55267 1636 55276
rect 1584 55233 1593 55267
rect 1593 55233 1627 55267
rect 1627 55233 1636 55267
rect 1584 55224 1636 55233
rect 43444 55267 43496 55276
rect 43444 55233 43453 55267
rect 43453 55233 43487 55267
rect 43487 55233 43496 55267
rect 43444 55224 43496 55233
rect 43812 55224 43864 55276
rect 47952 55224 48004 55276
rect 43904 55199 43956 55208
rect 43904 55165 43913 55199
rect 43913 55165 43947 55199
rect 43947 55165 43956 55199
rect 43904 55156 43956 55165
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 58348 54655 58400 54664
rect 58348 54621 58357 54655
rect 58357 54621 58391 54655
rect 58391 54621 58400 54655
rect 58348 54612 58400 54621
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 1676 54179 1728 54188
rect 1676 54145 1685 54179
rect 1685 54145 1719 54179
rect 1719 54145 1728 54179
rect 1676 54136 1728 54145
rect 43260 54179 43312 54188
rect 43260 54145 43269 54179
rect 43269 54145 43303 54179
rect 43303 54145 43312 54179
rect 43260 54136 43312 54145
rect 46940 54136 46992 54188
rect 42708 54111 42760 54120
rect 42708 54077 42717 54111
rect 42717 54077 42751 54111
rect 42751 54077 42760 54111
rect 42708 54068 42760 54077
rect 43904 54068 43956 54120
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 1584 53567 1636 53576
rect 1584 53533 1593 53567
rect 1593 53533 1627 53567
rect 1627 53533 1636 53567
rect 1584 53524 1636 53533
rect 18604 53388 18656 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 1952 53116 2004 53168
rect 19340 53116 19392 53168
rect 1584 53091 1636 53100
rect 1584 53057 1593 53091
rect 1593 53057 1627 53091
rect 1627 53057 1636 53091
rect 1584 53048 1636 53057
rect 1860 52844 1912 52896
rect 58348 52887 58400 52896
rect 58348 52853 58357 52887
rect 58357 52853 58391 52887
rect 58391 52853 58400 52887
rect 58348 52844 58400 52853
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 44088 52640 44140 52692
rect 46020 52640 46072 52692
rect 5448 52436 5500 52488
rect 1676 52411 1728 52420
rect 1676 52377 1685 52411
rect 1685 52377 1719 52411
rect 1719 52377 1728 52411
rect 1676 52368 1728 52377
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 5448 52071 5500 52080
rect 5448 52037 5457 52071
rect 5457 52037 5491 52071
rect 5491 52037 5500 52071
rect 5448 52028 5500 52037
rect 5172 52003 5224 52012
rect 5172 51969 5181 52003
rect 5181 51969 5215 52003
rect 5215 51969 5224 52003
rect 5172 51960 5224 51969
rect 4620 51892 4672 51944
rect 15568 51960 15620 52012
rect 20444 51960 20496 52012
rect 5724 51799 5776 51808
rect 5724 51765 5733 51799
rect 5733 51765 5767 51799
rect 5767 51765 5776 51799
rect 5724 51756 5776 51765
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 22192 51484 22244 51536
rect 1676 51323 1728 51332
rect 1676 51289 1685 51323
rect 1685 51289 1719 51323
rect 1719 51289 1728 51323
rect 1676 51280 1728 51289
rect 22192 51348 22244 51400
rect 22468 51391 22520 51400
rect 22468 51357 22477 51391
rect 22477 51357 22511 51391
rect 22511 51357 22520 51391
rect 22468 51348 22520 51357
rect 23020 51348 23072 51400
rect 58348 51391 58400 51400
rect 58348 51357 58357 51391
rect 58357 51357 58391 51391
rect 58391 51357 58400 51391
rect 58348 51348 58400 51357
rect 20444 51280 20496 51332
rect 43720 51280 43772 51332
rect 23112 51255 23164 51264
rect 23112 51221 23121 51255
rect 23121 51221 23155 51255
rect 23155 51221 23164 51255
rect 23112 51212 23164 51221
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 1676 50915 1728 50924
rect 1676 50881 1685 50915
rect 1685 50881 1719 50915
rect 1719 50881 1728 50915
rect 1676 50872 1728 50881
rect 8944 50736 8996 50788
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 57796 50260 57848 50312
rect 1676 50235 1728 50244
rect 1676 50201 1685 50235
rect 1685 50201 1719 50235
rect 1719 50201 1728 50235
rect 1676 50192 1728 50201
rect 20536 50124 20588 50176
rect 57888 50124 57940 50176
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 20444 49852 20496 49904
rect 20812 49895 20864 49904
rect 1676 49827 1728 49836
rect 1676 49793 1685 49827
rect 1685 49793 1719 49827
rect 1719 49793 1728 49827
rect 1676 49784 1728 49793
rect 20536 49827 20588 49836
rect 20536 49793 20545 49827
rect 20545 49793 20579 49827
rect 20579 49793 20588 49827
rect 20536 49784 20588 49793
rect 20812 49861 20821 49895
rect 20821 49861 20855 49895
rect 20855 49861 20864 49895
rect 20812 49852 20864 49861
rect 17868 49716 17920 49768
rect 20628 49716 20680 49768
rect 22008 49580 22060 49632
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 21640 49376 21692 49428
rect 17868 49172 17920 49224
rect 21548 49215 21600 49224
rect 21548 49181 21557 49215
rect 21557 49181 21591 49215
rect 21591 49181 21600 49215
rect 21548 49172 21600 49181
rect 20444 49104 20496 49156
rect 21456 49147 21508 49156
rect 21456 49113 21465 49147
rect 21465 49113 21499 49147
rect 21499 49113 21508 49147
rect 57980 49147 58032 49156
rect 21456 49104 21508 49113
rect 57980 49113 57989 49147
rect 57989 49113 58023 49147
rect 58023 49113 58032 49147
rect 57980 49104 58032 49113
rect 58900 49104 58952 49156
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 3332 48764 3384 48816
rect 20352 48764 20404 48816
rect 1676 48739 1728 48748
rect 1676 48705 1685 48739
rect 1685 48705 1719 48739
rect 1719 48705 1728 48739
rect 1676 48696 1728 48705
rect 20076 48739 20128 48748
rect 20076 48705 20085 48739
rect 20085 48705 20119 48739
rect 20119 48705 20128 48739
rect 20076 48696 20128 48705
rect 20628 48696 20680 48748
rect 22008 48739 22060 48748
rect 22008 48705 22017 48739
rect 22017 48705 22051 48739
rect 22051 48705 22060 48739
rect 22008 48696 22060 48705
rect 20444 48628 20496 48680
rect 20720 48628 20772 48680
rect 21548 48628 21600 48680
rect 19984 48560 20036 48612
rect 39304 48628 39356 48680
rect 24768 48560 24820 48612
rect 20260 48535 20312 48544
rect 20260 48501 20269 48535
rect 20269 48501 20303 48535
rect 20303 48501 20312 48535
rect 20260 48492 20312 48501
rect 22376 48492 22428 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 21732 48220 21784 48272
rect 22284 48220 22336 48272
rect 56876 48084 56928 48136
rect 1676 48059 1728 48068
rect 1676 48025 1685 48059
rect 1685 48025 1719 48059
rect 1719 48025 1728 48059
rect 1676 48016 1728 48025
rect 57336 48016 57388 48068
rect 57980 48059 58032 48068
rect 57980 48025 57989 48059
rect 57989 48025 58023 48059
rect 58023 48025 58032 48059
rect 57980 48016 58032 48025
rect 58348 48059 58400 48068
rect 58348 48025 58357 48059
rect 58357 48025 58391 48059
rect 58391 48025 58400 48059
rect 58348 48016 58400 48025
rect 16580 47948 16632 48000
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 1676 47651 1728 47660
rect 1676 47617 1685 47651
rect 1685 47617 1719 47651
rect 1719 47617 1728 47651
rect 1676 47608 1728 47617
rect 21456 47608 21508 47660
rect 41604 47608 41656 47660
rect 20352 47540 20404 47592
rect 57060 47540 57112 47592
rect 1492 47404 1544 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 17224 46996 17276 47048
rect 57612 46996 57664 47048
rect 1676 46971 1728 46980
rect 1676 46937 1685 46971
rect 1685 46937 1719 46971
rect 1719 46937 1728 46971
rect 1676 46928 1728 46937
rect 57888 46860 57940 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 21640 45976 21692 46028
rect 28356 45976 28408 46028
rect 1676 45883 1728 45892
rect 1676 45849 1685 45883
rect 1685 45849 1719 45883
rect 1719 45849 1728 45883
rect 1676 45840 1728 45849
rect 23204 45951 23256 45960
rect 23204 45917 23213 45951
rect 23213 45917 23247 45951
rect 23247 45917 23256 45951
rect 23204 45908 23256 45917
rect 56784 45840 56836 45892
rect 57980 45883 58032 45892
rect 57980 45849 57989 45883
rect 57989 45849 58023 45883
rect 58023 45849 58032 45883
rect 57980 45840 58032 45849
rect 58716 45840 58768 45892
rect 23296 45772 23348 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 21548 45568 21600 45620
rect 23204 45568 23256 45620
rect 1584 45475 1636 45484
rect 1584 45441 1593 45475
rect 1593 45441 1627 45475
rect 1627 45441 1636 45475
rect 1584 45432 1636 45441
rect 24124 45228 24176 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 9036 44956 9088 45008
rect 31484 44888 31536 44940
rect 45928 44888 45980 44940
rect 9128 44820 9180 44872
rect 19432 44820 19484 44872
rect 21272 44820 21324 44872
rect 54484 44820 54536 44872
rect 55956 44820 56008 44872
rect 1676 44795 1728 44804
rect 1676 44761 1685 44795
rect 1685 44761 1719 44795
rect 1719 44761 1728 44795
rect 1676 44752 1728 44761
rect 57244 44795 57296 44804
rect 57244 44761 57253 44795
rect 57253 44761 57287 44795
rect 57287 44761 57296 44795
rect 57244 44752 57296 44761
rect 57888 44752 57940 44804
rect 58440 44752 58492 44804
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 1676 44387 1728 44396
rect 1676 44353 1685 44387
rect 1685 44353 1719 44387
rect 1719 44353 1728 44387
rect 1676 44344 1728 44353
rect 15476 44140 15528 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 15476 43843 15528 43852
rect 15476 43809 15485 43843
rect 15485 43809 15519 43843
rect 15519 43809 15528 43843
rect 15476 43800 15528 43809
rect 16028 43775 16080 43784
rect 16028 43741 16037 43775
rect 16037 43741 16071 43775
rect 16071 43741 16080 43775
rect 16028 43732 16080 43741
rect 20076 43732 20128 43784
rect 47584 43732 47636 43784
rect 20444 43664 20496 43716
rect 20628 43664 20680 43716
rect 58164 43707 58216 43716
rect 58164 43673 58173 43707
rect 58173 43673 58207 43707
rect 58207 43673 58216 43707
rect 58164 43664 58216 43673
rect 15108 43639 15160 43648
rect 15108 43605 15117 43639
rect 15117 43605 15151 43639
rect 15151 43605 15160 43639
rect 15108 43596 15160 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 1584 43299 1636 43308
rect 1584 43265 1593 43299
rect 1593 43265 1627 43299
rect 1627 43265 1636 43299
rect 1584 43256 1636 43265
rect 4068 43052 4120 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 30564 42780 30616 42832
rect 32220 42780 32272 42832
rect 20076 42712 20128 42764
rect 22836 42712 22888 42764
rect 22744 42644 22796 42696
rect 31852 42644 31904 42696
rect 56968 42687 57020 42696
rect 56968 42653 56977 42687
rect 56977 42653 57011 42687
rect 57011 42653 57020 42687
rect 56968 42644 57020 42653
rect 57888 42687 57940 42696
rect 57888 42653 57897 42687
rect 57897 42653 57931 42687
rect 57931 42653 57940 42687
rect 57888 42644 57940 42653
rect 1676 42619 1728 42628
rect 1676 42585 1685 42619
rect 1685 42585 1719 42619
rect 1719 42585 1728 42619
rect 1676 42576 1728 42585
rect 5540 42576 5592 42628
rect 31760 42576 31812 42628
rect 58624 42576 58676 42628
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 3792 42304 3844 42356
rect 1676 42211 1728 42220
rect 1676 42177 1685 42211
rect 1685 42177 1719 42211
rect 1719 42177 1728 42211
rect 1676 42168 1728 42177
rect 4620 42211 4672 42220
rect 4620 42177 4629 42211
rect 4629 42177 4663 42211
rect 4663 42177 4672 42211
rect 4620 42168 4672 42177
rect 22652 42168 22704 42220
rect 23112 42211 23164 42220
rect 23112 42177 23121 42211
rect 23121 42177 23155 42211
rect 23155 42177 23164 42211
rect 23112 42168 23164 42177
rect 4896 42100 4948 42152
rect 27528 42100 27580 42152
rect 4068 42032 4120 42084
rect 32772 42032 32824 42084
rect 4988 42007 5040 42016
rect 4988 41973 4997 42007
rect 4997 41973 5031 42007
rect 5031 41973 5040 42007
rect 4988 41964 5040 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 22652 41803 22704 41812
rect 22652 41769 22661 41803
rect 22661 41769 22695 41803
rect 22695 41769 22704 41803
rect 22652 41760 22704 41769
rect 4988 41692 5040 41744
rect 22836 41599 22888 41608
rect 22836 41565 22845 41599
rect 22845 41565 22879 41599
rect 22879 41565 22888 41599
rect 22836 41556 22888 41565
rect 22928 41599 22980 41608
rect 22928 41565 22937 41599
rect 22937 41565 22971 41599
rect 22971 41565 22980 41599
rect 22928 41556 22980 41565
rect 24860 41556 24912 41608
rect 49148 41556 49200 41608
rect 1676 41531 1728 41540
rect 1676 41497 1685 41531
rect 1685 41497 1719 41531
rect 1719 41497 1728 41531
rect 1676 41488 1728 41497
rect 3976 41488 4028 41540
rect 57244 41531 57296 41540
rect 57244 41497 57253 41531
rect 57253 41497 57287 41531
rect 57287 41497 57296 41531
rect 57244 41488 57296 41497
rect 57888 41488 57940 41540
rect 58808 41488 58860 41540
rect 3884 41420 3936 41472
rect 4620 41420 4672 41472
rect 31852 41420 31904 41472
rect 32404 41420 32456 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 2964 41216 3016 41268
rect 3792 41216 3844 41268
rect 3976 41191 4028 41200
rect 3976 41157 3985 41191
rect 3985 41157 4019 41191
rect 4019 41157 4028 41191
rect 3976 41148 4028 41157
rect 1400 41080 1452 41132
rect 3884 41123 3936 41132
rect 3884 41089 3893 41123
rect 3893 41089 3927 41123
rect 3927 41089 3936 41123
rect 3884 41080 3936 41089
rect 4804 41012 4856 41064
rect 5540 41012 5592 41064
rect 18604 41012 18656 41064
rect 22560 41012 22612 41064
rect 11704 40876 11756 40928
rect 34428 40944 34480 40996
rect 22652 40876 22704 40928
rect 27620 40876 27672 40928
rect 34336 40876 34388 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 11704 40672 11756 40724
rect 18052 40672 18104 40724
rect 22652 40511 22704 40520
rect 22652 40477 22661 40511
rect 22661 40477 22695 40511
rect 22695 40477 22704 40511
rect 22652 40468 22704 40477
rect 23020 40511 23072 40520
rect 23020 40477 23029 40511
rect 23029 40477 23063 40511
rect 23063 40477 23072 40511
rect 23020 40468 23072 40477
rect 48228 40468 48280 40520
rect 1676 40443 1728 40452
rect 1676 40409 1685 40443
rect 1685 40409 1719 40443
rect 1719 40409 1728 40443
rect 1676 40400 1728 40409
rect 22836 40443 22888 40452
rect 22836 40409 22845 40443
rect 22845 40409 22879 40443
rect 22879 40409 22888 40443
rect 22836 40400 22888 40409
rect 28264 40400 28316 40452
rect 2780 40332 2832 40384
rect 23480 40332 23532 40384
rect 57888 40332 57940 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 1584 40060 1636 40112
rect 2412 40060 2464 40112
rect 3884 40128 3936 40180
rect 2780 40103 2832 40112
rect 2780 40069 2789 40103
rect 2789 40069 2823 40103
rect 2823 40069 2832 40103
rect 2780 40060 2832 40069
rect 58164 40103 58216 40112
rect 58164 40069 58173 40103
rect 58173 40069 58207 40103
rect 58207 40069 58216 40103
rect 58164 40060 58216 40069
rect 2688 40035 2740 40044
rect 2688 40001 2697 40035
rect 2697 40001 2731 40035
rect 2731 40001 2740 40035
rect 2964 40035 3016 40044
rect 2688 39992 2740 40001
rect 2964 40001 2967 40035
rect 2967 40001 3016 40035
rect 2964 39992 3016 40001
rect 3056 39831 3108 39840
rect 3056 39797 3065 39831
rect 3065 39797 3099 39831
rect 3099 39797 3108 39831
rect 3056 39788 3108 39797
rect 22652 39788 22704 39840
rect 56048 39788 56100 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 3056 39584 3108 39636
rect 22284 39584 22336 39636
rect 16580 39516 16632 39568
rect 21916 39516 21968 39568
rect 23020 39448 23072 39500
rect 23112 39423 23164 39432
rect 23112 39389 23121 39423
rect 23121 39389 23155 39423
rect 23155 39389 23164 39423
rect 23112 39380 23164 39389
rect 1400 39312 1452 39364
rect 2504 39312 2556 39364
rect 24860 39312 24912 39364
rect 42524 39312 42576 39364
rect 57060 39355 57112 39364
rect 57060 39321 57069 39355
rect 57069 39321 57103 39355
rect 57103 39321 57112 39355
rect 57060 39312 57112 39321
rect 57980 39355 58032 39364
rect 57980 39321 57989 39355
rect 57989 39321 58023 39355
rect 58023 39321 58032 39355
rect 57980 39312 58032 39321
rect 58532 39312 58584 39364
rect 29644 39244 29696 39296
rect 31760 39244 31812 39296
rect 37924 39244 37976 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 20536 39040 20588 39092
rect 22744 39040 22796 39092
rect 10324 38972 10376 39024
rect 26884 38972 26936 39024
rect 1676 38947 1728 38956
rect 1676 38913 1685 38947
rect 1685 38913 1719 38947
rect 1719 38913 1728 38947
rect 1676 38904 1728 38913
rect 20444 38947 20496 38956
rect 20444 38913 20453 38947
rect 20453 38913 20487 38947
rect 20487 38913 20496 38947
rect 20444 38904 20496 38913
rect 20720 38947 20772 38956
rect 20720 38913 20729 38947
rect 20729 38913 20763 38947
rect 20763 38913 20772 38947
rect 20720 38904 20772 38913
rect 20996 38904 21048 38956
rect 22652 38947 22704 38956
rect 22652 38913 22661 38947
rect 22661 38913 22695 38947
rect 22695 38913 22704 38947
rect 22652 38904 22704 38913
rect 22836 38947 22888 38956
rect 22836 38913 22845 38947
rect 22845 38913 22879 38947
rect 22879 38913 22888 38947
rect 22836 38904 22888 38913
rect 23020 38947 23072 38956
rect 23020 38913 23034 38947
rect 23034 38913 23068 38947
rect 23068 38913 23072 38947
rect 23020 38904 23072 38913
rect 26148 38836 26200 38888
rect 20720 38768 20772 38820
rect 24952 38768 25004 38820
rect 11704 38700 11756 38752
rect 21088 38743 21140 38752
rect 21088 38709 21097 38743
rect 21097 38709 21131 38743
rect 21131 38709 21140 38743
rect 21088 38700 21140 38709
rect 23848 38700 23900 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 2964 38428 3016 38480
rect 3700 38428 3752 38480
rect 21088 38428 21140 38480
rect 21640 38428 21692 38480
rect 2596 38360 2648 38412
rect 2504 38335 2556 38344
rect 2504 38301 2513 38335
rect 2513 38301 2547 38335
rect 2547 38301 2556 38335
rect 2504 38292 2556 38301
rect 2688 38292 2740 38344
rect 2872 38292 2924 38344
rect 18880 38360 18932 38412
rect 20628 38360 20680 38412
rect 21364 38335 21416 38344
rect 21364 38301 21373 38335
rect 21373 38301 21407 38335
rect 21407 38301 21416 38335
rect 21364 38292 21416 38301
rect 21456 38292 21508 38344
rect 21640 38335 21692 38344
rect 21640 38301 21649 38335
rect 21649 38301 21683 38335
rect 21683 38301 21692 38335
rect 21640 38292 21692 38301
rect 57888 38335 57940 38344
rect 13912 38224 13964 38276
rect 20996 38224 21048 38276
rect 14004 38156 14056 38208
rect 21824 38199 21876 38208
rect 21824 38165 21833 38199
rect 21833 38165 21867 38199
rect 21867 38165 21876 38199
rect 21824 38156 21876 38165
rect 57888 38301 57897 38335
rect 57897 38301 57931 38335
rect 57931 38301 57940 38335
rect 57888 38292 57940 38301
rect 57244 38267 57296 38276
rect 57244 38233 57253 38267
rect 57253 38233 57287 38267
rect 57287 38233 57296 38267
rect 57244 38224 57296 38233
rect 59084 38224 59136 38276
rect 58256 38156 58308 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 2688 37995 2740 38004
rect 2688 37961 2697 37995
rect 2697 37961 2731 37995
rect 2731 37961 2740 37995
rect 2688 37952 2740 37961
rect 1952 37884 2004 37936
rect 56324 37952 56376 38004
rect 11980 37927 12032 37936
rect 2320 37859 2372 37868
rect 2320 37825 2329 37859
rect 2329 37825 2363 37859
rect 2363 37825 2372 37859
rect 2320 37816 2372 37825
rect 2504 37859 2556 37868
rect 2504 37825 2513 37859
rect 2513 37825 2547 37859
rect 2547 37825 2556 37859
rect 2504 37816 2556 37825
rect 11980 37893 11989 37927
rect 11989 37893 12023 37927
rect 12023 37893 12032 37927
rect 11980 37884 12032 37893
rect 3700 37816 3752 37868
rect 11704 37859 11756 37868
rect 11704 37825 11713 37859
rect 11713 37825 11747 37859
rect 11747 37825 11756 37859
rect 11704 37816 11756 37825
rect 13912 37884 13964 37936
rect 14004 37884 14056 37936
rect 11336 37748 11388 37800
rect 17224 37816 17276 37868
rect 18880 37859 18932 37868
rect 18880 37825 18889 37859
rect 18889 37825 18923 37859
rect 18923 37825 18932 37859
rect 18880 37816 18932 37825
rect 18972 37859 19024 37868
rect 18972 37825 18981 37859
rect 18981 37825 19015 37859
rect 19015 37825 19024 37859
rect 18972 37816 19024 37825
rect 19708 37859 19760 37868
rect 19708 37825 19717 37859
rect 19717 37825 19751 37859
rect 19751 37825 19760 37859
rect 21456 37859 21508 37868
rect 19708 37816 19760 37825
rect 21456 37825 21465 37859
rect 21465 37825 21499 37859
rect 21499 37825 21508 37859
rect 21456 37816 21508 37825
rect 22192 37816 22244 37868
rect 22652 37816 22704 37868
rect 26148 37884 26200 37936
rect 41512 37884 41564 37936
rect 23204 37859 23256 37868
rect 20812 37748 20864 37800
rect 20904 37748 20956 37800
rect 23204 37825 23213 37859
rect 23213 37825 23247 37859
rect 23247 37825 23256 37859
rect 23204 37816 23256 37825
rect 18788 37680 18840 37732
rect 20444 37680 20496 37732
rect 17960 37612 18012 37664
rect 18880 37612 18932 37664
rect 19708 37612 19760 37664
rect 20352 37612 20404 37664
rect 26516 37748 26568 37800
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 20628 37408 20680 37460
rect 21364 37408 21416 37460
rect 23204 37408 23256 37460
rect 41696 37408 41748 37460
rect 48228 37408 48280 37460
rect 18972 37340 19024 37392
rect 46940 37340 46992 37392
rect 1584 37247 1636 37256
rect 1584 37213 1593 37247
rect 1593 37213 1627 37247
rect 1627 37213 1636 37247
rect 1584 37204 1636 37213
rect 19708 37247 19760 37256
rect 19708 37213 19717 37247
rect 19717 37213 19751 37247
rect 19751 37213 19760 37247
rect 19708 37204 19760 37213
rect 20536 37247 20588 37256
rect 20536 37213 20545 37247
rect 20545 37213 20579 37247
rect 20579 37213 20588 37247
rect 20536 37204 20588 37213
rect 20812 37272 20864 37324
rect 21548 37204 21600 37256
rect 21916 37247 21968 37256
rect 21916 37213 21925 37247
rect 21925 37213 21959 37247
rect 21959 37213 21968 37247
rect 21916 37204 21968 37213
rect 23020 37204 23072 37256
rect 24124 37204 24176 37256
rect 25596 37204 25648 37256
rect 36452 37204 36504 37256
rect 45192 37247 45244 37256
rect 45192 37213 45201 37247
rect 45201 37213 45235 37247
rect 45235 37213 45244 37247
rect 45192 37204 45244 37213
rect 45376 37272 45428 37324
rect 2412 37179 2464 37188
rect 2412 37145 2421 37179
rect 2421 37145 2455 37179
rect 2455 37145 2464 37179
rect 2412 37136 2464 37145
rect 11336 37136 11388 37188
rect 2136 37068 2188 37120
rect 20720 37068 20772 37120
rect 21364 37136 21416 37188
rect 22192 37179 22244 37188
rect 22192 37145 22201 37179
rect 22201 37145 22235 37179
rect 22235 37145 22244 37179
rect 22192 37136 22244 37145
rect 44088 37136 44140 37188
rect 22836 37068 22888 37120
rect 43904 37068 43956 37120
rect 45652 37068 45704 37120
rect 57704 37204 57756 37256
rect 46296 37179 46348 37188
rect 46296 37145 46305 37179
rect 46305 37145 46339 37179
rect 46339 37145 46348 37179
rect 46296 37136 46348 37145
rect 58164 37179 58216 37188
rect 58164 37145 58173 37179
rect 58173 37145 58207 37179
rect 58207 37145 58216 37179
rect 58164 37136 58216 37145
rect 59176 37068 59228 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 18420 36864 18472 36916
rect 20536 36864 20588 36916
rect 1768 36796 1820 36848
rect 1400 36728 1452 36780
rect 21088 36839 21140 36848
rect 20720 36771 20772 36780
rect 20720 36737 20729 36771
rect 20729 36737 20763 36771
rect 20763 36737 20772 36771
rect 20720 36728 20772 36737
rect 21088 36805 21097 36839
rect 21097 36805 21131 36839
rect 21131 36805 21140 36839
rect 21088 36796 21140 36805
rect 21640 36864 21692 36916
rect 26884 36864 26936 36916
rect 38936 36864 38988 36916
rect 45376 36864 45428 36916
rect 22192 36796 22244 36848
rect 20996 36771 21048 36780
rect 20996 36737 21005 36771
rect 21005 36737 21039 36771
rect 21039 36737 21048 36771
rect 20996 36728 21048 36737
rect 21180 36771 21232 36780
rect 21180 36737 21194 36771
rect 21194 36737 21228 36771
rect 21228 36737 21232 36771
rect 21180 36728 21232 36737
rect 23020 36728 23072 36780
rect 23388 36771 23440 36780
rect 23388 36737 23397 36771
rect 23397 36737 23431 36771
rect 23431 36737 23440 36771
rect 23388 36728 23440 36737
rect 23480 36771 23532 36780
rect 23480 36737 23489 36771
rect 23489 36737 23523 36771
rect 23523 36737 23532 36771
rect 23480 36728 23532 36737
rect 43168 36728 43220 36780
rect 45652 36839 45704 36848
rect 45652 36805 45661 36839
rect 45661 36805 45695 36839
rect 45695 36805 45704 36839
rect 45652 36796 45704 36805
rect 48688 36728 48740 36780
rect 12348 36524 12400 36576
rect 36544 36660 36596 36712
rect 16764 36592 16816 36644
rect 21088 36592 21140 36644
rect 26884 36592 26936 36644
rect 58992 36592 59044 36644
rect 21640 36524 21692 36576
rect 22652 36524 22704 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 1768 36363 1820 36372
rect 1768 36329 1777 36363
rect 1777 36329 1811 36363
rect 1811 36329 1820 36363
rect 1768 36320 1820 36329
rect 1860 36252 1912 36304
rect 2320 36184 2372 36236
rect 2596 36184 2648 36236
rect 27344 36320 27396 36372
rect 46296 36320 46348 36372
rect 25136 36295 25188 36304
rect 25136 36261 25145 36295
rect 25145 36261 25179 36295
rect 25179 36261 25188 36295
rect 25136 36252 25188 36261
rect 32956 36252 33008 36304
rect 1676 36091 1728 36100
rect 1676 36057 1685 36091
rect 1685 36057 1719 36091
rect 1719 36057 1728 36091
rect 1676 36048 1728 36057
rect 18604 36159 18656 36168
rect 18604 36125 18613 36159
rect 18613 36125 18647 36159
rect 18647 36125 18656 36159
rect 18604 36116 18656 36125
rect 21272 36116 21324 36168
rect 21640 36159 21692 36168
rect 21640 36125 21649 36159
rect 21649 36125 21683 36159
rect 21683 36125 21692 36159
rect 21640 36116 21692 36125
rect 22376 36159 22428 36168
rect 20996 36048 21048 36100
rect 21456 36048 21508 36100
rect 22376 36125 22385 36159
rect 22385 36125 22419 36159
rect 22419 36125 22428 36159
rect 22376 36116 22428 36125
rect 22652 36159 22704 36168
rect 22652 36125 22661 36159
rect 22661 36125 22695 36159
rect 22695 36125 22704 36159
rect 22652 36116 22704 36125
rect 24952 36159 25004 36168
rect 24952 36125 24961 36159
rect 24961 36125 24995 36159
rect 24995 36125 25004 36159
rect 24952 36116 25004 36125
rect 20444 35980 20496 36032
rect 21272 35980 21324 36032
rect 24768 36091 24820 36100
rect 24768 36057 24777 36091
rect 24777 36057 24811 36091
rect 24811 36057 24820 36091
rect 24768 36048 24820 36057
rect 40868 36048 40920 36100
rect 57980 36091 58032 36100
rect 57980 36057 57989 36091
rect 57989 36057 58023 36091
rect 58023 36057 58032 36091
rect 57980 36048 58032 36057
rect 59176 36048 59228 36100
rect 26424 35980 26476 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 2228 35776 2280 35828
rect 17960 35776 18012 35828
rect 1860 35708 1912 35760
rect 20628 35776 20680 35828
rect 22192 35776 22244 35828
rect 35440 35776 35492 35828
rect 38936 35776 38988 35828
rect 2044 35683 2096 35692
rect 2044 35649 2053 35683
rect 2053 35649 2087 35683
rect 2087 35649 2096 35683
rect 2044 35640 2096 35649
rect 2412 35683 2464 35692
rect 2412 35649 2426 35683
rect 2426 35649 2460 35683
rect 2460 35649 2464 35683
rect 2412 35640 2464 35649
rect 2688 35572 2740 35624
rect 20076 35708 20128 35760
rect 20996 35708 21048 35760
rect 18512 35683 18564 35692
rect 18512 35649 18521 35683
rect 18521 35649 18555 35683
rect 18555 35649 18564 35683
rect 18512 35640 18564 35649
rect 18604 35572 18656 35624
rect 4712 35436 4764 35488
rect 18788 35683 18840 35692
rect 18788 35649 18797 35683
rect 18797 35649 18831 35683
rect 18831 35649 18840 35683
rect 20812 35683 20864 35692
rect 18788 35640 18840 35649
rect 20812 35649 20821 35683
rect 20821 35649 20855 35683
rect 20855 35649 20864 35683
rect 20812 35640 20864 35649
rect 20996 35572 21048 35624
rect 21272 35683 21324 35692
rect 21272 35649 21286 35683
rect 21286 35649 21320 35683
rect 21320 35649 21324 35683
rect 21272 35640 21324 35649
rect 36360 35708 36412 35760
rect 22008 35683 22060 35692
rect 22008 35649 22017 35683
rect 22017 35649 22051 35683
rect 22051 35649 22060 35683
rect 22008 35640 22060 35649
rect 24860 35640 24912 35692
rect 25136 35640 25188 35692
rect 25320 35683 25372 35692
rect 25320 35649 25329 35683
rect 25329 35649 25363 35683
rect 25363 35649 25372 35683
rect 25320 35640 25372 35649
rect 21456 35572 21508 35624
rect 24032 35572 24084 35624
rect 25412 35615 25464 35624
rect 25412 35581 25421 35615
rect 25421 35581 25455 35615
rect 25455 35581 25464 35615
rect 25412 35572 25464 35581
rect 26884 35504 26936 35556
rect 23572 35436 23624 35488
rect 24308 35436 24360 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4712 35232 4764 35284
rect 16396 35096 16448 35148
rect 1492 35028 1544 35080
rect 2228 35071 2280 35080
rect 2228 35037 2237 35071
rect 2237 35037 2271 35071
rect 2271 35037 2280 35071
rect 2228 35028 2280 35037
rect 2412 35071 2464 35080
rect 2412 35037 2426 35071
rect 2426 35037 2460 35071
rect 2460 35037 2464 35071
rect 16212 35071 16264 35080
rect 2412 35028 2464 35037
rect 16212 35037 16221 35071
rect 16221 35037 16255 35071
rect 16255 35037 16264 35071
rect 16212 35028 16264 35037
rect 16304 35071 16356 35080
rect 16304 35037 16313 35071
rect 16313 35037 16347 35071
rect 16347 35037 16356 35071
rect 21548 35096 21600 35148
rect 22192 35232 22244 35284
rect 22376 35275 22428 35284
rect 22376 35241 22385 35275
rect 22385 35241 22419 35275
rect 22419 35241 22428 35275
rect 24860 35275 24912 35284
rect 22376 35232 22428 35241
rect 24860 35241 24869 35275
rect 24869 35241 24903 35275
rect 24903 35241 24912 35275
rect 24860 35232 24912 35241
rect 24952 35164 25004 35216
rect 22468 35139 22520 35148
rect 16304 35028 16356 35037
rect 2320 35003 2372 35012
rect 2320 34969 2329 35003
rect 2329 34969 2363 35003
rect 2363 34969 2372 35003
rect 2320 34960 2372 34969
rect 15384 34960 15436 35012
rect 15844 34935 15896 34944
rect 15844 34901 15853 34935
rect 15853 34901 15887 34935
rect 15887 34901 15896 34935
rect 15844 34892 15896 34901
rect 22100 35071 22152 35080
rect 22100 35037 22109 35071
rect 22109 35037 22143 35071
rect 22143 35037 22152 35071
rect 22468 35105 22477 35139
rect 22477 35105 22511 35139
rect 22511 35105 22520 35139
rect 22468 35096 22520 35105
rect 22100 35028 22152 35037
rect 18696 34960 18748 35012
rect 24768 35096 24820 35148
rect 24032 35071 24084 35080
rect 24032 35037 24041 35071
rect 24041 35037 24075 35071
rect 24075 35037 24084 35071
rect 24032 35028 24084 35037
rect 24860 35028 24912 35080
rect 25228 35232 25280 35284
rect 25504 35096 25556 35148
rect 36544 35164 36596 35216
rect 49884 35164 49936 35216
rect 21180 34935 21232 34944
rect 21180 34901 21189 34935
rect 21189 34901 21223 34935
rect 21223 34901 21232 34935
rect 21180 34892 21232 34901
rect 22744 34935 22796 34944
rect 22744 34901 22753 34935
rect 22753 34901 22787 34935
rect 22787 34901 22796 34935
rect 22744 34892 22796 34901
rect 24124 34960 24176 35012
rect 24216 34960 24268 35012
rect 47676 35028 47728 35080
rect 51724 35028 51776 35080
rect 25504 34960 25556 35012
rect 58072 35028 58124 35080
rect 58164 35003 58216 35012
rect 58164 34969 58173 35003
rect 58173 34969 58207 35003
rect 58207 34969 58216 35003
rect 58164 34960 58216 34969
rect 24768 34892 24820 34944
rect 57152 34892 57204 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 15844 34688 15896 34740
rect 27620 34688 27672 34740
rect 20996 34620 21048 34672
rect 1676 34595 1728 34604
rect 1676 34561 1685 34595
rect 1685 34561 1719 34595
rect 1719 34561 1728 34595
rect 1676 34552 1728 34561
rect 16212 34552 16264 34604
rect 17960 34552 18012 34604
rect 21272 34620 21324 34672
rect 21180 34552 21232 34604
rect 24768 34620 24820 34672
rect 24860 34620 24912 34672
rect 35440 34620 35492 34672
rect 18696 34484 18748 34536
rect 21916 34484 21968 34536
rect 23112 34484 23164 34536
rect 23388 34552 23440 34604
rect 23664 34595 23716 34604
rect 23664 34561 23673 34595
rect 23673 34561 23707 34595
rect 23707 34561 23716 34595
rect 23664 34552 23716 34561
rect 23848 34595 23900 34604
rect 23848 34561 23857 34595
rect 23857 34561 23891 34595
rect 23891 34561 23900 34595
rect 23848 34552 23900 34561
rect 24952 34595 25004 34604
rect 20076 34416 20128 34468
rect 23664 34416 23716 34468
rect 24216 34416 24268 34468
rect 24492 34484 24544 34536
rect 24952 34561 24961 34595
rect 24961 34561 24995 34595
rect 24995 34561 25004 34595
rect 24952 34552 25004 34561
rect 25688 34484 25740 34536
rect 26884 34484 26936 34536
rect 56416 34484 56468 34536
rect 25412 34416 25464 34468
rect 32956 34348 33008 34400
rect 34612 34348 34664 34400
rect 43260 34348 43312 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 20260 34144 20312 34196
rect 21180 34144 21232 34196
rect 21640 34144 21692 34196
rect 1860 34119 1912 34128
rect 1860 34085 1869 34119
rect 1869 34085 1903 34119
rect 1903 34085 1912 34119
rect 1860 34076 1912 34085
rect 5724 34076 5776 34128
rect 22468 34144 22520 34196
rect 12348 34008 12400 34060
rect 17776 34008 17828 34060
rect 21640 34008 21692 34060
rect 17224 33983 17276 33992
rect 17224 33949 17233 33983
rect 17233 33949 17267 33983
rect 17267 33949 17276 33983
rect 17224 33940 17276 33949
rect 17868 33940 17920 33992
rect 19340 33940 19392 33992
rect 20260 33940 20312 33992
rect 1676 33915 1728 33924
rect 1676 33881 1685 33915
rect 1685 33881 1719 33915
rect 1719 33881 1728 33915
rect 1676 33872 1728 33881
rect 17316 33915 17368 33924
rect 17316 33881 17325 33915
rect 17325 33881 17359 33915
rect 17359 33881 17368 33915
rect 17316 33872 17368 33881
rect 17960 33872 18012 33924
rect 18972 33804 19024 33856
rect 19340 33804 19392 33856
rect 20076 33847 20128 33856
rect 20076 33813 20085 33847
rect 20085 33813 20119 33847
rect 20119 33813 20128 33847
rect 20076 33804 20128 33813
rect 20352 33847 20404 33856
rect 20352 33813 20361 33847
rect 20361 33813 20395 33847
rect 20395 33813 20404 33847
rect 22928 33940 22980 33992
rect 25044 34076 25096 34128
rect 25780 34076 25832 34128
rect 24768 34008 24820 34060
rect 22836 33872 22888 33924
rect 24676 33983 24728 33992
rect 24676 33949 24686 33983
rect 24686 33949 24720 33983
rect 24720 33949 24728 33983
rect 24676 33940 24728 33949
rect 24860 33983 24912 33992
rect 24860 33949 24869 33983
rect 24869 33949 24903 33983
rect 24903 33949 24912 33983
rect 24860 33940 24912 33949
rect 25412 33940 25464 33992
rect 26056 33940 26108 33992
rect 20352 33804 20404 33813
rect 23940 33804 23992 33856
rect 25228 33847 25280 33856
rect 25228 33813 25237 33847
rect 25237 33813 25271 33847
rect 25271 33813 25280 33847
rect 25228 33804 25280 33813
rect 40040 33940 40092 33992
rect 40592 33983 40644 33992
rect 40592 33949 40606 33983
rect 40606 33949 40640 33983
rect 40640 33949 40644 33983
rect 40592 33940 40644 33949
rect 40500 33915 40552 33924
rect 40500 33881 40509 33915
rect 40509 33881 40543 33915
rect 40543 33881 40552 33915
rect 40500 33872 40552 33881
rect 57980 33983 58032 33992
rect 57980 33949 57989 33983
rect 57989 33949 58023 33983
rect 58023 33949 58032 33983
rect 57980 33940 58032 33949
rect 50988 33872 51040 33924
rect 58992 33872 59044 33924
rect 44088 33804 44140 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 19064 33600 19116 33652
rect 20536 33600 20588 33652
rect 1952 33532 2004 33584
rect 20076 33532 20128 33584
rect 32864 33600 32916 33652
rect 21180 33532 21232 33584
rect 25320 33575 25372 33584
rect 1676 33507 1728 33516
rect 1676 33473 1685 33507
rect 1685 33473 1719 33507
rect 1719 33473 1728 33507
rect 1676 33464 1728 33473
rect 18880 33464 18932 33516
rect 19432 33464 19484 33516
rect 20260 33464 20312 33516
rect 23572 33507 23624 33516
rect 23572 33473 23581 33507
rect 23581 33473 23615 33507
rect 23615 33473 23624 33507
rect 23572 33464 23624 33473
rect 25320 33541 25329 33575
rect 25329 33541 25363 33575
rect 25363 33541 25372 33575
rect 35348 33600 35400 33652
rect 25320 33532 25372 33541
rect 17960 33439 18012 33448
rect 17960 33405 17969 33439
rect 17969 33405 18003 33439
rect 18003 33405 18012 33439
rect 17960 33396 18012 33405
rect 23664 33396 23716 33448
rect 23940 33439 23992 33448
rect 23940 33405 23949 33439
rect 23949 33405 23983 33439
rect 23983 33405 23992 33439
rect 23940 33396 23992 33405
rect 25412 33507 25464 33516
rect 25412 33473 25421 33507
rect 25421 33473 25455 33507
rect 25455 33473 25464 33507
rect 25412 33464 25464 33473
rect 25780 33464 25832 33516
rect 27344 33507 27396 33516
rect 27344 33473 27353 33507
rect 27353 33473 27387 33507
rect 27387 33473 27396 33507
rect 27344 33464 27396 33473
rect 27528 33507 27580 33516
rect 27528 33473 27537 33507
rect 27537 33473 27571 33507
rect 27571 33473 27580 33507
rect 27528 33464 27580 33473
rect 27620 33464 27672 33516
rect 28448 33507 28500 33516
rect 28448 33473 28457 33507
rect 28457 33473 28491 33507
rect 28491 33473 28500 33507
rect 28448 33464 28500 33473
rect 32128 33464 32180 33516
rect 32772 33507 32824 33516
rect 32772 33473 32781 33507
rect 32781 33473 32815 33507
rect 32815 33473 32824 33507
rect 32772 33464 32824 33473
rect 32956 33507 33008 33516
rect 32956 33473 32965 33507
rect 32965 33473 32999 33507
rect 32999 33473 33008 33507
rect 32956 33464 33008 33473
rect 33048 33507 33100 33516
rect 33048 33473 33065 33507
rect 33065 33473 33099 33507
rect 33099 33473 33100 33507
rect 33048 33464 33100 33473
rect 34060 33464 34112 33516
rect 36084 33464 36136 33516
rect 40592 33464 40644 33516
rect 26608 33396 26660 33448
rect 32772 33328 32824 33380
rect 32864 33328 32916 33380
rect 34704 33328 34756 33380
rect 17316 33260 17368 33312
rect 17960 33260 18012 33312
rect 19432 33260 19484 33312
rect 20352 33260 20404 33312
rect 25688 33303 25740 33312
rect 25688 33269 25697 33303
rect 25697 33269 25731 33303
rect 25731 33269 25740 33303
rect 25688 33260 25740 33269
rect 29552 33260 29604 33312
rect 33416 33260 33468 33312
rect 46940 33260 46992 33312
rect 48964 33260 49016 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 17224 33056 17276 33108
rect 17316 33056 17368 33108
rect 19616 32988 19668 33040
rect 14464 32920 14516 32972
rect 17224 32920 17276 32972
rect 18972 32920 19024 32972
rect 8944 32852 8996 32904
rect 17868 32895 17920 32904
rect 17868 32861 17877 32895
rect 17877 32861 17911 32895
rect 17911 32861 17920 32895
rect 17868 32852 17920 32861
rect 17960 32895 18012 32904
rect 17960 32861 17969 32895
rect 17969 32861 18003 32895
rect 18003 32861 18012 32895
rect 17960 32852 18012 32861
rect 18328 32852 18380 32904
rect 18788 32852 18840 32904
rect 19340 32852 19392 32904
rect 19524 32784 19576 32836
rect 17224 32716 17276 32768
rect 18052 32716 18104 32768
rect 19340 32716 19392 32768
rect 19432 32716 19484 32768
rect 20076 32852 20128 32904
rect 20260 32895 20312 32904
rect 20260 32861 20269 32895
rect 20269 32861 20303 32895
rect 20303 32861 20312 32895
rect 20812 32920 20864 32972
rect 33508 33056 33560 33108
rect 34060 33099 34112 33108
rect 34060 33065 34069 33099
rect 34069 33065 34103 33099
rect 34103 33065 34112 33099
rect 34060 33056 34112 33065
rect 27528 32988 27580 33040
rect 32772 32988 32824 33040
rect 43996 32988 44048 33040
rect 58164 32963 58216 32972
rect 20260 32852 20312 32861
rect 19892 32784 19944 32836
rect 21180 32895 21232 32904
rect 21180 32861 21189 32895
rect 21189 32861 21223 32895
rect 21223 32861 21232 32895
rect 21180 32852 21232 32861
rect 21548 32895 21600 32904
rect 21548 32861 21557 32895
rect 21557 32861 21591 32895
rect 21591 32861 21600 32895
rect 21548 32852 21600 32861
rect 21732 32895 21784 32904
rect 21732 32861 21741 32895
rect 21741 32861 21775 32895
rect 21775 32861 21784 32895
rect 21732 32852 21784 32861
rect 21916 32895 21968 32904
rect 21916 32861 21925 32895
rect 21925 32861 21959 32895
rect 21959 32861 21968 32895
rect 21916 32852 21968 32861
rect 23572 32852 23624 32904
rect 25504 32895 25556 32904
rect 25504 32861 25513 32895
rect 25513 32861 25547 32895
rect 25547 32861 25556 32895
rect 25504 32852 25556 32861
rect 25596 32895 25648 32904
rect 25596 32861 25606 32895
rect 25606 32861 25640 32895
rect 25640 32861 25648 32895
rect 25596 32852 25648 32861
rect 25964 32895 26016 32904
rect 25964 32861 25978 32895
rect 25978 32861 26012 32895
rect 26012 32861 26016 32895
rect 25964 32852 26016 32861
rect 26148 32852 26200 32904
rect 20812 32784 20864 32836
rect 21364 32784 21416 32836
rect 27344 32852 27396 32904
rect 27528 32852 27580 32904
rect 33048 32895 33100 32904
rect 33048 32861 33057 32895
rect 33057 32861 33091 32895
rect 33091 32861 33100 32895
rect 33048 32852 33100 32861
rect 58164 32929 58173 32963
rect 58173 32929 58207 32963
rect 58207 32929 58216 32963
rect 58164 32920 58216 32929
rect 27620 32784 27672 32836
rect 33416 32895 33468 32904
rect 33416 32861 33425 32895
rect 33425 32861 33459 32895
rect 33459 32861 33468 32895
rect 42892 32895 42944 32904
rect 33416 32852 33468 32861
rect 42892 32861 42901 32895
rect 42901 32861 42935 32895
rect 42935 32861 42944 32895
rect 42892 32852 42944 32861
rect 43076 32895 43128 32904
rect 43076 32861 43083 32895
rect 43083 32861 43128 32895
rect 43076 32852 43128 32861
rect 43352 32895 43404 32904
rect 43352 32861 43366 32895
rect 43366 32861 43400 32895
rect 43400 32861 43404 32895
rect 43352 32852 43404 32861
rect 57520 32852 57572 32904
rect 33968 32827 34020 32836
rect 25504 32716 25556 32768
rect 33968 32793 33977 32827
rect 33977 32793 34011 32827
rect 34011 32793 34020 32827
rect 33968 32784 34020 32793
rect 35348 32784 35400 32836
rect 44272 32784 44324 32836
rect 57060 32827 57112 32836
rect 57060 32793 57069 32827
rect 57069 32793 57103 32827
rect 57103 32793 57112 32827
rect 57060 32784 57112 32793
rect 33784 32716 33836 32768
rect 36544 32716 36596 32768
rect 48044 32716 48096 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 17960 32512 18012 32564
rect 18788 32512 18840 32564
rect 19340 32512 19392 32564
rect 19984 32512 20036 32564
rect 2320 32444 2372 32496
rect 17868 32444 17920 32496
rect 19432 32444 19484 32496
rect 1676 32419 1728 32428
rect 1676 32385 1685 32419
rect 1685 32385 1719 32419
rect 1719 32385 1728 32419
rect 1676 32376 1728 32385
rect 17408 32376 17460 32428
rect 18236 32308 18288 32360
rect 18420 32308 18472 32360
rect 18788 32419 18840 32428
rect 18788 32385 18797 32419
rect 18797 32385 18831 32419
rect 18831 32385 18840 32419
rect 20628 32444 20680 32496
rect 25228 32444 25280 32496
rect 27344 32444 27396 32496
rect 18788 32376 18840 32385
rect 19984 32376 20036 32428
rect 20260 32419 20312 32428
rect 20260 32385 20269 32419
rect 20269 32385 20303 32419
rect 20303 32385 20312 32419
rect 20260 32376 20312 32385
rect 22192 32419 22244 32428
rect 19248 32351 19300 32360
rect 19248 32317 19257 32351
rect 19257 32317 19291 32351
rect 19291 32317 19300 32351
rect 19248 32308 19300 32317
rect 19892 32351 19944 32360
rect 19892 32317 19901 32351
rect 19901 32317 19935 32351
rect 19935 32317 19944 32351
rect 19892 32308 19944 32317
rect 19432 32240 19484 32292
rect 22192 32385 22201 32419
rect 22201 32385 22235 32419
rect 22235 32385 22244 32419
rect 22192 32376 22244 32385
rect 22560 32419 22612 32428
rect 19064 32172 19116 32224
rect 20536 32240 20588 32292
rect 22560 32385 22569 32419
rect 22569 32385 22603 32419
rect 22603 32385 22612 32419
rect 22560 32376 22612 32385
rect 36544 32512 36596 32564
rect 42800 32512 42852 32564
rect 44088 32444 44140 32496
rect 46112 32444 46164 32496
rect 33508 32419 33560 32428
rect 33508 32385 33517 32419
rect 33517 32385 33551 32419
rect 33551 32385 33560 32419
rect 33508 32376 33560 32385
rect 33876 32376 33928 32428
rect 44732 32419 44784 32428
rect 23020 32240 23072 32292
rect 25964 32240 26016 32292
rect 27160 32240 27212 32292
rect 27528 32240 27580 32292
rect 24768 32172 24820 32224
rect 34152 32308 34204 32360
rect 44732 32385 44741 32419
rect 44741 32385 44775 32419
rect 44775 32385 44784 32419
rect 44732 32376 44784 32385
rect 43352 32308 43404 32360
rect 44456 32308 44508 32360
rect 45744 32308 45796 32360
rect 33508 32240 33560 32292
rect 37004 32240 37056 32292
rect 42616 32240 42668 32292
rect 49700 32240 49752 32292
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 17500 31968 17552 32020
rect 19800 31968 19852 32020
rect 19892 31968 19944 32020
rect 20444 31968 20496 32020
rect 20904 31968 20956 32020
rect 38660 31968 38712 32020
rect 16488 31900 16540 31952
rect 16764 31832 16816 31884
rect 1676 31807 1728 31816
rect 1676 31773 1685 31807
rect 1685 31773 1719 31807
rect 1719 31773 1728 31807
rect 1676 31764 1728 31773
rect 17408 31807 17460 31816
rect 17408 31773 17417 31807
rect 17417 31773 17451 31807
rect 17451 31773 17460 31807
rect 17408 31764 17460 31773
rect 17500 31696 17552 31748
rect 17960 31832 18012 31884
rect 19340 31832 19392 31884
rect 22652 31900 22704 31952
rect 25872 31900 25924 31952
rect 33508 31900 33560 31952
rect 36176 31900 36228 31952
rect 23020 31832 23072 31884
rect 24400 31832 24452 31884
rect 18144 31696 18196 31748
rect 18328 31696 18380 31748
rect 19248 31696 19300 31748
rect 20720 31764 20772 31816
rect 20812 31764 20864 31816
rect 21916 31807 21968 31816
rect 20536 31696 20588 31748
rect 21916 31773 21925 31807
rect 21925 31773 21959 31807
rect 21959 31773 21968 31807
rect 21916 31764 21968 31773
rect 22192 31764 22244 31816
rect 22560 31696 22612 31748
rect 23296 31764 23348 31816
rect 25964 31832 26016 31884
rect 33876 31832 33928 31884
rect 42340 31900 42392 31952
rect 44456 31900 44508 31952
rect 44732 31900 44784 31952
rect 49240 31900 49292 31952
rect 23572 31696 23624 31748
rect 14372 31628 14424 31680
rect 25780 31696 25832 31748
rect 25964 31696 26016 31748
rect 31760 31696 31812 31748
rect 33968 31764 34020 31816
rect 34704 31764 34756 31816
rect 42432 31807 42484 31816
rect 42432 31773 42439 31807
rect 42439 31773 42484 31807
rect 42432 31764 42484 31773
rect 42616 31807 42668 31816
rect 42616 31773 42625 31807
rect 42625 31773 42659 31807
rect 42659 31773 42668 31807
rect 42616 31764 42668 31773
rect 26056 31628 26108 31680
rect 32036 31628 32088 31680
rect 33508 31696 33560 31748
rect 33048 31628 33100 31680
rect 33600 31628 33652 31680
rect 38476 31696 38528 31748
rect 43444 31764 43496 31816
rect 43996 31807 44048 31816
rect 43996 31773 44005 31807
rect 44005 31773 44039 31807
rect 44039 31773 44048 31807
rect 43996 31764 44048 31773
rect 44088 31807 44140 31816
rect 44088 31773 44098 31807
rect 44098 31773 44132 31807
rect 44132 31773 44140 31807
rect 44088 31764 44140 31773
rect 44180 31696 44232 31748
rect 46756 31832 46808 31884
rect 45836 31764 45888 31816
rect 47584 31764 47636 31816
rect 57428 31764 57480 31816
rect 58164 31807 58216 31816
rect 58164 31773 58173 31807
rect 58173 31773 58207 31807
rect 58207 31773 58216 31807
rect 58164 31764 58216 31773
rect 34060 31628 34112 31680
rect 53932 31628 53984 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 24584 31424 24636 31476
rect 17960 31356 18012 31408
rect 1676 31331 1728 31340
rect 1676 31297 1685 31331
rect 1685 31297 1719 31331
rect 1719 31297 1728 31331
rect 1676 31288 1728 31297
rect 18144 31331 18196 31340
rect 18144 31297 18153 31331
rect 18153 31297 18187 31331
rect 18187 31297 18196 31331
rect 18144 31288 18196 31297
rect 19064 31331 19116 31340
rect 19064 31297 19073 31331
rect 19073 31297 19107 31331
rect 19107 31297 19116 31331
rect 19064 31288 19116 31297
rect 19432 31288 19484 31340
rect 20444 31288 20496 31340
rect 25136 31399 25188 31408
rect 25136 31365 25145 31399
rect 25145 31365 25179 31399
rect 25179 31365 25188 31399
rect 25872 31399 25924 31408
rect 25136 31356 25188 31365
rect 25872 31365 25881 31399
rect 25881 31365 25915 31399
rect 25915 31365 25924 31399
rect 25872 31356 25924 31365
rect 32404 31424 32456 31476
rect 20536 31263 20588 31272
rect 20536 31229 20545 31263
rect 20545 31229 20579 31263
rect 20579 31229 20588 31263
rect 20536 31220 20588 31229
rect 22100 31220 22152 31272
rect 24952 31331 25004 31340
rect 24952 31297 24959 31331
rect 24959 31297 25004 31331
rect 24584 31220 24636 31272
rect 21548 31152 21600 31204
rect 24952 31288 25004 31297
rect 26056 31331 26108 31340
rect 25780 31220 25832 31272
rect 26056 31297 26065 31331
rect 26065 31297 26099 31331
rect 26099 31297 26108 31331
rect 26056 31288 26108 31297
rect 32036 31288 32088 31340
rect 33600 31288 33652 31340
rect 33784 31331 33836 31340
rect 33784 31297 33793 31331
rect 33793 31297 33827 31331
rect 33827 31297 33836 31331
rect 33784 31288 33836 31297
rect 34060 31331 34112 31340
rect 34060 31297 34069 31331
rect 34069 31297 34103 31331
rect 34103 31297 34112 31331
rect 34060 31288 34112 31297
rect 34796 31356 34848 31408
rect 35256 31399 35308 31408
rect 35256 31365 35265 31399
rect 35265 31365 35299 31399
rect 35299 31365 35308 31399
rect 35256 31356 35308 31365
rect 25964 31220 26016 31272
rect 26332 31263 26384 31272
rect 26332 31229 26341 31263
rect 26341 31229 26375 31263
rect 26375 31229 26384 31263
rect 26332 31220 26384 31229
rect 33140 31220 33192 31272
rect 35164 31331 35216 31340
rect 35164 31297 35171 31331
rect 35171 31297 35216 31331
rect 35164 31288 35216 31297
rect 35348 31331 35400 31340
rect 35348 31297 35357 31331
rect 35357 31297 35391 31331
rect 35391 31297 35400 31331
rect 35348 31288 35400 31297
rect 36268 31220 36320 31272
rect 37464 31220 37516 31272
rect 43076 31220 43128 31272
rect 52276 31220 52328 31272
rect 31116 31152 31168 31204
rect 44088 31152 44140 31204
rect 53012 31152 53064 31204
rect 23296 31084 23348 31136
rect 24584 31084 24636 31136
rect 29828 31084 29880 31136
rect 37280 31084 37332 31136
rect 42432 31084 42484 31136
rect 52920 31084 52972 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 6920 30880 6972 30932
rect 35348 30880 35400 30932
rect 35808 30880 35860 30932
rect 17960 30812 18012 30864
rect 18880 30812 18932 30864
rect 23572 30855 23624 30864
rect 17500 30787 17552 30796
rect 17500 30753 17509 30787
rect 17509 30753 17543 30787
rect 17543 30753 17552 30787
rect 17500 30744 17552 30753
rect 1676 30651 1728 30660
rect 1676 30617 1685 30651
rect 1685 30617 1719 30651
rect 1719 30617 1728 30651
rect 1676 30608 1728 30617
rect 17408 30608 17460 30660
rect 17776 30608 17828 30660
rect 18328 30676 18380 30728
rect 19432 30676 19484 30728
rect 20076 30744 20128 30796
rect 21548 30787 21600 30796
rect 21548 30753 21557 30787
rect 21557 30753 21591 30787
rect 21591 30753 21600 30787
rect 21548 30744 21600 30753
rect 19984 30719 20036 30728
rect 19984 30685 19993 30719
rect 19993 30685 20027 30719
rect 20027 30685 20036 30719
rect 19984 30676 20036 30685
rect 20536 30676 20588 30728
rect 20628 30676 20680 30728
rect 22192 30719 22244 30728
rect 16304 30540 16356 30592
rect 18144 30540 18196 30592
rect 18788 30540 18840 30592
rect 19340 30540 19392 30592
rect 20536 30540 20588 30592
rect 20996 30540 21048 30592
rect 22192 30685 22201 30719
rect 22201 30685 22235 30719
rect 22235 30685 22244 30719
rect 22192 30676 22244 30685
rect 23020 30719 23072 30728
rect 23020 30685 23029 30719
rect 23029 30685 23063 30719
rect 23063 30685 23072 30719
rect 23020 30676 23072 30685
rect 23296 30719 23348 30728
rect 23296 30685 23305 30719
rect 23305 30685 23339 30719
rect 23339 30685 23348 30719
rect 23296 30676 23348 30685
rect 23572 30821 23581 30855
rect 23581 30821 23615 30855
rect 23615 30821 23624 30855
rect 23572 30812 23624 30821
rect 30472 30787 30524 30796
rect 30472 30753 30481 30787
rect 30481 30753 30515 30787
rect 30515 30753 30524 30787
rect 30472 30744 30524 30753
rect 24584 30719 24636 30728
rect 24584 30685 24593 30719
rect 24593 30685 24627 30719
rect 24627 30685 24636 30719
rect 24584 30676 24636 30685
rect 24768 30719 24820 30728
rect 24768 30685 24777 30719
rect 24777 30685 24811 30719
rect 24811 30685 24820 30719
rect 24768 30676 24820 30685
rect 28540 30676 28592 30728
rect 29736 30651 29788 30660
rect 29736 30617 29745 30651
rect 29745 30617 29779 30651
rect 29779 30617 29788 30651
rect 29736 30608 29788 30617
rect 43812 30812 43864 30864
rect 31116 30744 31168 30796
rect 31760 30676 31812 30728
rect 35624 30676 35676 30728
rect 35900 30719 35952 30728
rect 35900 30685 35910 30719
rect 35910 30685 35944 30719
rect 35944 30685 35952 30719
rect 35900 30676 35952 30685
rect 36084 30719 36136 30728
rect 36084 30685 36093 30719
rect 36093 30685 36127 30719
rect 36127 30685 36136 30719
rect 36084 30676 36136 30685
rect 36268 30719 36320 30728
rect 36268 30685 36282 30719
rect 36282 30685 36316 30719
rect 36316 30685 36320 30719
rect 36912 30719 36964 30728
rect 36268 30676 36320 30685
rect 36912 30685 36921 30719
rect 36921 30685 36955 30719
rect 36955 30685 36964 30719
rect 36912 30676 36964 30685
rect 37004 30719 37056 30728
rect 37004 30685 37014 30719
rect 37014 30685 37048 30719
rect 37048 30685 37056 30719
rect 37004 30676 37056 30685
rect 37280 30719 37332 30728
rect 37280 30685 37289 30719
rect 37289 30685 37323 30719
rect 37323 30685 37332 30719
rect 37280 30676 37332 30685
rect 37464 30676 37516 30728
rect 38660 30676 38712 30728
rect 57980 30719 58032 30728
rect 57980 30685 57989 30719
rect 57989 30685 58023 30719
rect 58023 30685 58032 30719
rect 57980 30676 58032 30685
rect 22100 30540 22152 30592
rect 24860 30583 24912 30592
rect 24860 30549 24869 30583
rect 24869 30549 24903 30583
rect 24903 30549 24912 30583
rect 24860 30540 24912 30549
rect 27436 30540 27488 30592
rect 37556 30583 37608 30592
rect 37556 30549 37565 30583
rect 37565 30549 37599 30583
rect 37599 30549 37608 30583
rect 37556 30540 37608 30549
rect 58072 30583 58124 30592
rect 58072 30549 58081 30583
rect 58081 30549 58115 30583
rect 58115 30549 58124 30583
rect 58072 30540 58124 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 19616 30379 19668 30388
rect 19616 30345 19625 30379
rect 19625 30345 19659 30379
rect 19659 30345 19668 30379
rect 19616 30336 19668 30345
rect 20076 30336 20128 30388
rect 33784 30336 33836 30388
rect 36268 30336 36320 30388
rect 17500 30268 17552 30320
rect 17868 30311 17920 30320
rect 17868 30277 17877 30311
rect 17877 30277 17911 30311
rect 17911 30277 17920 30311
rect 20628 30311 20680 30320
rect 17868 30268 17920 30277
rect 18328 30243 18380 30252
rect 18328 30209 18337 30243
rect 18337 30209 18371 30243
rect 18371 30209 18380 30243
rect 18328 30200 18380 30209
rect 20076 30200 20128 30252
rect 20628 30277 20637 30311
rect 20637 30277 20671 30311
rect 20671 30277 20680 30311
rect 20628 30268 20680 30277
rect 23480 30268 23532 30320
rect 35624 30268 35676 30320
rect 36912 30336 36964 30388
rect 42892 30336 42944 30388
rect 43168 30336 43220 30388
rect 37556 30268 37608 30320
rect 19432 30132 19484 30184
rect 19984 30132 20036 30184
rect 19616 30064 19668 30116
rect 22192 30200 22244 30252
rect 42340 30200 42392 30252
rect 21916 30132 21968 30184
rect 23020 30132 23072 30184
rect 20996 30064 21048 30116
rect 37648 29996 37700 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 20444 29792 20496 29844
rect 34796 29792 34848 29844
rect 36820 29792 36872 29844
rect 43812 29835 43864 29844
rect 43812 29801 43821 29835
rect 43821 29801 43855 29835
rect 43855 29801 43864 29835
rect 43812 29792 43864 29801
rect 53472 29724 53524 29776
rect 6184 29656 6236 29708
rect 17684 29656 17736 29708
rect 22836 29656 22888 29708
rect 34796 29656 34848 29708
rect 34980 29656 35032 29708
rect 43076 29656 43128 29708
rect 15200 29631 15252 29640
rect 1860 29563 1912 29572
rect 1860 29529 1869 29563
rect 1869 29529 1903 29563
rect 1903 29529 1912 29563
rect 1860 29520 1912 29529
rect 15200 29597 15209 29631
rect 15209 29597 15243 29631
rect 15243 29597 15252 29631
rect 15200 29588 15252 29597
rect 17868 29588 17920 29640
rect 19156 29588 19208 29640
rect 19340 29588 19392 29640
rect 20444 29631 20496 29640
rect 18788 29520 18840 29572
rect 20444 29597 20453 29631
rect 20453 29597 20487 29631
rect 20487 29597 20496 29631
rect 20444 29588 20496 29597
rect 20996 29631 21048 29640
rect 20996 29597 21005 29631
rect 21005 29597 21039 29631
rect 21039 29597 21048 29631
rect 20996 29588 21048 29597
rect 34888 29631 34940 29640
rect 34888 29597 34897 29631
rect 34897 29597 34931 29631
rect 34931 29597 34940 29631
rect 34888 29588 34940 29597
rect 20720 29520 20772 29572
rect 34244 29520 34296 29572
rect 36176 29588 36228 29640
rect 43168 29631 43220 29640
rect 43168 29597 43177 29631
rect 43177 29597 43211 29631
rect 43211 29597 43220 29631
rect 43168 29588 43220 29597
rect 47216 29656 47268 29708
rect 58164 29699 58216 29708
rect 58164 29665 58173 29699
rect 58173 29665 58207 29699
rect 58207 29665 58216 29699
rect 58164 29656 58216 29665
rect 43444 29631 43496 29640
rect 43444 29597 43453 29631
rect 43453 29597 43487 29631
rect 43487 29597 43496 29631
rect 43444 29588 43496 29597
rect 46112 29588 46164 29640
rect 35072 29563 35124 29572
rect 35072 29529 35081 29563
rect 35081 29529 35115 29563
rect 35115 29529 35124 29563
rect 35072 29520 35124 29529
rect 44640 29520 44692 29572
rect 57060 29563 57112 29572
rect 57060 29529 57069 29563
rect 57069 29529 57103 29563
rect 57103 29529 57112 29563
rect 57060 29520 57112 29529
rect 18880 29452 18932 29504
rect 43628 29452 43680 29504
rect 57152 29495 57204 29504
rect 57152 29461 57161 29495
rect 57161 29461 57195 29495
rect 57195 29461 57204 29495
rect 57152 29452 57204 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 19432 29248 19484 29300
rect 24400 29291 24452 29300
rect 24400 29257 24409 29291
rect 24409 29257 24443 29291
rect 24443 29257 24452 29291
rect 24400 29248 24452 29257
rect 32864 29248 32916 29300
rect 35072 29248 35124 29300
rect 43076 29248 43128 29300
rect 49056 29248 49108 29300
rect 20444 29180 20496 29232
rect 34888 29180 34940 29232
rect 37280 29180 37332 29232
rect 2872 29112 2924 29164
rect 18420 29112 18472 29164
rect 18788 29155 18840 29164
rect 18788 29121 18797 29155
rect 18797 29121 18831 29155
rect 18831 29121 18840 29155
rect 18788 29112 18840 29121
rect 1768 29087 1820 29096
rect 1768 29053 1777 29087
rect 1777 29053 1811 29087
rect 1811 29053 1820 29087
rect 1768 29044 1820 29053
rect 18144 29044 18196 29096
rect 18328 29044 18380 29096
rect 19524 29112 19576 29164
rect 24124 29155 24176 29164
rect 24124 29121 24133 29155
rect 24133 29121 24167 29155
rect 24167 29121 24176 29155
rect 24124 29112 24176 29121
rect 24216 29155 24268 29164
rect 24216 29121 24225 29155
rect 24225 29121 24259 29155
rect 24259 29121 24268 29155
rect 24216 29112 24268 29121
rect 25320 29112 25372 29164
rect 31300 29112 31352 29164
rect 57152 29112 57204 29164
rect 19156 29044 19208 29096
rect 19616 29044 19668 29096
rect 26424 29044 26476 29096
rect 31024 29044 31076 29096
rect 18420 28908 18472 28960
rect 19064 28908 19116 28960
rect 20996 28976 21048 29028
rect 24308 28976 24360 29028
rect 27712 28976 27764 29028
rect 32956 28976 33008 29028
rect 39856 28976 39908 29028
rect 34152 28908 34204 28960
rect 41696 28908 41748 28960
rect 47216 28908 47268 28960
rect 52736 28908 52788 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 26148 28704 26200 28756
rect 41144 28704 41196 28756
rect 2872 28679 2924 28688
rect 2872 28645 2881 28679
rect 2881 28645 2915 28679
rect 2915 28645 2924 28679
rect 2872 28636 2924 28645
rect 16304 28636 16356 28688
rect 27160 28636 27212 28688
rect 35716 28636 35768 28688
rect 47584 28636 47636 28688
rect 37004 28568 37056 28620
rect 47952 28568 48004 28620
rect 1584 28543 1636 28552
rect 1584 28509 1593 28543
rect 1593 28509 1627 28543
rect 1627 28509 1636 28543
rect 1584 28500 1636 28509
rect 2504 28543 2556 28552
rect 2504 28509 2513 28543
rect 2513 28509 2547 28543
rect 2547 28509 2556 28543
rect 2504 28500 2556 28509
rect 18236 28500 18288 28552
rect 25412 28500 25464 28552
rect 42892 28500 42944 28552
rect 43996 28500 44048 28552
rect 1860 28475 1912 28484
rect 1860 28441 1869 28475
rect 1869 28441 1903 28475
rect 1903 28441 1912 28475
rect 1860 28432 1912 28441
rect 24952 28432 25004 28484
rect 31852 28432 31904 28484
rect 58164 28475 58216 28484
rect 58164 28441 58173 28475
rect 58173 28441 58207 28475
rect 58207 28441 58216 28475
rect 58164 28432 58216 28441
rect 23020 28364 23072 28416
rect 54760 28364 54812 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 1584 28160 1636 28212
rect 31852 28160 31904 28212
rect 44180 28160 44232 28212
rect 55312 28160 55364 28212
rect 56048 28160 56100 28212
rect 1400 28067 1452 28076
rect 1400 28033 1409 28067
rect 1409 28033 1443 28067
rect 1443 28033 1452 28067
rect 1400 28024 1452 28033
rect 2504 28067 2556 28076
rect 2504 28033 2513 28067
rect 2513 28033 2547 28067
rect 2547 28033 2556 28067
rect 2504 28024 2556 28033
rect 17960 28024 18012 28076
rect 1584 27999 1636 28008
rect 1584 27965 1593 27999
rect 1593 27965 1627 27999
rect 1627 27965 1636 27999
rect 1584 27956 1636 27965
rect 30380 27820 30432 27872
rect 33048 27820 33100 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 1400 27616 1452 27668
rect 18052 27616 18104 27668
rect 22008 27616 22060 27668
rect 44824 27616 44876 27668
rect 45652 27616 45704 27668
rect 17960 27548 18012 27600
rect 18880 27548 18932 27600
rect 18420 27480 18472 27532
rect 2228 27455 2280 27464
rect 2228 27421 2241 27455
rect 2241 27421 2280 27455
rect 2228 27412 2280 27421
rect 17960 27412 18012 27464
rect 19340 27480 19392 27532
rect 20536 27548 20588 27600
rect 24032 27548 24084 27600
rect 31944 27480 31996 27532
rect 32864 27480 32916 27532
rect 35900 27480 35952 27532
rect 42064 27480 42116 27532
rect 18788 27412 18840 27464
rect 57980 27455 58032 27464
rect 57980 27421 57989 27455
rect 57989 27421 58023 27455
rect 58023 27421 58032 27455
rect 57980 27412 58032 27421
rect 2504 27344 2556 27396
rect 18604 27387 18656 27396
rect 18604 27353 18613 27387
rect 18613 27353 18647 27387
rect 18647 27353 18656 27387
rect 18604 27344 18656 27353
rect 17868 27276 17920 27328
rect 20720 27344 20772 27396
rect 25320 27276 25372 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 37280 27072 37332 27124
rect 39580 27072 39632 27124
rect 18052 27047 18104 27056
rect 18052 27013 18061 27047
rect 18061 27013 18095 27047
rect 18095 27013 18104 27047
rect 18052 27004 18104 27013
rect 2504 26979 2556 26988
rect 2504 26945 2513 26979
rect 2513 26945 2547 26979
rect 2547 26945 2556 26979
rect 2504 26936 2556 26945
rect 1768 26911 1820 26920
rect 1768 26877 1777 26911
rect 1777 26877 1811 26911
rect 1811 26877 1820 26911
rect 1768 26868 1820 26877
rect 17868 26936 17920 26988
rect 18604 27004 18656 27056
rect 18236 26868 18288 26920
rect 19340 26936 19392 26988
rect 35716 27004 35768 27056
rect 48044 27004 48096 27056
rect 19248 26868 19300 26920
rect 20168 26936 20220 26988
rect 20720 26936 20772 26988
rect 24676 26936 24728 26988
rect 46480 26936 46532 26988
rect 17592 26800 17644 26852
rect 26608 26868 26660 26920
rect 49792 26868 49844 26920
rect 21456 26800 21508 26852
rect 22192 26732 22244 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 18604 26435 18656 26444
rect 18604 26401 18613 26435
rect 18613 26401 18647 26435
rect 18647 26401 18656 26435
rect 18604 26392 18656 26401
rect 20168 26435 20220 26444
rect 20168 26401 20177 26435
rect 20177 26401 20211 26435
rect 20211 26401 20220 26435
rect 20168 26392 20220 26401
rect 25872 26392 25924 26444
rect 2504 26367 2556 26376
rect 2504 26333 2513 26367
rect 2513 26333 2547 26367
rect 2547 26333 2556 26367
rect 2504 26324 2556 26333
rect 2596 26367 2648 26376
rect 2596 26333 2606 26367
rect 2606 26333 2640 26367
rect 2640 26333 2648 26367
rect 2596 26324 2648 26333
rect 18328 26324 18380 26376
rect 19432 26367 19484 26376
rect 19432 26333 19441 26367
rect 19441 26333 19475 26367
rect 19475 26333 19484 26367
rect 19432 26324 19484 26333
rect 20076 26324 20128 26376
rect 58716 26460 58768 26512
rect 28356 26392 28408 26444
rect 58164 26435 58216 26444
rect 58164 26401 58173 26435
rect 58173 26401 58207 26435
rect 58207 26401 58216 26435
rect 58164 26392 58216 26401
rect 1860 26299 1912 26308
rect 1860 26265 1869 26299
rect 1869 26265 1903 26299
rect 1903 26265 1912 26299
rect 1860 26256 1912 26265
rect 26148 26299 26200 26308
rect 26148 26265 26157 26299
rect 26157 26265 26191 26299
rect 26191 26265 26200 26299
rect 26148 26256 26200 26265
rect 26792 26256 26844 26308
rect 40408 26324 40460 26376
rect 27436 26299 27488 26308
rect 27436 26265 27445 26299
rect 27445 26265 27479 26299
rect 27479 26265 27488 26299
rect 27436 26256 27488 26265
rect 25688 26231 25740 26240
rect 25688 26197 25697 26231
rect 25697 26197 25731 26231
rect 25731 26197 25740 26231
rect 25688 26188 25740 26197
rect 26884 26188 26936 26240
rect 58348 26188 58400 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 23388 25984 23440 26036
rect 24860 25984 24912 26036
rect 25872 25916 25924 25968
rect 2688 25848 2740 25900
rect 20536 25891 20588 25900
rect 20536 25857 20545 25891
rect 20545 25857 20579 25891
rect 20579 25857 20588 25891
rect 20536 25848 20588 25857
rect 21088 25848 21140 25900
rect 28448 25916 28500 25968
rect 29828 25916 29880 25968
rect 1768 25823 1820 25832
rect 1768 25789 1777 25823
rect 1777 25789 1811 25823
rect 1811 25789 1820 25823
rect 1768 25780 1820 25789
rect 20444 25780 20496 25832
rect 25872 25780 25924 25832
rect 26056 25823 26108 25832
rect 26056 25789 26065 25823
rect 26065 25789 26099 25823
rect 26099 25789 26108 25823
rect 27988 25848 28040 25900
rect 58072 25891 58124 25900
rect 58072 25857 58081 25891
rect 58081 25857 58115 25891
rect 58115 25857 58124 25891
rect 58072 25848 58124 25857
rect 26056 25780 26108 25789
rect 29092 25780 29144 25832
rect 58440 25712 58492 25764
rect 20076 25644 20128 25696
rect 25596 25687 25648 25696
rect 25596 25653 25605 25687
rect 25605 25653 25639 25687
rect 25639 25653 25648 25687
rect 25596 25644 25648 25653
rect 27804 25687 27856 25696
rect 27804 25653 27813 25687
rect 27813 25653 27847 25687
rect 27847 25653 27856 25687
rect 27804 25644 27856 25653
rect 31576 25644 31628 25696
rect 58256 25687 58308 25696
rect 58256 25653 58265 25687
rect 58265 25653 58299 25687
rect 58299 25653 58308 25687
rect 58256 25644 58308 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 2688 25483 2740 25492
rect 2688 25449 2697 25483
rect 2697 25449 2731 25483
rect 2731 25449 2740 25483
rect 2688 25440 2740 25449
rect 19248 25440 19300 25492
rect 19984 25440 20036 25492
rect 2504 25372 2556 25424
rect 1584 25279 1636 25288
rect 1584 25245 1593 25279
rect 1593 25245 1627 25279
rect 1627 25245 1636 25279
rect 1584 25236 1636 25245
rect 15200 25304 15252 25356
rect 16488 25347 16540 25356
rect 16488 25313 16497 25347
rect 16497 25313 16531 25347
rect 16531 25313 16540 25347
rect 16488 25304 16540 25313
rect 20444 25304 20496 25356
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 17224 25236 17276 25288
rect 20168 25236 20220 25288
rect 26884 25440 26936 25492
rect 27804 25440 27856 25492
rect 55496 25440 55548 25492
rect 55588 25440 55640 25492
rect 58900 25440 58952 25492
rect 36636 25372 36688 25424
rect 58256 25372 58308 25424
rect 30196 25304 30248 25356
rect 24952 25279 25004 25288
rect 24952 25245 24961 25279
rect 24961 25245 24995 25279
rect 24995 25245 25004 25279
rect 24952 25236 25004 25245
rect 29000 25279 29052 25288
rect 29000 25245 29009 25279
rect 29009 25245 29043 25279
rect 29043 25245 29052 25279
rect 29000 25236 29052 25245
rect 29460 25236 29512 25288
rect 29828 25236 29880 25288
rect 55772 25236 55824 25288
rect 56048 25279 56100 25288
rect 56048 25245 56057 25279
rect 56057 25245 56091 25279
rect 56091 25245 56100 25279
rect 56048 25236 56100 25245
rect 56876 25279 56928 25288
rect 56876 25245 56885 25279
rect 56885 25245 56919 25279
rect 56919 25245 56928 25279
rect 56876 25236 56928 25245
rect 19984 25168 20036 25220
rect 21272 25168 21324 25220
rect 25688 25168 25740 25220
rect 26240 25168 26292 25220
rect 27528 25168 27580 25220
rect 29092 25168 29144 25220
rect 53840 25168 53892 25220
rect 58164 25211 58216 25220
rect 58164 25177 58173 25211
rect 58173 25177 58207 25211
rect 58207 25177 58216 25211
rect 58164 25168 58216 25177
rect 19248 25100 19300 25152
rect 20628 25100 20680 25152
rect 21364 25143 21416 25152
rect 21364 25109 21373 25143
rect 21373 25109 21407 25143
rect 21407 25109 21416 25143
rect 21364 25100 21416 25109
rect 22836 25100 22888 25152
rect 26148 25100 26200 25152
rect 28540 25143 28592 25152
rect 28540 25109 28549 25143
rect 28549 25109 28583 25143
rect 28583 25109 28592 25143
rect 28540 25100 28592 25109
rect 30104 25143 30156 25152
rect 30104 25109 30113 25143
rect 30113 25109 30147 25143
rect 30147 25109 30156 25143
rect 30104 25100 30156 25109
rect 56324 25100 56376 25152
rect 57152 25100 57204 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 1584 24896 1636 24948
rect 15200 24760 15252 24812
rect 15568 24760 15620 24812
rect 16120 24760 16172 24812
rect 16488 24760 16540 24812
rect 19340 24803 19392 24812
rect 19340 24769 19349 24803
rect 19349 24769 19383 24803
rect 19383 24769 19392 24803
rect 19340 24760 19392 24769
rect 20352 24896 20404 24948
rect 20536 24896 20588 24948
rect 56048 24939 56100 24948
rect 20168 24760 20220 24812
rect 21364 24760 21416 24812
rect 22468 24803 22520 24812
rect 19708 24692 19760 24744
rect 22468 24769 22477 24803
rect 22477 24769 22511 24803
rect 22511 24769 22520 24803
rect 22468 24760 22520 24769
rect 23572 24803 23624 24812
rect 23204 24692 23256 24744
rect 23572 24769 23581 24803
rect 23581 24769 23615 24803
rect 23615 24769 23624 24803
rect 23572 24760 23624 24769
rect 26424 24803 26476 24812
rect 26424 24769 26433 24803
rect 26433 24769 26467 24803
rect 26467 24769 26476 24803
rect 26424 24760 26476 24769
rect 23940 24692 23992 24744
rect 19156 24556 19208 24608
rect 19432 24556 19484 24608
rect 22560 24624 22612 24676
rect 24216 24624 24268 24676
rect 24308 24624 24360 24676
rect 27252 24760 27304 24812
rect 29920 24828 29972 24880
rect 31392 24871 31444 24880
rect 31392 24837 31401 24871
rect 31401 24837 31435 24871
rect 31435 24837 31444 24871
rect 31392 24828 31444 24837
rect 56048 24905 56057 24939
rect 56057 24905 56091 24939
rect 56091 24905 56100 24939
rect 56048 24896 56100 24905
rect 56876 24896 56928 24948
rect 27620 24692 27672 24744
rect 21272 24556 21324 24608
rect 22744 24556 22796 24608
rect 24676 24556 24728 24608
rect 26056 24556 26108 24608
rect 27620 24556 27672 24608
rect 29828 24803 29880 24812
rect 29828 24769 29862 24803
rect 29862 24769 29880 24803
rect 29828 24760 29880 24769
rect 32588 24803 32640 24812
rect 28908 24692 28960 24744
rect 32588 24769 32597 24803
rect 32597 24769 32631 24803
rect 32631 24769 32640 24803
rect 32588 24760 32640 24769
rect 55588 24828 55640 24880
rect 31668 24692 31720 24744
rect 31852 24692 31904 24744
rect 32864 24760 32916 24812
rect 36084 24760 36136 24812
rect 37004 24760 37056 24812
rect 45284 24760 45336 24812
rect 45468 24803 45520 24812
rect 45468 24769 45477 24803
rect 45477 24769 45511 24803
rect 45511 24769 45520 24803
rect 45468 24760 45520 24769
rect 51172 24760 51224 24812
rect 55312 24760 55364 24812
rect 55496 24803 55548 24812
rect 55496 24769 55505 24803
rect 55505 24769 55539 24803
rect 55539 24769 55548 24803
rect 55496 24760 55548 24769
rect 33048 24692 33100 24744
rect 45744 24692 45796 24744
rect 28908 24556 28960 24608
rect 29092 24599 29144 24608
rect 29092 24565 29101 24599
rect 29101 24565 29135 24599
rect 29135 24565 29144 24599
rect 29092 24556 29144 24565
rect 32588 24624 32640 24676
rect 30472 24556 30524 24608
rect 30840 24556 30892 24608
rect 32312 24599 32364 24608
rect 32312 24565 32321 24599
rect 32321 24565 32355 24599
rect 32355 24565 32364 24599
rect 32312 24556 32364 24565
rect 46204 24624 46256 24676
rect 45008 24556 45060 24608
rect 45284 24556 45336 24608
rect 51816 24692 51868 24744
rect 54116 24692 54168 24744
rect 55128 24692 55180 24744
rect 56232 24760 56284 24812
rect 56508 24803 56560 24812
rect 56508 24769 56517 24803
rect 56517 24769 56551 24803
rect 56551 24769 56560 24803
rect 56508 24760 56560 24769
rect 56692 24803 56744 24812
rect 56692 24769 56701 24803
rect 56701 24769 56735 24803
rect 56735 24769 56744 24803
rect 56876 24803 56928 24812
rect 56692 24760 56744 24769
rect 56876 24769 56885 24803
rect 56885 24769 56919 24803
rect 56919 24769 56928 24803
rect 56876 24760 56928 24769
rect 58072 24803 58124 24812
rect 46388 24624 46440 24676
rect 55036 24624 55088 24676
rect 57428 24692 57480 24744
rect 58072 24769 58081 24803
rect 58081 24769 58115 24803
rect 58115 24769 58124 24803
rect 58072 24760 58124 24769
rect 58348 24692 58400 24744
rect 50068 24556 50120 24608
rect 54484 24556 54536 24608
rect 55772 24556 55824 24608
rect 56232 24624 56284 24676
rect 56876 24624 56928 24676
rect 56692 24556 56744 24608
rect 58256 24599 58308 24608
rect 58256 24565 58265 24599
rect 58265 24565 58299 24599
rect 58299 24565 58308 24599
rect 58256 24556 58308 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19432 24216 19484 24268
rect 20168 24352 20220 24404
rect 13084 24148 13136 24200
rect 17500 24191 17552 24200
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 17500 24148 17552 24157
rect 17684 24148 17736 24200
rect 19248 24148 19300 24200
rect 20076 24148 20128 24200
rect 1860 24123 1912 24132
rect 1860 24089 1869 24123
rect 1869 24089 1903 24123
rect 1903 24089 1912 24123
rect 1860 24080 1912 24089
rect 16856 24123 16908 24132
rect 16856 24089 16865 24123
rect 16865 24089 16899 24123
rect 16899 24089 16908 24123
rect 16856 24080 16908 24089
rect 17776 24080 17828 24132
rect 22560 24284 22612 24336
rect 22652 24284 22704 24336
rect 21456 24216 21508 24268
rect 21180 24148 21232 24200
rect 21548 24191 21600 24200
rect 21548 24157 21557 24191
rect 21557 24157 21591 24191
rect 21591 24157 21600 24191
rect 21548 24148 21600 24157
rect 23020 24148 23072 24200
rect 19708 24012 19760 24064
rect 21088 24012 21140 24064
rect 24952 24352 25004 24404
rect 26424 24352 26476 24404
rect 29000 24352 29052 24404
rect 30012 24352 30064 24404
rect 30748 24352 30800 24404
rect 30932 24352 30984 24404
rect 40040 24352 40092 24404
rect 27160 24284 27212 24336
rect 29736 24284 29788 24336
rect 29920 24284 29972 24336
rect 35624 24284 35676 24336
rect 58256 24352 58308 24404
rect 44640 24327 44692 24336
rect 44640 24293 44649 24327
rect 44649 24293 44683 24327
rect 44683 24293 44692 24327
rect 44640 24284 44692 24293
rect 27068 24216 27120 24268
rect 29644 24216 29696 24268
rect 44824 24216 44876 24268
rect 45008 24216 45060 24268
rect 25596 24148 25648 24200
rect 27528 24148 27580 24200
rect 34796 24148 34848 24200
rect 44548 24148 44600 24200
rect 50068 24148 50120 24200
rect 50896 24148 50948 24200
rect 51540 24216 51592 24268
rect 51632 24191 51684 24200
rect 21824 24012 21876 24064
rect 22284 24012 22336 24064
rect 23020 24012 23072 24064
rect 23204 24055 23256 24064
rect 23204 24021 23213 24055
rect 23213 24021 23247 24055
rect 23247 24021 23256 24055
rect 23204 24012 23256 24021
rect 23296 24055 23348 24064
rect 23296 24021 23305 24055
rect 23305 24021 23339 24055
rect 23339 24021 23348 24055
rect 23296 24012 23348 24021
rect 25136 24012 25188 24064
rect 25228 24012 25280 24064
rect 25964 24055 26016 24064
rect 25964 24021 25973 24055
rect 25973 24021 26007 24055
rect 26007 24021 26016 24055
rect 25964 24012 26016 24021
rect 31116 24080 31168 24132
rect 32312 24080 32364 24132
rect 44456 24080 44508 24132
rect 50804 24080 50856 24132
rect 51356 24080 51408 24132
rect 51632 24157 51641 24191
rect 51641 24157 51675 24191
rect 51675 24157 51684 24191
rect 51632 24148 51684 24157
rect 52552 24191 52604 24200
rect 52552 24157 52561 24191
rect 52561 24157 52595 24191
rect 52595 24157 52604 24191
rect 52552 24148 52604 24157
rect 55864 24284 55916 24336
rect 57428 24327 57480 24336
rect 57428 24293 57437 24327
rect 57437 24293 57471 24327
rect 57471 24293 57480 24327
rect 57428 24284 57480 24293
rect 54484 24259 54536 24268
rect 54484 24225 54493 24259
rect 54493 24225 54527 24259
rect 54527 24225 54536 24259
rect 54484 24216 54536 24225
rect 54668 24191 54720 24200
rect 54668 24157 54677 24191
rect 54677 24157 54711 24191
rect 54711 24157 54720 24191
rect 54668 24148 54720 24157
rect 56048 24191 56100 24200
rect 56048 24157 56057 24191
rect 56057 24157 56091 24191
rect 56091 24157 56100 24191
rect 56048 24148 56100 24157
rect 56324 24191 56376 24200
rect 56324 24157 56358 24191
rect 56358 24157 56376 24191
rect 56324 24148 56376 24157
rect 57888 24191 57940 24200
rect 57888 24157 57897 24191
rect 57897 24157 57931 24191
rect 57931 24157 57940 24191
rect 57888 24148 57940 24157
rect 51816 24123 51868 24132
rect 51816 24089 51825 24123
rect 51825 24089 51859 24123
rect 51859 24089 51868 24123
rect 51816 24080 51868 24089
rect 53288 24080 53340 24132
rect 54024 24080 54076 24132
rect 27988 24012 28040 24064
rect 32680 24012 32732 24064
rect 43352 24012 43404 24064
rect 44640 24012 44692 24064
rect 50620 24012 50672 24064
rect 53104 24012 53156 24064
rect 54852 24055 54904 24064
rect 54852 24021 54861 24055
rect 54861 24021 54895 24055
rect 54895 24021 54904 24055
rect 54852 24012 54904 24021
rect 55036 24080 55088 24132
rect 59084 24148 59136 24200
rect 58164 24123 58216 24132
rect 58164 24089 58173 24123
rect 58173 24089 58207 24123
rect 58207 24089 58216 24123
rect 58164 24080 58216 24089
rect 57980 24012 58032 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 19984 23808 20036 23860
rect 20628 23851 20680 23860
rect 20628 23817 20637 23851
rect 20637 23817 20671 23851
rect 20671 23817 20680 23851
rect 20628 23808 20680 23817
rect 22284 23851 22336 23860
rect 22284 23817 22293 23851
rect 22293 23817 22327 23851
rect 22327 23817 22336 23851
rect 22284 23808 22336 23817
rect 15200 23740 15252 23792
rect 1768 23647 1820 23656
rect 1768 23613 1777 23647
rect 1777 23613 1811 23647
rect 1811 23613 1820 23647
rect 1768 23604 1820 23613
rect 17592 23740 17644 23792
rect 19064 23740 19116 23792
rect 19248 23740 19300 23792
rect 27068 23808 27120 23860
rect 27252 23851 27304 23860
rect 27252 23817 27261 23851
rect 27261 23817 27295 23851
rect 27295 23817 27304 23851
rect 27252 23808 27304 23817
rect 27528 23808 27580 23860
rect 29920 23808 29972 23860
rect 31116 23851 31168 23860
rect 15568 23715 15620 23724
rect 15568 23681 15577 23715
rect 15577 23681 15611 23715
rect 15611 23681 15620 23715
rect 15568 23672 15620 23681
rect 17776 23672 17828 23724
rect 18144 23715 18196 23724
rect 18144 23681 18153 23715
rect 18153 23681 18187 23715
rect 18187 23681 18196 23715
rect 18144 23672 18196 23681
rect 21824 23672 21876 23724
rect 13912 23647 13964 23656
rect 13912 23613 13921 23647
rect 13921 23613 13955 23647
rect 13955 23613 13964 23647
rect 13912 23604 13964 23613
rect 20444 23604 20496 23656
rect 22100 23604 22152 23656
rect 22744 23715 22796 23724
rect 22744 23681 22753 23715
rect 22753 23681 22787 23715
rect 22787 23681 22796 23715
rect 22744 23672 22796 23681
rect 23204 23672 23256 23724
rect 24216 23740 24268 23792
rect 27160 23740 27212 23792
rect 30104 23740 30156 23792
rect 31116 23817 31125 23851
rect 31125 23817 31159 23851
rect 31159 23817 31168 23851
rect 31116 23808 31168 23817
rect 32680 23783 32732 23792
rect 32680 23749 32689 23783
rect 32689 23749 32723 23783
rect 32723 23749 32732 23783
rect 32680 23740 32732 23749
rect 22652 23647 22704 23656
rect 22652 23613 22661 23647
rect 22661 23613 22695 23647
rect 22695 23613 22704 23647
rect 22652 23604 22704 23613
rect 25044 23604 25096 23656
rect 20536 23536 20588 23588
rect 19800 23468 19852 23520
rect 21456 23468 21508 23520
rect 21732 23468 21784 23520
rect 24308 23468 24360 23520
rect 27896 23715 27948 23724
rect 27896 23681 27905 23715
rect 27905 23681 27939 23715
rect 27939 23681 27948 23715
rect 27896 23672 27948 23681
rect 27988 23672 28040 23724
rect 29000 23672 29052 23724
rect 31300 23672 31352 23724
rect 29736 23604 29788 23656
rect 30104 23604 30156 23656
rect 31576 23715 31628 23724
rect 31576 23681 31585 23715
rect 31585 23681 31619 23715
rect 31619 23681 31628 23715
rect 31576 23672 31628 23681
rect 31760 23715 31812 23724
rect 31760 23681 31769 23715
rect 31769 23681 31803 23715
rect 31803 23681 31812 23715
rect 31760 23672 31812 23681
rect 32864 23672 32916 23724
rect 31852 23604 31904 23656
rect 32128 23604 32180 23656
rect 36176 23808 36228 23860
rect 40408 23851 40460 23860
rect 40408 23817 40417 23851
rect 40417 23817 40451 23851
rect 40451 23817 40460 23851
rect 40408 23808 40460 23817
rect 56508 23808 56560 23860
rect 57520 23851 57572 23860
rect 57520 23817 57529 23851
rect 57529 23817 57563 23851
rect 57563 23817 57572 23851
rect 57520 23808 57572 23817
rect 28264 23579 28316 23588
rect 28264 23545 28273 23579
rect 28273 23545 28307 23579
rect 28307 23545 28316 23579
rect 28264 23536 28316 23545
rect 30932 23536 30984 23588
rect 29092 23468 29144 23520
rect 31668 23468 31720 23520
rect 32680 23536 32732 23588
rect 34704 23672 34756 23724
rect 36452 23715 36504 23724
rect 36452 23681 36461 23715
rect 36461 23681 36495 23715
rect 36495 23681 36504 23715
rect 36452 23672 36504 23681
rect 38384 23715 38436 23724
rect 35900 23604 35952 23656
rect 38384 23681 38393 23715
rect 38393 23681 38427 23715
rect 38427 23681 38436 23715
rect 38384 23672 38436 23681
rect 39120 23672 39172 23724
rect 41880 23715 41932 23724
rect 41880 23681 41889 23715
rect 41889 23681 41923 23715
rect 41923 23681 41932 23715
rect 41880 23672 41932 23681
rect 44364 23672 44416 23724
rect 44640 23715 44692 23724
rect 44640 23681 44649 23715
rect 44649 23681 44683 23715
rect 44683 23681 44692 23715
rect 44640 23672 44692 23681
rect 52552 23740 52604 23792
rect 50620 23715 50672 23724
rect 50620 23681 50654 23715
rect 50654 23681 50672 23715
rect 37832 23604 37884 23656
rect 38752 23604 38804 23656
rect 38936 23604 38988 23656
rect 40408 23604 40460 23656
rect 44548 23604 44600 23656
rect 50620 23672 50672 23681
rect 53104 23715 53156 23724
rect 53104 23681 53113 23715
rect 53113 23681 53147 23715
rect 53147 23681 53156 23715
rect 53104 23672 53156 23681
rect 53288 23715 53340 23724
rect 53288 23681 53297 23715
rect 53297 23681 53331 23715
rect 53331 23681 53340 23715
rect 53288 23672 53340 23681
rect 56048 23740 56100 23792
rect 54852 23672 54904 23724
rect 56876 23740 56928 23792
rect 56416 23715 56468 23724
rect 56416 23681 56450 23715
rect 56450 23681 56468 23715
rect 56416 23672 56468 23681
rect 52000 23604 52052 23656
rect 35072 23579 35124 23588
rect 35072 23545 35081 23579
rect 35081 23545 35115 23579
rect 35115 23545 35124 23579
rect 35072 23536 35124 23545
rect 35440 23536 35492 23588
rect 35808 23536 35860 23588
rect 40040 23536 40092 23588
rect 51724 23579 51776 23588
rect 34796 23468 34848 23520
rect 36728 23468 36780 23520
rect 39028 23468 39080 23520
rect 43996 23511 44048 23520
rect 43996 23477 44005 23511
rect 44005 23477 44039 23511
rect 44039 23477 44048 23511
rect 43996 23468 44048 23477
rect 44456 23511 44508 23520
rect 44456 23477 44465 23511
rect 44465 23477 44499 23511
rect 44499 23477 44508 23511
rect 44456 23468 44508 23477
rect 51724 23545 51733 23579
rect 51733 23545 51767 23579
rect 51767 23545 51776 23579
rect 51724 23536 51776 23545
rect 54024 23468 54076 23520
rect 54392 23468 54444 23520
rect 57796 23468 57848 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19800 23307 19852 23316
rect 19800 23273 19809 23307
rect 19809 23273 19843 23307
rect 19843 23273 19852 23307
rect 19800 23264 19852 23273
rect 22468 23264 22520 23316
rect 24768 23264 24820 23316
rect 26240 23264 26292 23316
rect 19340 23196 19392 23248
rect 20536 23196 20588 23248
rect 17592 23128 17644 23180
rect 18880 23171 18932 23180
rect 13912 23060 13964 23112
rect 15936 23103 15988 23112
rect 15936 23069 15945 23103
rect 15945 23069 15979 23103
rect 15979 23069 15988 23103
rect 15936 23060 15988 23069
rect 1860 23035 1912 23044
rect 1860 23001 1869 23035
rect 1869 23001 1903 23035
rect 1903 23001 1912 23035
rect 1860 22992 1912 23001
rect 17776 22992 17828 23044
rect 18880 23137 18889 23171
rect 18889 23137 18923 23171
rect 18923 23137 18932 23171
rect 18880 23128 18932 23137
rect 19800 23060 19852 23112
rect 21180 23128 21232 23180
rect 20812 23060 20864 23112
rect 25044 23196 25096 23248
rect 29828 23264 29880 23316
rect 24768 23128 24820 23180
rect 24584 23103 24636 23112
rect 24584 23069 24593 23103
rect 24593 23069 24627 23103
rect 24627 23069 24636 23103
rect 24584 23060 24636 23069
rect 25320 23103 25372 23112
rect 25320 23069 25329 23103
rect 25329 23069 25363 23103
rect 25363 23069 25372 23103
rect 25320 23060 25372 23069
rect 25688 23060 25740 23112
rect 26148 23128 26200 23180
rect 26056 23103 26108 23112
rect 26056 23069 26065 23103
rect 26065 23069 26099 23103
rect 26099 23069 26108 23103
rect 26056 23060 26108 23069
rect 27896 23196 27948 23248
rect 29920 23196 29972 23248
rect 30104 23196 30156 23248
rect 37832 23196 37884 23248
rect 38108 23196 38160 23248
rect 38384 23264 38436 23316
rect 40592 23264 40644 23316
rect 41880 23264 41932 23316
rect 42524 23307 42576 23316
rect 42524 23273 42533 23307
rect 42533 23273 42567 23307
rect 42567 23273 42576 23307
rect 42524 23264 42576 23273
rect 44364 23264 44416 23316
rect 50896 23307 50948 23316
rect 50896 23273 50905 23307
rect 50905 23273 50939 23307
rect 50939 23273 50948 23307
rect 50896 23264 50948 23273
rect 54668 23264 54720 23316
rect 58348 23264 58400 23316
rect 19432 22924 19484 22976
rect 20352 22992 20404 23044
rect 20444 22992 20496 23044
rect 20536 22924 20588 22976
rect 20904 22992 20956 23044
rect 21548 22992 21600 23044
rect 23848 22992 23900 23044
rect 28540 23060 28592 23112
rect 29644 23060 29696 23112
rect 30196 23103 30248 23112
rect 30196 23069 30210 23103
rect 30210 23069 30244 23103
rect 30244 23069 30248 23103
rect 30196 23060 30248 23069
rect 30380 23103 30432 23112
rect 30380 23069 30389 23103
rect 30389 23069 30423 23103
rect 30423 23069 30432 23103
rect 31760 23128 31812 23180
rect 31024 23103 31076 23112
rect 30380 23060 30432 23069
rect 31024 23069 31033 23103
rect 31033 23069 31067 23103
rect 31067 23069 31076 23103
rect 31024 23060 31076 23069
rect 35440 23060 35492 23112
rect 36176 23128 36228 23180
rect 40316 23196 40368 23248
rect 53840 23196 53892 23248
rect 22284 22924 22336 22976
rect 22928 22967 22980 22976
rect 22928 22933 22937 22967
rect 22937 22933 22971 22967
rect 22971 22933 22980 22967
rect 22928 22924 22980 22933
rect 25596 22924 25648 22976
rect 33876 22992 33928 23044
rect 34336 22992 34388 23044
rect 34612 22992 34664 23044
rect 26884 22924 26936 22976
rect 34152 22967 34204 22976
rect 34152 22933 34161 22967
rect 34161 22933 34195 22967
rect 34195 22933 34204 22967
rect 34152 22924 34204 22933
rect 36544 23103 36596 23112
rect 36544 23069 36553 23103
rect 36553 23069 36587 23103
rect 36587 23069 36596 23103
rect 36544 23060 36596 23069
rect 37832 23060 37884 23112
rect 39488 23060 39540 23112
rect 40500 23128 40552 23180
rect 36268 22992 36320 23044
rect 37004 22992 37056 23044
rect 37280 22992 37332 23044
rect 38844 23035 38896 23044
rect 38844 23001 38853 23035
rect 38853 23001 38887 23035
rect 38887 23001 38896 23035
rect 38844 22992 38896 23001
rect 36176 22924 36228 22976
rect 39672 22924 39724 22976
rect 39764 22924 39816 22976
rect 40224 22924 40276 22976
rect 43996 23128 44048 23180
rect 54392 23171 54444 23180
rect 42800 23060 42852 23112
rect 43352 23103 43404 23112
rect 43352 23069 43394 23103
rect 43394 23069 43404 23103
rect 43352 23060 43404 23069
rect 43720 23060 43772 23112
rect 43904 23103 43956 23112
rect 43904 23069 43913 23103
rect 43913 23069 43947 23103
rect 43947 23069 43956 23103
rect 43904 23060 43956 23069
rect 44364 23060 44416 23112
rect 48136 23060 48188 23112
rect 50712 23103 50764 23112
rect 50712 23069 50721 23103
rect 50721 23069 50755 23103
rect 50755 23069 50764 23103
rect 50712 23060 50764 23069
rect 53932 23103 53984 23112
rect 53932 23069 53941 23103
rect 53941 23069 53975 23103
rect 53975 23069 53984 23103
rect 53932 23060 53984 23069
rect 54116 23103 54168 23112
rect 54116 23069 54125 23103
rect 54125 23069 54159 23103
rect 54159 23069 54168 23103
rect 54116 23060 54168 23069
rect 54392 23137 54401 23171
rect 54401 23137 54435 23171
rect 54435 23137 54444 23171
rect 54392 23128 54444 23137
rect 56508 23128 56560 23180
rect 56876 23171 56928 23180
rect 56876 23137 56885 23171
rect 56885 23137 56919 23171
rect 56919 23137 56928 23171
rect 56876 23128 56928 23137
rect 56048 23060 56100 23112
rect 40500 23035 40552 23044
rect 40500 23001 40535 23035
rect 40535 23001 40552 23035
rect 40500 22992 40552 23001
rect 47860 22992 47912 23044
rect 40684 22924 40736 22976
rect 41420 22924 41472 22976
rect 49976 22992 50028 23044
rect 51724 22992 51776 23044
rect 55956 23035 56008 23044
rect 55956 23001 55965 23035
rect 55965 23001 55999 23035
rect 55999 23001 56008 23035
rect 55956 22992 56008 23001
rect 50712 22924 50764 22976
rect 53380 22967 53432 22976
rect 53380 22933 53389 22967
rect 53389 22933 53423 22967
rect 53423 22933 53432 22967
rect 53380 22924 53432 22933
rect 53932 22924 53984 22976
rect 55128 22924 55180 22976
rect 56324 23103 56376 23112
rect 56324 23069 56338 23103
rect 56338 23069 56372 23103
rect 56372 23069 56376 23103
rect 57152 23103 57204 23112
rect 56324 23060 56376 23069
rect 57152 23069 57186 23103
rect 57186 23069 57204 23103
rect 57152 23060 57204 23069
rect 57520 22992 57572 23044
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 17316 22720 17368 22772
rect 17500 22763 17552 22772
rect 17500 22729 17509 22763
rect 17509 22729 17543 22763
rect 17543 22729 17552 22763
rect 17500 22720 17552 22729
rect 19432 22720 19484 22772
rect 23848 22763 23900 22772
rect 13544 22584 13596 22636
rect 19340 22652 19392 22704
rect 20352 22652 20404 22704
rect 1768 22559 1820 22568
rect 1768 22525 1777 22559
rect 1777 22525 1811 22559
rect 1811 22525 1820 22559
rect 1768 22516 1820 22525
rect 17500 22584 17552 22636
rect 17684 22584 17736 22636
rect 17868 22584 17920 22636
rect 18880 22584 18932 22636
rect 21364 22627 21416 22636
rect 21364 22593 21373 22627
rect 21373 22593 21407 22627
rect 21407 22593 21416 22627
rect 21364 22584 21416 22593
rect 18236 22516 18288 22568
rect 20536 22516 20588 22568
rect 21824 22584 21876 22636
rect 22928 22652 22980 22704
rect 23848 22729 23857 22763
rect 23857 22729 23891 22763
rect 23891 22729 23900 22763
rect 23848 22720 23900 22729
rect 24584 22720 24636 22772
rect 26240 22720 26292 22772
rect 26424 22720 26476 22772
rect 27068 22720 27120 22772
rect 29368 22720 29420 22772
rect 31024 22720 31076 22772
rect 34704 22720 34756 22772
rect 29000 22652 29052 22704
rect 23296 22584 23348 22636
rect 24308 22627 24360 22636
rect 22376 22516 22428 22568
rect 17960 22380 18012 22432
rect 23572 22380 23624 22432
rect 24308 22593 24317 22627
rect 24317 22593 24351 22627
rect 24351 22593 24360 22627
rect 24308 22584 24360 22593
rect 27436 22627 27488 22636
rect 27436 22593 27445 22627
rect 27445 22593 27479 22627
rect 27479 22593 27488 22627
rect 27436 22584 27488 22593
rect 27712 22627 27764 22636
rect 27712 22593 27721 22627
rect 27721 22593 27755 22627
rect 27755 22593 27764 22627
rect 27712 22584 27764 22593
rect 27988 22627 28040 22636
rect 27988 22593 27997 22627
rect 27997 22593 28031 22627
rect 28031 22593 28040 22627
rect 27988 22584 28040 22593
rect 28356 22627 28408 22636
rect 28356 22593 28365 22627
rect 28365 22593 28399 22627
rect 28399 22593 28408 22627
rect 28356 22584 28408 22593
rect 28540 22584 28592 22636
rect 29644 22584 29696 22636
rect 30380 22584 30432 22636
rect 30840 22584 30892 22636
rect 34060 22584 34112 22636
rect 35624 22720 35676 22772
rect 35716 22720 35768 22772
rect 35900 22720 35952 22772
rect 36268 22763 36320 22772
rect 36268 22729 36277 22763
rect 36277 22729 36311 22763
rect 36311 22729 36320 22763
rect 36268 22720 36320 22729
rect 36636 22720 36688 22772
rect 36728 22720 36780 22772
rect 37832 22763 37884 22772
rect 37832 22729 37841 22763
rect 37841 22729 37875 22763
rect 37875 22729 37884 22763
rect 37832 22720 37884 22729
rect 40316 22763 40368 22772
rect 40316 22729 40325 22763
rect 40325 22729 40359 22763
rect 40359 22729 40368 22763
rect 40316 22720 40368 22729
rect 43260 22720 43312 22772
rect 44732 22720 44784 22772
rect 45560 22720 45612 22772
rect 45836 22763 45888 22772
rect 45836 22729 45845 22763
rect 45845 22729 45879 22763
rect 45879 22729 45888 22763
rect 45836 22720 45888 22729
rect 49148 22763 49200 22772
rect 49148 22729 49157 22763
rect 49157 22729 49191 22763
rect 49191 22729 49200 22763
rect 49148 22720 49200 22729
rect 33600 22516 33652 22568
rect 35624 22584 35676 22636
rect 36084 22584 36136 22636
rect 36268 22584 36320 22636
rect 37556 22652 37608 22704
rect 38936 22652 38988 22704
rect 40408 22652 40460 22704
rect 40592 22652 40644 22704
rect 48136 22652 48188 22704
rect 27252 22448 27304 22500
rect 30380 22448 30432 22500
rect 30472 22448 30524 22500
rect 33140 22448 33192 22500
rect 36912 22627 36964 22636
rect 36912 22593 36921 22627
rect 36921 22593 36955 22627
rect 36955 22593 36964 22627
rect 37464 22627 37516 22636
rect 36912 22584 36964 22593
rect 37464 22593 37473 22627
rect 37473 22593 37507 22627
rect 37507 22593 37516 22627
rect 37464 22584 37516 22593
rect 39028 22584 39080 22636
rect 43812 22627 43864 22636
rect 43812 22593 43821 22627
rect 43821 22593 43855 22627
rect 43855 22593 43864 22627
rect 43812 22584 43864 22593
rect 37188 22516 37240 22568
rect 38936 22559 38988 22568
rect 38936 22525 38945 22559
rect 38945 22525 38979 22559
rect 38979 22525 38988 22559
rect 38936 22516 38988 22525
rect 43168 22516 43220 22568
rect 44548 22584 44600 22636
rect 44732 22627 44784 22636
rect 44732 22593 44766 22627
rect 44766 22593 44784 22627
rect 44732 22584 44784 22593
rect 48872 22584 48924 22636
rect 56508 22627 56560 22636
rect 56508 22593 56517 22627
rect 56517 22593 56551 22627
rect 56551 22593 56560 22627
rect 56508 22584 56560 22593
rect 56784 22584 56836 22636
rect 58072 22627 58124 22636
rect 58072 22593 58081 22627
rect 58081 22593 58115 22627
rect 58115 22593 58124 22627
rect 58072 22584 58124 22593
rect 34612 22380 34664 22432
rect 35900 22380 35952 22432
rect 36176 22380 36228 22432
rect 36452 22380 36504 22432
rect 43720 22448 43772 22500
rect 44272 22380 44324 22432
rect 56416 22448 56468 22500
rect 48136 22380 48188 22432
rect 56324 22380 56376 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 13544 22219 13596 22228
rect 13544 22185 13553 22219
rect 13553 22185 13587 22219
rect 13587 22185 13596 22219
rect 13544 22176 13596 22185
rect 14280 22176 14332 22228
rect 16856 22176 16908 22228
rect 53380 22176 53432 22228
rect 26976 22108 27028 22160
rect 27988 22108 28040 22160
rect 13360 22015 13412 22024
rect 13360 21981 13369 22015
rect 13369 21981 13403 22015
rect 13403 21981 13412 22015
rect 13360 21972 13412 21981
rect 14372 22015 14424 22024
rect 14372 21981 14381 22015
rect 14381 21981 14415 22015
rect 14415 21981 14424 22015
rect 14372 21972 14424 21981
rect 16672 21972 16724 22024
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 24400 22040 24452 22092
rect 29736 22040 29788 22092
rect 31484 22108 31536 22160
rect 33140 22108 33192 22160
rect 34152 22151 34204 22160
rect 34152 22117 34161 22151
rect 34161 22117 34195 22151
rect 34195 22117 34204 22151
rect 34152 22108 34204 22117
rect 37096 22151 37148 22160
rect 37096 22117 37105 22151
rect 37105 22117 37139 22151
rect 37139 22117 37148 22151
rect 37096 22108 37148 22117
rect 40040 22108 40092 22160
rect 22284 21972 22336 22024
rect 22376 21972 22428 22024
rect 25136 21972 25188 22024
rect 20720 21904 20772 21956
rect 26516 21904 26568 21956
rect 26884 22015 26936 22024
rect 26884 21981 26893 22015
rect 26893 21981 26927 22015
rect 26927 21981 26936 22015
rect 26884 21972 26936 21981
rect 29276 21972 29328 22024
rect 30012 21972 30064 22024
rect 30656 22040 30708 22092
rect 31116 22040 31168 22092
rect 30932 21972 30984 22024
rect 31576 21972 31628 22024
rect 36544 22040 36596 22092
rect 37188 22040 37240 22092
rect 39120 22083 39172 22092
rect 33968 22015 34020 22024
rect 33968 21981 34000 22015
rect 34000 21981 34020 22015
rect 33968 21972 34020 21981
rect 35440 21972 35492 22024
rect 35624 21972 35676 22024
rect 39120 22049 39129 22083
rect 39129 22049 39163 22083
rect 39163 22049 39172 22083
rect 39120 22040 39172 22049
rect 45376 22108 45428 22160
rect 15936 21836 15988 21888
rect 16212 21836 16264 21888
rect 16580 21836 16632 21888
rect 22008 21836 22060 21888
rect 22928 21879 22980 21888
rect 22928 21845 22937 21879
rect 22937 21845 22971 21879
rect 22971 21845 22980 21879
rect 22928 21836 22980 21845
rect 27252 21836 27304 21888
rect 31760 21904 31812 21956
rect 34152 21904 34204 21956
rect 36544 21904 36596 21956
rect 37464 21972 37516 22024
rect 38108 22015 38160 22024
rect 38108 21981 38117 22015
rect 38117 21981 38151 22015
rect 38151 21981 38160 22015
rect 38108 21972 38160 21981
rect 38844 22015 38896 22024
rect 38844 21981 38853 22015
rect 38853 21981 38887 22015
rect 38887 21981 38896 22015
rect 38844 21972 38896 21981
rect 39672 21972 39724 22024
rect 40040 22015 40092 22024
rect 40040 21981 40049 22015
rect 40049 21981 40083 22015
rect 40083 21981 40092 22015
rect 40316 22015 40368 22024
rect 40040 21972 40092 21981
rect 40316 21981 40325 22015
rect 40325 21981 40359 22015
rect 40359 21981 40368 22015
rect 40316 21972 40368 21981
rect 40592 21972 40644 22024
rect 43352 22015 43404 22024
rect 43352 21981 43361 22015
rect 43361 21981 43395 22015
rect 43395 21981 43404 22015
rect 43352 21972 43404 21981
rect 43996 22015 44048 22024
rect 43996 21981 44002 22015
rect 44002 21981 44036 22015
rect 44036 21981 44048 22015
rect 43996 21972 44048 21981
rect 44364 21972 44416 22024
rect 37280 21947 37332 21956
rect 37280 21913 37289 21947
rect 37289 21913 37323 21947
rect 37323 21913 37332 21947
rect 37280 21904 37332 21913
rect 39488 21904 39540 21956
rect 43260 21947 43312 21956
rect 43260 21913 43269 21947
rect 43269 21913 43303 21947
rect 43303 21913 43312 21947
rect 43260 21904 43312 21913
rect 45560 21972 45612 22024
rect 47492 22015 47544 22024
rect 47492 21981 47501 22015
rect 47501 21981 47535 22015
rect 47535 21981 47544 22015
rect 47492 21972 47544 21981
rect 47860 22015 47912 22024
rect 47860 21981 47869 22015
rect 47869 21981 47903 22015
rect 47903 21981 47912 22015
rect 47860 21972 47912 21981
rect 49148 22108 49200 22160
rect 48872 22083 48924 22092
rect 48872 22049 48881 22083
rect 48881 22049 48915 22083
rect 48915 22049 48924 22083
rect 48872 22040 48924 22049
rect 51632 22040 51684 22092
rect 53932 22040 53984 22092
rect 48504 22015 48556 22024
rect 48504 21981 48513 22015
rect 48513 21981 48547 22015
rect 48547 21981 48556 22015
rect 48504 21972 48556 21981
rect 29828 21879 29880 21888
rect 29828 21845 29837 21879
rect 29837 21845 29871 21879
rect 29871 21845 29880 21879
rect 29828 21836 29880 21845
rect 30196 21836 30248 21888
rect 33876 21836 33928 21888
rect 34336 21836 34388 21888
rect 43812 21879 43864 21888
rect 43812 21845 43821 21879
rect 43821 21845 43855 21879
rect 43855 21845 43864 21879
rect 43812 21836 43864 21845
rect 43904 21836 43956 21888
rect 47860 21836 47912 21888
rect 51724 21972 51776 22024
rect 58164 21947 58216 21956
rect 58164 21913 58173 21947
rect 58173 21913 58207 21947
rect 58207 21913 58216 21947
rect 58164 21904 58216 21913
rect 48780 21836 48832 21888
rect 57888 21836 57940 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 13360 21632 13412 21684
rect 15568 21632 15620 21684
rect 7656 21564 7708 21616
rect 13728 21564 13780 21616
rect 15936 21564 15988 21616
rect 15200 21496 15252 21548
rect 15660 21539 15712 21548
rect 1860 21471 1912 21480
rect 1860 21437 1869 21471
rect 1869 21437 1903 21471
rect 1903 21437 1912 21471
rect 1860 21428 1912 21437
rect 15660 21505 15669 21539
rect 15669 21505 15703 21539
rect 15703 21505 15712 21539
rect 15660 21496 15712 21505
rect 20444 21632 20496 21684
rect 21180 21632 21232 21684
rect 27160 21675 27212 21684
rect 27160 21641 27169 21675
rect 27169 21641 27203 21675
rect 27203 21641 27212 21675
rect 27160 21632 27212 21641
rect 27436 21632 27488 21684
rect 30656 21632 30708 21684
rect 34612 21632 34664 21684
rect 35440 21675 35492 21684
rect 16212 21564 16264 21616
rect 19432 21564 19484 21616
rect 22928 21564 22980 21616
rect 29736 21564 29788 21616
rect 29828 21564 29880 21616
rect 33416 21564 33468 21616
rect 35440 21641 35449 21675
rect 35449 21641 35483 21675
rect 35483 21641 35492 21675
rect 35440 21632 35492 21641
rect 35716 21632 35768 21684
rect 16028 21428 16080 21480
rect 17960 21496 18012 21548
rect 19156 21539 19208 21548
rect 19156 21505 19165 21539
rect 19165 21505 19199 21539
rect 19199 21505 19208 21539
rect 19156 21496 19208 21505
rect 22376 21539 22428 21548
rect 22376 21505 22385 21539
rect 22385 21505 22419 21539
rect 22419 21505 22428 21539
rect 22376 21496 22428 21505
rect 24308 21539 24360 21548
rect 24308 21505 24317 21539
rect 24317 21505 24351 21539
rect 24351 21505 24360 21539
rect 27344 21539 27396 21548
rect 24308 21496 24360 21505
rect 27344 21505 27350 21539
rect 27350 21505 27384 21539
rect 27384 21505 27396 21539
rect 27344 21496 27396 21505
rect 27620 21496 27672 21548
rect 30196 21496 30248 21548
rect 31392 21539 31444 21548
rect 31392 21505 31401 21539
rect 31401 21505 31435 21539
rect 31435 21505 31444 21539
rect 31392 21496 31444 21505
rect 31576 21539 31628 21548
rect 31576 21505 31585 21539
rect 31585 21505 31619 21539
rect 31619 21505 31628 21539
rect 31576 21496 31628 21505
rect 24400 21428 24452 21480
rect 26148 21428 26200 21480
rect 16948 21360 17000 21412
rect 19156 21360 19208 21412
rect 19340 21360 19392 21412
rect 18604 21335 18656 21344
rect 18604 21301 18613 21335
rect 18613 21301 18647 21335
rect 18647 21301 18656 21335
rect 18604 21292 18656 21301
rect 20904 21292 20956 21344
rect 21272 21292 21324 21344
rect 28908 21428 28960 21480
rect 30380 21360 30432 21412
rect 31300 21360 31352 21412
rect 31576 21360 31628 21412
rect 26700 21292 26752 21344
rect 27712 21335 27764 21344
rect 27712 21301 27721 21335
rect 27721 21301 27755 21335
rect 27755 21301 27764 21335
rect 27712 21292 27764 21301
rect 27804 21292 27856 21344
rect 34336 21496 34388 21548
rect 35440 21496 35492 21548
rect 35716 21539 35768 21548
rect 35716 21505 35725 21539
rect 35725 21505 35759 21539
rect 35759 21505 35768 21539
rect 35716 21496 35768 21505
rect 36452 21632 36504 21684
rect 37004 21564 37056 21616
rect 36084 21539 36136 21548
rect 36084 21505 36093 21539
rect 36093 21505 36127 21539
rect 36127 21505 36136 21539
rect 36084 21496 36136 21505
rect 36268 21496 36320 21548
rect 37372 21496 37424 21548
rect 33968 21428 34020 21480
rect 36912 21428 36964 21480
rect 37648 21428 37700 21480
rect 38844 21564 38896 21616
rect 47860 21632 47912 21684
rect 51632 21632 51684 21684
rect 40408 21539 40460 21548
rect 40408 21505 40417 21539
rect 40417 21505 40451 21539
rect 40451 21505 40460 21539
rect 40408 21496 40460 21505
rect 40500 21496 40552 21548
rect 44272 21539 44324 21548
rect 44272 21505 44306 21539
rect 44306 21505 44324 21539
rect 58808 21564 58860 21616
rect 44272 21496 44324 21505
rect 48504 21496 48556 21548
rect 43352 21428 43404 21480
rect 50160 21496 50212 21548
rect 56232 21496 56284 21548
rect 56784 21496 56836 21548
rect 57152 21539 57204 21548
rect 57152 21505 57161 21539
rect 57161 21505 57195 21539
rect 57195 21505 57204 21539
rect 57152 21496 57204 21505
rect 52000 21428 52052 21480
rect 37004 21292 37056 21344
rect 37464 21335 37516 21344
rect 37464 21301 37473 21335
rect 37473 21301 37507 21335
rect 37507 21301 37516 21335
rect 37464 21292 37516 21301
rect 38292 21360 38344 21412
rect 41788 21335 41840 21344
rect 41788 21301 41797 21335
rect 41797 21301 41831 21335
rect 41831 21301 41840 21335
rect 41788 21292 41840 21301
rect 55956 21360 56008 21412
rect 45376 21335 45428 21344
rect 45376 21301 45385 21335
rect 45385 21301 45419 21335
rect 45419 21301 45428 21335
rect 45376 21292 45428 21301
rect 48780 21292 48832 21344
rect 50436 21335 50488 21344
rect 50436 21301 50445 21335
rect 50445 21301 50479 21335
rect 50479 21301 50488 21335
rect 50436 21292 50488 21301
rect 56968 21292 57020 21344
rect 57244 21335 57296 21344
rect 57244 21301 57253 21335
rect 57253 21301 57287 21335
rect 57287 21301 57296 21335
rect 57244 21292 57296 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 17776 21131 17828 21140
rect 17776 21097 17785 21131
rect 17785 21097 17819 21131
rect 17819 21097 17828 21131
rect 17776 21088 17828 21097
rect 18604 21088 18656 21140
rect 29368 21088 29420 21140
rect 29460 21088 29512 21140
rect 29920 21088 29972 21140
rect 31024 21088 31076 21140
rect 31300 21088 31352 21140
rect 31392 21088 31444 21140
rect 31760 21088 31812 21140
rect 36268 21088 36320 21140
rect 36360 21088 36412 21140
rect 44456 21088 44508 21140
rect 51724 21131 51776 21140
rect 51724 21097 51733 21131
rect 51733 21097 51767 21131
rect 51767 21097 51776 21131
rect 51724 21088 51776 21097
rect 57796 21088 57848 21140
rect 19340 21020 19392 21072
rect 24308 21020 24360 21072
rect 15936 20952 15988 21004
rect 27252 21020 27304 21072
rect 27804 21020 27856 21072
rect 35808 21020 35860 21072
rect 37464 21020 37516 21072
rect 47492 21020 47544 21072
rect 10784 20884 10836 20936
rect 15200 20884 15252 20936
rect 16580 20927 16632 20936
rect 16580 20893 16589 20927
rect 16589 20893 16623 20927
rect 16623 20893 16632 20927
rect 16580 20884 16632 20893
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 21732 20927 21784 20936
rect 1860 20859 1912 20868
rect 1860 20825 1869 20859
rect 1869 20825 1903 20859
rect 1903 20825 1912 20859
rect 1860 20816 1912 20825
rect 13728 20748 13780 20800
rect 18144 20816 18196 20868
rect 18420 20816 18472 20868
rect 21732 20893 21741 20927
rect 21741 20893 21775 20927
rect 21775 20893 21784 20927
rect 21732 20884 21784 20893
rect 22652 20884 22704 20936
rect 24860 20884 24912 20936
rect 32312 20952 32364 21004
rect 35440 20952 35492 21004
rect 36084 20952 36136 21004
rect 26148 20884 26200 20936
rect 28356 20884 28408 20936
rect 28540 20927 28592 20936
rect 28540 20893 28549 20927
rect 28549 20893 28583 20927
rect 28583 20893 28592 20927
rect 28540 20884 28592 20893
rect 28816 20927 28868 20936
rect 28816 20893 28825 20927
rect 28825 20893 28859 20927
rect 28859 20893 28868 20927
rect 28816 20884 28868 20893
rect 30380 20927 30432 20936
rect 20996 20816 21048 20868
rect 17040 20748 17092 20800
rect 30380 20893 30389 20927
rect 30389 20893 30423 20927
rect 30423 20893 30432 20927
rect 30380 20884 30432 20893
rect 35348 20884 35400 20936
rect 36268 20884 36320 20936
rect 36452 20884 36504 20936
rect 36912 20927 36964 20936
rect 36912 20893 36921 20927
rect 36921 20893 36955 20927
rect 36955 20893 36964 20927
rect 36912 20884 36964 20893
rect 30472 20816 30524 20868
rect 22928 20791 22980 20800
rect 22928 20757 22937 20791
rect 22937 20757 22971 20791
rect 22971 20757 22980 20791
rect 22928 20748 22980 20757
rect 25320 20748 25372 20800
rect 26700 20748 26752 20800
rect 27344 20748 27396 20800
rect 27712 20748 27764 20800
rect 28448 20748 28500 20800
rect 33968 20816 34020 20868
rect 35440 20859 35492 20868
rect 32680 20748 32732 20800
rect 35440 20825 35449 20859
rect 35449 20825 35483 20859
rect 35483 20825 35492 20859
rect 35440 20816 35492 20825
rect 35624 20816 35676 20868
rect 36268 20791 36320 20800
rect 36268 20757 36277 20791
rect 36277 20757 36311 20791
rect 36311 20757 36320 20791
rect 36268 20748 36320 20757
rect 37004 20816 37056 20868
rect 40224 20952 40276 21004
rect 38200 20927 38252 20936
rect 38200 20893 38209 20927
rect 38209 20893 38243 20927
rect 38243 20893 38252 20927
rect 38200 20884 38252 20893
rect 41788 20952 41840 21004
rect 43352 20995 43404 21004
rect 43352 20961 43361 20995
rect 43361 20961 43395 20995
rect 43395 20961 43404 20995
rect 43352 20952 43404 20961
rect 43444 20952 43496 21004
rect 44640 20952 44692 21004
rect 48228 20952 48280 21004
rect 56232 20995 56284 21004
rect 56232 20961 56241 20995
rect 56241 20961 56275 20995
rect 56275 20961 56284 20995
rect 56232 20952 56284 20961
rect 56876 20995 56928 21004
rect 56876 20961 56885 20995
rect 56885 20961 56919 20995
rect 56919 20961 56928 20995
rect 56876 20952 56928 20961
rect 41328 20884 41380 20936
rect 42800 20884 42852 20936
rect 48136 20884 48188 20936
rect 52368 20884 52420 20936
rect 56048 20884 56100 20936
rect 37556 20859 37608 20868
rect 37556 20825 37565 20859
rect 37565 20825 37599 20859
rect 37599 20825 37608 20859
rect 37556 20816 37608 20825
rect 37648 20816 37700 20868
rect 40684 20816 40736 20868
rect 46848 20859 46900 20868
rect 46848 20825 46857 20859
rect 46857 20825 46891 20859
rect 46891 20825 46900 20859
rect 46848 20816 46900 20825
rect 50436 20816 50488 20868
rect 37924 20748 37976 20800
rect 38384 20791 38436 20800
rect 38384 20757 38393 20791
rect 38393 20757 38427 20791
rect 38427 20757 38436 20791
rect 38384 20748 38436 20757
rect 40316 20748 40368 20800
rect 40592 20791 40644 20800
rect 40592 20757 40601 20791
rect 40601 20757 40635 20791
rect 40635 20757 40644 20791
rect 40592 20748 40644 20757
rect 45560 20748 45612 20800
rect 46112 20748 46164 20800
rect 48320 20748 48372 20800
rect 56140 20859 56192 20868
rect 56140 20825 56149 20859
rect 56149 20825 56183 20859
rect 56183 20825 56192 20859
rect 56140 20816 56192 20825
rect 56968 20884 57020 20936
rect 53932 20748 53984 20800
rect 56416 20816 56468 20868
rect 57704 20748 57756 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 16672 20544 16724 20596
rect 15660 20476 15712 20528
rect 15108 20408 15160 20460
rect 18236 20476 18288 20528
rect 1768 20383 1820 20392
rect 1768 20349 1777 20383
rect 1777 20349 1811 20383
rect 1811 20349 1820 20383
rect 1768 20340 1820 20349
rect 16028 20383 16080 20392
rect 16028 20349 16037 20383
rect 16037 20349 16071 20383
rect 16071 20349 16080 20383
rect 16028 20340 16080 20349
rect 16948 20383 17000 20392
rect 16948 20349 16957 20383
rect 16957 20349 16991 20383
rect 16991 20349 17000 20383
rect 16948 20340 17000 20349
rect 17868 20408 17920 20460
rect 20812 20476 20864 20528
rect 22928 20476 22980 20528
rect 24860 20544 24912 20596
rect 27344 20544 27396 20596
rect 27712 20544 27764 20596
rect 26976 20476 27028 20528
rect 27252 20476 27304 20528
rect 27436 20519 27488 20528
rect 27436 20485 27445 20519
rect 27445 20485 27479 20519
rect 27479 20485 27488 20519
rect 27436 20476 27488 20485
rect 28540 20476 28592 20528
rect 37648 20544 37700 20596
rect 38844 20544 38896 20596
rect 30380 20476 30432 20528
rect 30840 20476 30892 20528
rect 18420 20451 18472 20460
rect 18420 20417 18429 20451
rect 18429 20417 18463 20451
rect 18463 20417 18472 20451
rect 19156 20451 19208 20460
rect 18420 20408 18472 20417
rect 19156 20417 19165 20451
rect 19165 20417 19199 20451
rect 19199 20417 19208 20451
rect 19156 20408 19208 20417
rect 22376 20451 22428 20460
rect 22376 20417 22385 20451
rect 22385 20417 22419 20451
rect 22419 20417 22428 20451
rect 22376 20408 22428 20417
rect 27344 20451 27396 20460
rect 17868 20272 17920 20324
rect 18236 20272 18288 20324
rect 18604 20383 18656 20392
rect 18604 20349 18613 20383
rect 18613 20349 18647 20383
rect 18647 20349 18656 20383
rect 20720 20383 20772 20392
rect 18604 20340 18656 20349
rect 20720 20349 20729 20383
rect 20729 20349 20763 20383
rect 20763 20349 20772 20383
rect 20720 20340 20772 20349
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 27528 20451 27580 20460
rect 27528 20417 27537 20451
rect 27537 20417 27571 20451
rect 27571 20417 27580 20451
rect 27528 20408 27580 20417
rect 29460 20408 29512 20460
rect 28816 20340 28868 20392
rect 31576 20408 31628 20460
rect 32496 20476 32548 20528
rect 32680 20476 32732 20528
rect 33324 20476 33376 20528
rect 36912 20476 36964 20528
rect 15936 20204 15988 20256
rect 19156 20204 19208 20256
rect 27620 20272 27672 20324
rect 27712 20315 27764 20324
rect 27712 20281 27721 20315
rect 27721 20281 27755 20315
rect 27755 20281 27764 20315
rect 27712 20272 27764 20281
rect 28632 20272 28684 20324
rect 30840 20340 30892 20392
rect 33968 20340 34020 20392
rect 36544 20340 36596 20392
rect 37188 20340 37240 20392
rect 37464 20451 37516 20460
rect 37464 20417 37473 20451
rect 37473 20417 37507 20451
rect 37507 20417 37516 20451
rect 37464 20408 37516 20417
rect 38384 20408 38436 20460
rect 39948 20476 40000 20528
rect 40500 20544 40552 20596
rect 48320 20544 48372 20596
rect 50160 20544 50212 20596
rect 54300 20544 54352 20596
rect 57612 20544 57664 20596
rect 38936 20408 38988 20460
rect 40316 20451 40368 20460
rect 40316 20417 40325 20451
rect 40325 20417 40359 20451
rect 40359 20417 40368 20451
rect 40316 20408 40368 20417
rect 43444 20408 43496 20460
rect 48044 20476 48096 20528
rect 48228 20476 48280 20528
rect 45560 20451 45612 20460
rect 45560 20417 45569 20451
rect 45569 20417 45603 20451
rect 45603 20417 45612 20451
rect 45560 20408 45612 20417
rect 45744 20451 45796 20460
rect 45744 20417 45753 20451
rect 45753 20417 45787 20451
rect 45787 20417 45796 20451
rect 45744 20408 45796 20417
rect 49700 20408 49752 20460
rect 49976 20451 50028 20460
rect 49976 20417 49985 20451
rect 49985 20417 50019 20451
rect 50019 20417 50028 20451
rect 49976 20408 50028 20417
rect 50712 20408 50764 20460
rect 30564 20272 30616 20324
rect 38844 20272 38896 20324
rect 24124 20204 24176 20256
rect 35900 20204 35952 20256
rect 36636 20204 36688 20256
rect 38016 20204 38068 20256
rect 38108 20204 38160 20256
rect 51724 20340 51776 20392
rect 52368 20408 52420 20460
rect 53196 20451 53248 20460
rect 53196 20417 53230 20451
rect 53230 20417 53248 20451
rect 53196 20408 53248 20417
rect 52552 20340 52604 20392
rect 52092 20272 52144 20324
rect 45836 20204 45888 20256
rect 51816 20204 51868 20256
rect 52368 20204 52420 20256
rect 54300 20247 54352 20256
rect 54300 20213 54309 20247
rect 54309 20213 54343 20247
rect 54343 20213 54352 20247
rect 54300 20204 54352 20213
rect 56784 20204 56836 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 15200 20000 15252 20052
rect 20996 20043 21048 20052
rect 20996 20009 21005 20043
rect 21005 20009 21039 20043
rect 21039 20009 21048 20043
rect 20996 20000 21048 20009
rect 22284 20000 22336 20052
rect 26516 20043 26568 20052
rect 26516 20009 26525 20043
rect 26525 20009 26559 20043
rect 26559 20009 26568 20043
rect 26516 20000 26568 20009
rect 28540 20043 28592 20052
rect 28540 20009 28549 20043
rect 28549 20009 28583 20043
rect 28583 20009 28592 20043
rect 28540 20000 28592 20009
rect 31852 20000 31904 20052
rect 32312 20000 32364 20052
rect 34152 20000 34204 20052
rect 39672 20000 39724 20052
rect 40224 20043 40276 20052
rect 40224 20009 40233 20043
rect 40233 20009 40267 20043
rect 40267 20009 40276 20043
rect 40224 20000 40276 20009
rect 41236 20000 41288 20052
rect 58624 20000 58676 20052
rect 17776 19932 17828 19984
rect 20260 19932 20312 19984
rect 27344 19932 27396 19984
rect 27896 19932 27948 19984
rect 1492 19796 1544 19848
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 20444 19864 20496 19916
rect 22376 19864 22428 19916
rect 1860 19771 1912 19780
rect 1860 19737 1869 19771
rect 1869 19737 1903 19771
rect 1903 19737 1912 19771
rect 1860 19728 1912 19737
rect 17868 19728 17920 19780
rect 18420 19728 18472 19780
rect 18972 19796 19024 19848
rect 27712 19864 27764 19916
rect 29460 19864 29512 19916
rect 30472 19907 30524 19916
rect 30472 19873 30481 19907
rect 30481 19873 30515 19907
rect 30515 19873 30524 19907
rect 30472 19864 30524 19873
rect 24676 19839 24728 19848
rect 24676 19805 24685 19839
rect 24685 19805 24719 19839
rect 24719 19805 24728 19839
rect 24676 19796 24728 19805
rect 24768 19796 24820 19848
rect 25320 19839 25372 19848
rect 25320 19805 25329 19839
rect 25329 19805 25363 19839
rect 25363 19805 25372 19839
rect 25320 19796 25372 19805
rect 28448 19796 28500 19848
rect 28816 19796 28868 19848
rect 21272 19728 21324 19780
rect 21824 19728 21876 19780
rect 22652 19728 22704 19780
rect 25504 19728 25556 19780
rect 29736 19771 29788 19780
rect 19340 19660 19392 19712
rect 28724 19703 28776 19712
rect 28724 19669 28733 19703
rect 28733 19669 28767 19703
rect 28767 19669 28776 19703
rect 28724 19660 28776 19669
rect 29736 19737 29745 19771
rect 29745 19737 29779 19771
rect 29779 19737 29788 19771
rect 29736 19728 29788 19737
rect 29828 19660 29880 19712
rect 30748 19839 30800 19848
rect 30748 19805 30757 19839
rect 30757 19805 30791 19839
rect 30791 19805 30800 19839
rect 30748 19796 30800 19805
rect 31116 19796 31168 19848
rect 34888 19839 34940 19848
rect 34888 19805 34897 19839
rect 34897 19805 34931 19839
rect 34931 19805 34940 19839
rect 37556 19864 37608 19916
rect 34888 19796 34940 19805
rect 37280 19796 37332 19848
rect 37648 19839 37700 19848
rect 37648 19805 37657 19839
rect 37657 19805 37691 19839
rect 37691 19805 37700 19839
rect 37648 19796 37700 19805
rect 37740 19796 37792 19848
rect 38016 19796 38068 19848
rect 41328 19864 41380 19916
rect 41880 19864 41932 19916
rect 45928 19907 45980 19916
rect 45928 19873 45937 19907
rect 45937 19873 45971 19907
rect 45971 19873 45980 19907
rect 45928 19864 45980 19873
rect 46388 19932 46440 19984
rect 39672 19796 39724 19848
rect 40592 19796 40644 19848
rect 41052 19839 41104 19848
rect 41052 19805 41061 19839
rect 41061 19805 41095 19839
rect 41095 19805 41104 19839
rect 41052 19796 41104 19805
rect 41236 19839 41288 19848
rect 41236 19805 41245 19839
rect 41245 19805 41279 19839
rect 41279 19805 41288 19839
rect 41236 19796 41288 19805
rect 45836 19839 45888 19848
rect 45836 19805 45845 19839
rect 45845 19805 45879 19839
rect 45879 19805 45888 19839
rect 45836 19796 45888 19805
rect 46204 19839 46256 19848
rect 46204 19805 46213 19839
rect 46213 19805 46247 19839
rect 46247 19805 46256 19839
rect 46204 19796 46256 19805
rect 31392 19728 31444 19780
rect 45100 19728 45152 19780
rect 45376 19728 45428 19780
rect 49976 19796 50028 19848
rect 54300 19864 54352 19916
rect 58164 19907 58216 19916
rect 58164 19873 58173 19907
rect 58173 19873 58207 19907
rect 58207 19873 58216 19907
rect 58164 19864 58216 19873
rect 47124 19728 47176 19780
rect 52368 19771 52420 19780
rect 52368 19737 52377 19771
rect 52377 19737 52411 19771
rect 52411 19737 52420 19771
rect 52368 19728 52420 19737
rect 52552 19728 52604 19780
rect 56324 19728 56376 19780
rect 56508 19728 56560 19780
rect 57060 19771 57112 19780
rect 57060 19737 57069 19771
rect 57069 19737 57103 19771
rect 57103 19737 57112 19771
rect 57060 19728 57112 19737
rect 30656 19660 30708 19712
rect 31116 19660 31168 19712
rect 33784 19660 33836 19712
rect 34336 19660 34388 19712
rect 46388 19660 46440 19712
rect 52184 19660 52236 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 15108 19499 15160 19508
rect 15108 19465 15117 19499
rect 15117 19465 15151 19499
rect 15151 19465 15160 19499
rect 15108 19456 15160 19465
rect 18328 19499 18380 19508
rect 18328 19465 18337 19499
rect 18337 19465 18371 19499
rect 18371 19465 18380 19499
rect 18328 19456 18380 19465
rect 19156 19456 19208 19508
rect 25504 19499 25556 19508
rect 25504 19465 25513 19499
rect 25513 19465 25547 19499
rect 25547 19465 25556 19499
rect 25504 19456 25556 19465
rect 17776 19388 17828 19440
rect 18604 19388 18656 19440
rect 14924 19252 14976 19304
rect 17592 19363 17644 19372
rect 17592 19329 17601 19363
rect 17601 19329 17635 19363
rect 17635 19329 17644 19363
rect 17592 19320 17644 19329
rect 18236 19363 18288 19372
rect 18236 19329 18245 19363
rect 18245 19329 18279 19363
rect 18279 19329 18288 19363
rect 18236 19320 18288 19329
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 14740 19184 14792 19236
rect 16396 19252 16448 19304
rect 18972 19252 19024 19304
rect 24124 19320 24176 19372
rect 24308 19363 24360 19372
rect 24308 19329 24317 19363
rect 24317 19329 24351 19363
rect 24351 19329 24360 19363
rect 24308 19320 24360 19329
rect 27528 19456 27580 19508
rect 28540 19456 28592 19508
rect 34704 19456 34756 19508
rect 37740 19456 37792 19508
rect 40040 19456 40092 19508
rect 45376 19499 45428 19508
rect 27344 19363 27396 19372
rect 22100 19252 22152 19304
rect 22376 19252 22428 19304
rect 22468 19295 22520 19304
rect 22468 19261 22477 19295
rect 22477 19261 22511 19295
rect 22511 19261 22520 19295
rect 22468 19252 22520 19261
rect 21180 19184 21232 19236
rect 21272 19184 21324 19236
rect 27344 19329 27354 19363
rect 27354 19329 27388 19363
rect 27388 19329 27396 19363
rect 27344 19320 27396 19329
rect 28264 19320 28316 19372
rect 28540 19363 28592 19372
rect 28540 19329 28549 19363
rect 28549 19329 28583 19363
rect 28583 19329 28592 19363
rect 28540 19320 28592 19329
rect 27436 19295 27488 19304
rect 27436 19261 27445 19295
rect 27445 19261 27479 19295
rect 27479 19261 27488 19295
rect 27436 19252 27488 19261
rect 27620 19295 27672 19304
rect 27620 19261 27629 19295
rect 27629 19261 27663 19295
rect 27663 19261 27672 19295
rect 27620 19252 27672 19261
rect 18604 19159 18656 19168
rect 18604 19125 18613 19159
rect 18613 19125 18647 19159
rect 18647 19125 18656 19159
rect 18604 19116 18656 19125
rect 21364 19159 21416 19168
rect 21364 19125 21373 19159
rect 21373 19125 21407 19159
rect 21407 19125 21416 19159
rect 21364 19116 21416 19125
rect 23388 19116 23440 19168
rect 27160 19159 27212 19168
rect 27160 19125 27169 19159
rect 27169 19125 27203 19159
rect 27203 19125 27212 19159
rect 27160 19116 27212 19125
rect 27896 19184 27948 19236
rect 28632 19184 28684 19236
rect 29000 19320 29052 19372
rect 29460 19363 29512 19372
rect 29460 19329 29469 19363
rect 29469 19329 29503 19363
rect 29503 19329 29512 19363
rect 29460 19320 29512 19329
rect 29828 19320 29880 19372
rect 37372 19388 37424 19440
rect 37556 19388 37608 19440
rect 37648 19388 37700 19440
rect 32588 19320 32640 19372
rect 34704 19320 34756 19372
rect 34796 19320 34848 19372
rect 35348 19363 35400 19372
rect 35348 19329 35382 19363
rect 35382 19329 35400 19363
rect 37740 19363 37792 19372
rect 35348 19320 35400 19329
rect 37740 19329 37749 19363
rect 37749 19329 37783 19363
rect 37783 19329 37792 19363
rect 37740 19320 37792 19329
rect 30656 19295 30708 19304
rect 30656 19261 30665 19295
rect 30665 19261 30699 19295
rect 30699 19261 30708 19295
rect 30656 19252 30708 19261
rect 31300 19252 31352 19304
rect 36084 19252 36136 19304
rect 37924 19363 37976 19372
rect 37924 19329 37933 19363
rect 37933 19329 37967 19363
rect 37967 19329 37976 19363
rect 37924 19320 37976 19329
rect 38660 19320 38712 19372
rect 38016 19252 38068 19304
rect 38384 19252 38436 19304
rect 42616 19320 42668 19372
rect 43352 19320 43404 19372
rect 44272 19363 44324 19372
rect 44272 19329 44306 19363
rect 44306 19329 44324 19363
rect 45376 19465 45385 19499
rect 45385 19465 45419 19499
rect 45419 19465 45428 19499
rect 45376 19456 45428 19465
rect 46204 19456 46256 19508
rect 45100 19388 45152 19440
rect 47124 19388 47176 19440
rect 44272 19320 44324 19329
rect 49976 19320 50028 19372
rect 52184 19363 52236 19372
rect 52184 19329 52193 19363
rect 52193 19329 52227 19363
rect 52227 19329 52236 19363
rect 52184 19320 52236 19329
rect 53196 19456 53248 19508
rect 58072 19456 58124 19508
rect 52460 19388 52512 19440
rect 53196 19320 53248 19372
rect 56784 19363 56836 19372
rect 56784 19329 56793 19363
rect 56793 19329 56827 19363
rect 56827 19329 56836 19363
rect 56784 19320 56836 19329
rect 52000 19295 52052 19304
rect 52000 19261 52009 19295
rect 52009 19261 52043 19295
rect 52043 19261 52052 19295
rect 52000 19252 52052 19261
rect 29092 19184 29144 19236
rect 31116 19184 31168 19236
rect 34888 19184 34940 19236
rect 30472 19116 30524 19168
rect 32772 19116 32824 19168
rect 33600 19116 33652 19168
rect 33784 19116 33836 19168
rect 36544 19116 36596 19168
rect 43444 19184 43496 19236
rect 46204 19184 46256 19236
rect 58992 19184 59044 19236
rect 39764 19116 39816 19168
rect 39948 19116 40000 19168
rect 44364 19116 44416 19168
rect 56968 19116 57020 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 10784 18955 10836 18964
rect 10784 18921 10793 18955
rect 10793 18921 10827 18955
rect 10827 18921 10836 18955
rect 10784 18912 10836 18921
rect 16212 18912 16264 18964
rect 17960 18912 18012 18964
rect 18328 18912 18380 18964
rect 17224 18844 17276 18896
rect 11152 18819 11204 18828
rect 11152 18785 11161 18819
rect 11161 18785 11195 18819
rect 11195 18785 11204 18819
rect 11152 18776 11204 18785
rect 14924 18776 14976 18828
rect 1952 18708 2004 18760
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 11244 18751 11296 18760
rect 11244 18717 11253 18751
rect 11253 18717 11287 18751
rect 11287 18717 11296 18751
rect 17684 18776 17736 18828
rect 11244 18708 11296 18717
rect 16212 18751 16264 18760
rect 16212 18717 16225 18751
rect 16225 18717 16264 18751
rect 16212 18708 16264 18717
rect 17132 18708 17184 18760
rect 15844 18640 15896 18692
rect 17500 18751 17552 18760
rect 17500 18717 17509 18751
rect 17509 18717 17543 18751
rect 17543 18717 17552 18751
rect 17500 18708 17552 18717
rect 18604 18819 18656 18828
rect 18604 18785 18613 18819
rect 18613 18785 18647 18819
rect 18647 18785 18656 18819
rect 18604 18776 18656 18785
rect 19432 18776 19484 18828
rect 19800 18819 19852 18828
rect 19800 18785 19809 18819
rect 19809 18785 19843 18819
rect 19843 18785 19852 18819
rect 19800 18776 19852 18785
rect 20904 18844 20956 18896
rect 25136 18912 25188 18964
rect 25688 18912 25740 18964
rect 28632 18912 28684 18964
rect 28816 18912 28868 18964
rect 34704 18912 34756 18964
rect 35348 18912 35400 18964
rect 22560 18844 22612 18896
rect 19432 18640 19484 18692
rect 20352 18640 20404 18692
rect 23664 18708 23716 18760
rect 27344 18776 27396 18828
rect 28080 18776 28132 18828
rect 27160 18708 27212 18760
rect 28540 18776 28592 18828
rect 30840 18844 30892 18896
rect 30472 18776 30524 18828
rect 27528 18640 27580 18692
rect 30380 18708 30432 18760
rect 30564 18751 30616 18760
rect 30564 18717 30573 18751
rect 30573 18717 30607 18751
rect 30607 18717 30616 18751
rect 30564 18708 30616 18717
rect 30748 18819 30800 18828
rect 30748 18785 30757 18819
rect 30757 18785 30791 18819
rect 30791 18785 30800 18819
rect 30748 18776 30800 18785
rect 31024 18708 31076 18760
rect 31576 18751 31628 18760
rect 31576 18717 31585 18751
rect 31585 18717 31619 18751
rect 31619 18717 31628 18751
rect 31576 18708 31628 18717
rect 33600 18844 33652 18896
rect 34888 18844 34940 18896
rect 35900 18912 35952 18964
rect 32772 18751 32824 18760
rect 30012 18640 30064 18692
rect 32220 18640 32272 18692
rect 32772 18717 32781 18751
rect 32781 18717 32815 18751
rect 32815 18717 32824 18751
rect 32772 18708 32824 18717
rect 32864 18751 32916 18760
rect 32864 18717 32873 18751
rect 32873 18717 32907 18751
rect 32907 18717 32916 18751
rect 33416 18751 33468 18760
rect 32864 18708 32916 18717
rect 33416 18717 33425 18751
rect 33425 18717 33459 18751
rect 33459 18717 33468 18751
rect 33416 18708 33468 18717
rect 33600 18751 33652 18760
rect 33600 18717 33609 18751
rect 33609 18717 33643 18751
rect 33643 18717 33652 18751
rect 33600 18708 33652 18717
rect 33876 18751 33928 18760
rect 33876 18717 33885 18751
rect 33885 18717 33919 18751
rect 33919 18717 33928 18751
rect 33876 18708 33928 18717
rect 35256 18708 35308 18760
rect 35348 18708 35400 18760
rect 36084 18844 36136 18896
rect 37464 18912 37516 18964
rect 37556 18912 37608 18964
rect 38384 18955 38436 18964
rect 38384 18921 38393 18955
rect 38393 18921 38427 18955
rect 38427 18921 38436 18955
rect 38384 18912 38436 18921
rect 37740 18844 37792 18896
rect 46204 18912 46256 18964
rect 57152 18912 57204 18964
rect 57888 18912 57940 18964
rect 38016 18776 38068 18828
rect 38752 18844 38804 18896
rect 33784 18640 33836 18692
rect 16856 18572 16908 18624
rect 17040 18615 17092 18624
rect 17040 18581 17049 18615
rect 17049 18581 17083 18615
rect 17083 18581 17092 18615
rect 17040 18572 17092 18581
rect 17224 18572 17276 18624
rect 21088 18572 21140 18624
rect 22560 18572 22612 18624
rect 22928 18615 22980 18624
rect 22928 18581 22937 18615
rect 22937 18581 22971 18615
rect 22971 18581 22980 18615
rect 22928 18572 22980 18581
rect 25320 18572 25372 18624
rect 25412 18572 25464 18624
rect 28080 18572 28132 18624
rect 28264 18572 28316 18624
rect 31300 18572 31352 18624
rect 31576 18572 31628 18624
rect 33692 18572 33744 18624
rect 36084 18751 36136 18760
rect 36084 18717 36093 18751
rect 36093 18717 36127 18751
rect 36127 18717 36136 18751
rect 36544 18751 36596 18760
rect 36084 18708 36136 18717
rect 36544 18717 36553 18751
rect 36553 18717 36587 18751
rect 36587 18717 36596 18751
rect 36544 18708 36596 18717
rect 37648 18708 37700 18760
rect 38568 18708 38620 18760
rect 41052 18776 41104 18828
rect 43996 18844 44048 18896
rect 44364 18887 44416 18896
rect 44364 18853 44373 18887
rect 44373 18853 44407 18887
rect 44407 18853 44416 18887
rect 44364 18844 44416 18853
rect 44272 18776 44324 18828
rect 36268 18640 36320 18692
rect 39028 18751 39080 18760
rect 39028 18717 39037 18751
rect 39037 18717 39071 18751
rect 39071 18717 39080 18751
rect 39028 18708 39080 18717
rect 43168 18751 43220 18760
rect 39212 18640 39264 18692
rect 43168 18717 43177 18751
rect 43177 18717 43211 18751
rect 43211 18717 43220 18751
rect 43168 18708 43220 18717
rect 45376 18776 45428 18828
rect 44456 18751 44508 18760
rect 44456 18717 44465 18751
rect 44465 18717 44499 18751
rect 44499 18717 44508 18751
rect 56876 18751 56928 18760
rect 44456 18708 44508 18717
rect 56876 18717 56885 18751
rect 56885 18717 56919 18751
rect 56919 18717 56928 18751
rect 56876 18708 56928 18717
rect 56968 18708 57020 18760
rect 38384 18572 38436 18624
rect 41880 18572 41932 18624
rect 42432 18572 42484 18624
rect 43444 18615 43496 18624
rect 43444 18581 43453 18615
rect 43453 18581 43487 18615
rect 43487 18581 43496 18615
rect 43444 18572 43496 18581
rect 43904 18640 43956 18692
rect 43996 18615 44048 18624
rect 43996 18581 44005 18615
rect 44005 18581 44039 18615
rect 44039 18581 44048 18615
rect 43996 18572 44048 18581
rect 59176 18572 59228 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 11244 18368 11296 18420
rect 13084 18368 13136 18420
rect 16856 18368 16908 18420
rect 18696 18368 18748 18420
rect 19248 18368 19300 18420
rect 19984 18368 20036 18420
rect 20352 18411 20404 18420
rect 11152 18300 11204 18352
rect 16120 18300 16172 18352
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 14924 18232 14976 18284
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 17132 18275 17184 18284
rect 17132 18241 17141 18275
rect 17141 18241 17175 18275
rect 17175 18241 17184 18275
rect 17132 18232 17184 18241
rect 17316 18232 17368 18284
rect 17500 18300 17552 18352
rect 7564 18096 7616 18148
rect 14740 18096 14792 18148
rect 15292 18207 15344 18216
rect 15292 18173 15301 18207
rect 15301 18173 15335 18207
rect 15335 18173 15344 18207
rect 15292 18164 15344 18173
rect 15568 18164 15620 18216
rect 16948 18164 17000 18216
rect 18052 18232 18104 18284
rect 20076 18300 20128 18352
rect 20352 18377 20361 18411
rect 20361 18377 20395 18411
rect 20395 18377 20404 18411
rect 20352 18368 20404 18377
rect 22468 18368 22520 18420
rect 27436 18368 27488 18420
rect 29736 18368 29788 18420
rect 22100 18300 22152 18352
rect 20996 18232 21048 18284
rect 22928 18300 22980 18352
rect 25136 18300 25188 18352
rect 27712 18300 27764 18352
rect 22468 18232 22520 18284
rect 25780 18232 25832 18284
rect 26332 18232 26384 18284
rect 26976 18232 27028 18284
rect 27160 18275 27212 18284
rect 27160 18241 27169 18275
rect 27169 18241 27203 18275
rect 27203 18241 27212 18275
rect 27160 18232 27212 18241
rect 28908 18300 28960 18352
rect 28080 18275 28132 18284
rect 28080 18241 28114 18275
rect 28114 18241 28132 18275
rect 20444 18164 20496 18216
rect 20628 18164 20680 18216
rect 25044 18164 25096 18216
rect 28080 18232 28132 18241
rect 28816 18232 28868 18284
rect 30380 18275 30432 18284
rect 30380 18241 30389 18275
rect 30389 18241 30423 18275
rect 30423 18241 30432 18275
rect 30380 18232 30432 18241
rect 33784 18368 33836 18420
rect 35348 18368 35400 18420
rect 35808 18368 35860 18420
rect 37740 18368 37792 18420
rect 52460 18368 52512 18420
rect 56784 18368 56836 18420
rect 58072 18368 58124 18420
rect 31024 18300 31076 18352
rect 31116 18275 31168 18284
rect 31116 18241 31125 18275
rect 31125 18241 31159 18275
rect 31159 18241 31168 18275
rect 31116 18232 31168 18241
rect 31668 18300 31720 18352
rect 31760 18300 31812 18352
rect 32312 18300 32364 18352
rect 32588 18343 32640 18352
rect 32588 18309 32597 18343
rect 32597 18309 32631 18343
rect 32631 18309 32640 18343
rect 32588 18300 32640 18309
rect 29000 18164 29052 18216
rect 30656 18164 30708 18216
rect 30748 18207 30800 18216
rect 30748 18173 30757 18207
rect 30757 18173 30791 18207
rect 30791 18173 30800 18207
rect 30748 18164 30800 18173
rect 23388 18096 23440 18148
rect 33140 18232 33192 18284
rect 33508 18275 33560 18284
rect 33508 18241 33517 18275
rect 33517 18241 33551 18275
rect 33551 18241 33560 18275
rect 33508 18232 33560 18241
rect 34244 18300 34296 18352
rect 34520 18300 34572 18352
rect 35624 18300 35676 18352
rect 39212 18343 39264 18352
rect 39212 18309 39221 18343
rect 39221 18309 39255 18343
rect 39255 18309 39264 18343
rect 39212 18300 39264 18309
rect 33876 18275 33928 18284
rect 33876 18241 33885 18275
rect 33885 18241 33919 18275
rect 33919 18241 33928 18275
rect 33876 18232 33928 18241
rect 33968 18164 34020 18216
rect 34428 18275 34480 18284
rect 34428 18241 34438 18275
rect 34438 18241 34472 18275
rect 34472 18241 34480 18275
rect 34428 18232 34480 18241
rect 34704 18275 34756 18284
rect 34704 18241 34713 18275
rect 34713 18241 34747 18275
rect 34747 18241 34756 18275
rect 34704 18232 34756 18241
rect 34888 18232 34940 18284
rect 35348 18232 35400 18284
rect 38108 18275 38160 18284
rect 38108 18241 38117 18275
rect 38117 18241 38151 18275
rect 38151 18241 38160 18275
rect 38108 18232 38160 18241
rect 38384 18275 38436 18284
rect 38384 18241 38393 18275
rect 38393 18241 38427 18275
rect 38427 18241 38436 18275
rect 38384 18232 38436 18241
rect 38844 18275 38896 18284
rect 38844 18241 38853 18275
rect 38853 18241 38887 18275
rect 38887 18241 38896 18275
rect 38844 18232 38896 18241
rect 39672 18232 39724 18284
rect 41236 18300 41288 18352
rect 56508 18300 56560 18352
rect 18420 18071 18472 18080
rect 18420 18037 18429 18071
rect 18429 18037 18463 18071
rect 18463 18037 18472 18071
rect 18420 18028 18472 18037
rect 18604 18028 18656 18080
rect 20628 18028 20680 18080
rect 23664 18028 23716 18080
rect 26332 18028 26384 18080
rect 26424 18028 26476 18080
rect 32680 18096 32732 18148
rect 36084 18164 36136 18216
rect 38568 18164 38620 18216
rect 41052 18232 41104 18284
rect 41788 18275 41840 18284
rect 41788 18241 41797 18275
rect 41797 18241 41831 18275
rect 41831 18241 41840 18275
rect 41788 18232 41840 18241
rect 42616 18275 42668 18284
rect 40040 18164 40092 18216
rect 42616 18241 42625 18275
rect 42625 18241 42659 18275
rect 42659 18241 42668 18275
rect 42616 18232 42668 18241
rect 43168 18232 43220 18284
rect 56692 18232 56744 18284
rect 57888 18300 57940 18352
rect 57980 18232 58032 18284
rect 35256 18096 35308 18148
rect 29184 18071 29236 18080
rect 29184 18037 29193 18071
rect 29193 18037 29227 18071
rect 29227 18037 29236 18071
rect 29184 18028 29236 18037
rect 30748 18028 30800 18080
rect 32772 18028 32824 18080
rect 33324 18071 33376 18080
rect 33324 18037 33333 18071
rect 33333 18037 33367 18071
rect 33367 18037 33376 18071
rect 33324 18028 33376 18037
rect 34704 18028 34756 18080
rect 36360 18028 36412 18080
rect 38844 18028 38896 18080
rect 40224 18028 40276 18080
rect 44272 18096 44324 18148
rect 43996 18071 44048 18080
rect 43996 18037 44005 18071
rect 44005 18037 44039 18071
rect 44039 18037 44048 18071
rect 43996 18028 44048 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 14832 17824 14884 17876
rect 17592 17756 17644 17808
rect 17684 17756 17736 17808
rect 19892 17756 19944 17808
rect 20260 17824 20312 17876
rect 33048 17824 33100 17876
rect 41788 17867 41840 17876
rect 25780 17799 25832 17808
rect 25780 17765 25789 17799
rect 25789 17765 25823 17799
rect 25823 17765 25832 17799
rect 25780 17756 25832 17765
rect 26148 17756 26200 17808
rect 30104 17756 30156 17808
rect 30288 17799 30340 17808
rect 30288 17765 30297 17799
rect 30297 17765 30331 17799
rect 30331 17765 30340 17799
rect 30288 17756 30340 17765
rect 32772 17756 32824 17808
rect 35348 17756 35400 17808
rect 2044 17620 2096 17672
rect 15660 17663 15712 17672
rect 15660 17629 15669 17663
rect 15669 17629 15703 17663
rect 15703 17629 15712 17663
rect 15660 17620 15712 17629
rect 17408 17663 17460 17672
rect 17408 17629 17417 17663
rect 17417 17629 17451 17663
rect 17451 17629 17460 17663
rect 17408 17620 17460 17629
rect 18144 17620 18196 17672
rect 1860 17595 1912 17604
rect 1860 17561 1869 17595
rect 1869 17561 1903 17595
rect 1903 17561 1912 17595
rect 1860 17552 1912 17561
rect 17132 17552 17184 17604
rect 17316 17552 17368 17604
rect 17960 17552 18012 17604
rect 19064 17620 19116 17672
rect 19340 17620 19392 17672
rect 22468 17688 22520 17740
rect 25320 17731 25372 17740
rect 25320 17697 25329 17731
rect 25329 17697 25363 17731
rect 25363 17697 25372 17731
rect 25320 17688 25372 17697
rect 27988 17688 28040 17740
rect 30748 17688 30800 17740
rect 23388 17620 23440 17672
rect 24860 17620 24912 17672
rect 13084 17484 13136 17536
rect 17684 17484 17736 17536
rect 18328 17484 18380 17536
rect 20352 17552 20404 17604
rect 22928 17552 22980 17604
rect 25504 17620 25556 17672
rect 29184 17620 29236 17672
rect 27896 17552 27948 17604
rect 29092 17552 29144 17604
rect 30564 17620 30616 17672
rect 30840 17663 30892 17672
rect 30840 17629 30849 17663
rect 30849 17629 30883 17663
rect 30883 17629 30892 17663
rect 31116 17663 31168 17672
rect 30840 17620 30892 17629
rect 31116 17629 31125 17663
rect 31125 17629 31159 17663
rect 31159 17629 31168 17663
rect 31116 17620 31168 17629
rect 31576 17620 31628 17672
rect 32036 17663 32088 17672
rect 32036 17629 32045 17663
rect 32045 17629 32079 17663
rect 32079 17629 32088 17663
rect 32036 17620 32088 17629
rect 32864 17620 32916 17672
rect 33508 17688 33560 17740
rect 33140 17663 33192 17672
rect 33140 17629 33149 17663
rect 33149 17629 33183 17663
rect 33183 17629 33192 17663
rect 33140 17620 33192 17629
rect 29460 17552 29512 17604
rect 30196 17552 30248 17604
rect 31944 17595 31996 17604
rect 31944 17561 31953 17595
rect 31953 17561 31987 17595
rect 31987 17561 31996 17595
rect 31944 17552 31996 17561
rect 32588 17552 32640 17604
rect 33232 17552 33284 17604
rect 36544 17620 36596 17672
rect 33968 17552 34020 17604
rect 41788 17833 41797 17867
rect 41797 17833 41831 17867
rect 41831 17833 41840 17867
rect 41788 17824 41840 17833
rect 42248 17756 42300 17808
rect 37924 17688 37976 17740
rect 58164 17731 58216 17740
rect 37832 17620 37884 17672
rect 38108 17620 38160 17672
rect 41236 17620 41288 17672
rect 58164 17697 58173 17731
rect 58173 17697 58207 17731
rect 58207 17697 58216 17731
rect 58164 17688 58216 17697
rect 37740 17552 37792 17604
rect 42432 17663 42484 17672
rect 42432 17629 42441 17663
rect 42441 17629 42475 17663
rect 42475 17629 42484 17663
rect 42432 17620 42484 17629
rect 43996 17620 44048 17672
rect 57060 17595 57112 17604
rect 57060 17561 57069 17595
rect 57069 17561 57103 17595
rect 57103 17561 57112 17595
rect 57060 17552 57112 17561
rect 18972 17484 19024 17536
rect 20444 17484 20496 17536
rect 21916 17484 21968 17536
rect 23940 17527 23992 17536
rect 23940 17493 23949 17527
rect 23949 17493 23983 17527
rect 23983 17493 23992 17527
rect 23940 17484 23992 17493
rect 25044 17484 25096 17536
rect 25320 17484 25372 17536
rect 30104 17484 30156 17536
rect 30380 17484 30432 17536
rect 31760 17484 31812 17536
rect 32772 17484 32824 17536
rect 33048 17484 33100 17536
rect 41052 17484 41104 17536
rect 46204 17484 46256 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 15660 17280 15712 17332
rect 16948 17280 17000 17332
rect 2136 17212 2188 17264
rect 11612 17212 11664 17264
rect 12348 17144 12400 17196
rect 17040 17144 17092 17196
rect 17408 17187 17460 17196
rect 17408 17153 17417 17187
rect 17417 17153 17451 17187
rect 17451 17153 17460 17187
rect 17408 17144 17460 17153
rect 18420 17280 18472 17332
rect 19156 17280 19208 17332
rect 17684 17212 17736 17264
rect 18880 17212 18932 17264
rect 17868 17187 17920 17196
rect 17868 17153 17877 17187
rect 17877 17153 17911 17187
rect 17911 17153 17920 17187
rect 19064 17212 19116 17264
rect 24308 17280 24360 17332
rect 24400 17280 24452 17332
rect 30196 17280 30248 17332
rect 30380 17280 30432 17332
rect 30564 17280 30616 17332
rect 31852 17280 31904 17332
rect 33508 17280 33560 17332
rect 39396 17280 39448 17332
rect 40960 17280 41012 17332
rect 41052 17280 41104 17332
rect 41236 17280 41288 17332
rect 45560 17280 45612 17332
rect 21088 17212 21140 17264
rect 21180 17212 21232 17264
rect 17868 17144 17920 17153
rect 1768 17119 1820 17128
rect 1768 17085 1777 17119
rect 1777 17085 1811 17119
rect 1811 17085 1820 17119
rect 1768 17076 1820 17085
rect 14740 17076 14792 17128
rect 19892 17144 19944 17196
rect 20076 17144 20128 17196
rect 20352 17187 20404 17196
rect 19248 17119 19300 17128
rect 19248 17085 19257 17119
rect 19257 17085 19291 17119
rect 19291 17085 19300 17119
rect 19248 17076 19300 17085
rect 19432 17076 19484 17128
rect 20352 17153 20361 17187
rect 20361 17153 20395 17187
rect 20395 17153 20404 17187
rect 20352 17144 20404 17153
rect 21916 17144 21968 17196
rect 22652 17144 22704 17196
rect 23940 17212 23992 17264
rect 25504 17212 25556 17264
rect 25688 17212 25740 17264
rect 26148 17212 26200 17264
rect 26240 17187 26292 17196
rect 26240 17153 26249 17187
rect 26249 17153 26283 17187
rect 26283 17153 26292 17187
rect 26240 17144 26292 17153
rect 27068 17212 27120 17264
rect 28908 17255 28960 17264
rect 28908 17221 28917 17255
rect 28917 17221 28951 17255
rect 28951 17221 28960 17255
rect 28908 17212 28960 17221
rect 29460 17212 29512 17264
rect 26424 17187 26476 17196
rect 26424 17153 26433 17187
rect 26433 17153 26467 17187
rect 26467 17153 26476 17187
rect 26424 17144 26476 17153
rect 17132 17008 17184 17060
rect 17500 17008 17552 17060
rect 18880 17008 18932 17060
rect 25412 17076 25464 17128
rect 29828 17144 29880 17196
rect 31668 17212 31720 17264
rect 26884 17076 26936 17128
rect 29736 17076 29788 17128
rect 30472 17144 30524 17196
rect 31484 17144 31536 17196
rect 31944 17144 31996 17196
rect 33232 17212 33284 17264
rect 35900 17212 35952 17264
rect 38108 17212 38160 17264
rect 32312 17187 32364 17196
rect 32312 17153 32321 17187
rect 32321 17153 32355 17187
rect 32355 17153 32364 17187
rect 32312 17144 32364 17153
rect 32772 17144 32824 17196
rect 30932 17076 30984 17128
rect 32128 17076 32180 17128
rect 15200 16940 15252 16992
rect 16672 16940 16724 16992
rect 21180 16940 21232 16992
rect 25504 17008 25556 17060
rect 25688 16940 25740 16992
rect 29552 16940 29604 16992
rect 29736 16983 29788 16992
rect 29736 16949 29745 16983
rect 29745 16949 29779 16983
rect 29779 16949 29788 16983
rect 29736 16940 29788 16949
rect 30196 17008 30248 17060
rect 31116 17008 31168 17060
rect 31024 16940 31076 16992
rect 31852 16940 31904 16992
rect 32312 16940 32364 16992
rect 33784 17187 33836 17196
rect 33784 17153 33798 17187
rect 33798 17153 33832 17187
rect 33832 17153 33836 17187
rect 33784 17144 33836 17153
rect 33968 17144 34020 17196
rect 34704 17187 34756 17196
rect 34704 17153 34713 17187
rect 34713 17153 34747 17187
rect 34747 17153 34756 17187
rect 34704 17144 34756 17153
rect 39028 17187 39080 17196
rect 39028 17153 39037 17187
rect 39037 17153 39071 17187
rect 39071 17153 39080 17187
rect 39028 17144 39080 17153
rect 40040 17212 40092 17264
rect 40592 17212 40644 17264
rect 40408 17144 40460 17196
rect 41420 17144 41472 17196
rect 57060 17187 57112 17196
rect 57060 17153 57069 17187
rect 57069 17153 57103 17187
rect 57103 17153 57112 17187
rect 57060 17144 57112 17153
rect 36820 17076 36872 17128
rect 37004 17076 37056 17128
rect 46204 17076 46256 17128
rect 57336 17119 57388 17128
rect 57336 17085 57345 17119
rect 57345 17085 57379 17119
rect 57379 17085 57388 17119
rect 57336 17076 57388 17085
rect 33600 17008 33652 17060
rect 33968 17051 34020 17060
rect 33968 17017 33977 17051
rect 33977 17017 34011 17051
rect 34011 17017 34020 17051
rect 33968 17008 34020 17017
rect 40684 17008 40736 17060
rect 39764 16940 39816 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 14832 16736 14884 16788
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 2228 16600 2280 16652
rect 11336 16643 11388 16652
rect 11336 16609 11345 16643
rect 11345 16609 11379 16643
rect 11379 16609 11388 16643
rect 11336 16600 11388 16609
rect 14740 16643 14792 16652
rect 14740 16609 14749 16643
rect 14749 16609 14783 16643
rect 14783 16609 14792 16643
rect 14740 16600 14792 16609
rect 11244 16575 11296 16584
rect 11244 16541 11253 16575
rect 11253 16541 11287 16575
rect 11287 16541 11296 16575
rect 11244 16532 11296 16541
rect 11612 16575 11664 16584
rect 11612 16541 11621 16575
rect 11621 16541 11655 16575
rect 11655 16541 11664 16575
rect 11612 16532 11664 16541
rect 14924 16575 14976 16584
rect 14924 16541 14933 16575
rect 14933 16541 14967 16575
rect 14967 16541 14976 16575
rect 14924 16532 14976 16541
rect 10508 16464 10560 16516
rect 12348 16396 12400 16448
rect 14924 16396 14976 16448
rect 16212 16575 16264 16584
rect 16212 16541 16221 16575
rect 16221 16541 16255 16575
rect 16255 16541 16264 16575
rect 16212 16532 16264 16541
rect 16672 16575 16724 16584
rect 16672 16541 16681 16575
rect 16681 16541 16715 16575
rect 16715 16541 16724 16575
rect 16672 16532 16724 16541
rect 22560 16736 22612 16788
rect 22928 16779 22980 16788
rect 22928 16745 22937 16779
rect 22937 16745 22971 16779
rect 22971 16745 22980 16779
rect 22928 16736 22980 16745
rect 24584 16779 24636 16788
rect 24584 16745 24593 16779
rect 24593 16745 24627 16779
rect 24627 16745 24636 16779
rect 24584 16736 24636 16745
rect 24860 16736 24912 16788
rect 26148 16736 26200 16788
rect 21364 16668 21416 16720
rect 18972 16600 19024 16652
rect 19892 16600 19944 16652
rect 24400 16600 24452 16652
rect 24492 16600 24544 16652
rect 25688 16668 25740 16720
rect 17592 16575 17644 16584
rect 16580 16464 16632 16516
rect 16764 16464 16816 16516
rect 17592 16541 17601 16575
rect 17601 16541 17635 16575
rect 17635 16541 17644 16575
rect 17592 16532 17644 16541
rect 17776 16532 17828 16584
rect 18512 16575 18564 16584
rect 16028 16396 16080 16448
rect 18512 16541 18521 16575
rect 18521 16541 18555 16575
rect 18555 16541 18564 16575
rect 18512 16532 18564 16541
rect 18788 16575 18840 16584
rect 18788 16541 18797 16575
rect 18797 16541 18831 16575
rect 18831 16541 18840 16575
rect 18788 16532 18840 16541
rect 19064 16532 19116 16584
rect 19248 16532 19300 16584
rect 20628 16575 20680 16584
rect 20628 16541 20637 16575
rect 20637 16541 20671 16575
rect 20671 16541 20680 16575
rect 20628 16532 20680 16541
rect 21732 16575 21784 16584
rect 21732 16541 21741 16575
rect 21741 16541 21775 16575
rect 21775 16541 21784 16575
rect 21732 16532 21784 16541
rect 26884 16668 26936 16720
rect 25136 16575 25188 16584
rect 25136 16541 25145 16575
rect 25145 16541 25179 16575
rect 25179 16541 25188 16575
rect 25136 16532 25188 16541
rect 25412 16532 25464 16584
rect 26332 16600 26384 16652
rect 30472 16736 30524 16788
rect 28540 16668 28592 16720
rect 29368 16668 29420 16720
rect 37740 16736 37792 16788
rect 40040 16779 40092 16788
rect 40040 16745 40049 16779
rect 40049 16745 40083 16779
rect 40083 16745 40092 16779
rect 40040 16736 40092 16745
rect 34428 16668 34480 16720
rect 29828 16643 29880 16652
rect 26240 16575 26292 16584
rect 26240 16541 26249 16575
rect 26249 16541 26283 16575
rect 26283 16541 26292 16575
rect 26240 16532 26292 16541
rect 26884 16575 26936 16584
rect 26884 16541 26893 16575
rect 26893 16541 26927 16575
rect 26927 16541 26936 16575
rect 26884 16532 26936 16541
rect 18972 16464 19024 16516
rect 20444 16464 20496 16516
rect 21180 16464 21232 16516
rect 18788 16396 18840 16448
rect 20996 16396 21048 16448
rect 25412 16439 25464 16448
rect 25412 16405 25421 16439
rect 25421 16405 25455 16439
rect 25455 16405 25464 16439
rect 25412 16396 25464 16405
rect 27436 16396 27488 16448
rect 29828 16609 29837 16643
rect 29837 16609 29871 16643
rect 29871 16609 29880 16643
rect 29828 16600 29880 16609
rect 31760 16600 31812 16652
rect 29736 16532 29788 16584
rect 31576 16532 31628 16584
rect 32312 16600 32364 16652
rect 36728 16600 36780 16652
rect 37924 16600 37976 16652
rect 39120 16600 39172 16652
rect 40592 16643 40644 16652
rect 40592 16609 40601 16643
rect 40601 16609 40635 16643
rect 40635 16609 40644 16643
rect 40592 16600 40644 16609
rect 52000 16600 52052 16652
rect 56876 16643 56928 16652
rect 32036 16532 32088 16584
rect 36176 16532 36228 16584
rect 39672 16532 39724 16584
rect 42432 16532 42484 16584
rect 56600 16532 56652 16584
rect 56876 16609 56885 16643
rect 56885 16609 56919 16643
rect 56919 16609 56928 16643
rect 56876 16600 56928 16609
rect 30564 16464 30616 16516
rect 32404 16464 32456 16516
rect 30748 16396 30800 16448
rect 40868 16464 40920 16516
rect 56048 16464 56100 16516
rect 36268 16439 36320 16448
rect 36268 16405 36277 16439
rect 36277 16405 36311 16439
rect 36311 16405 36320 16439
rect 36268 16396 36320 16405
rect 36820 16396 36872 16448
rect 56968 16396 57020 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 12532 16192 12584 16244
rect 16764 16192 16816 16244
rect 17408 16192 17460 16244
rect 18972 16192 19024 16244
rect 19064 16192 19116 16244
rect 16580 16124 16632 16176
rect 2688 16056 2740 16108
rect 1768 16031 1820 16040
rect 1768 15997 1777 16031
rect 1777 15997 1811 16031
rect 1811 15997 1820 16031
rect 1768 15988 1820 15997
rect 16212 16056 16264 16108
rect 16856 16056 16908 16108
rect 17500 16124 17552 16176
rect 17316 16099 17368 16108
rect 17316 16065 17325 16099
rect 17325 16065 17359 16099
rect 17359 16065 17368 16099
rect 17316 16056 17368 16065
rect 17960 16056 18012 16108
rect 18236 16099 18288 16108
rect 18236 16065 18245 16099
rect 18245 16065 18279 16099
rect 18279 16065 18288 16099
rect 18236 16056 18288 16065
rect 18788 16099 18840 16108
rect 18788 16065 18797 16099
rect 18797 16065 18831 16099
rect 18831 16065 18840 16099
rect 18788 16056 18840 16065
rect 18880 16056 18932 16108
rect 17224 15988 17276 16040
rect 17592 15988 17644 16040
rect 22652 16192 22704 16244
rect 26884 16192 26936 16244
rect 19984 16056 20036 16108
rect 21180 16099 21232 16108
rect 21180 16065 21189 16099
rect 21189 16065 21223 16099
rect 21223 16065 21232 16099
rect 21180 16056 21232 16065
rect 21456 16099 21508 16108
rect 21456 16065 21465 16099
rect 21465 16065 21499 16099
rect 21499 16065 21508 16099
rect 21456 16056 21508 16065
rect 24860 16124 24912 16176
rect 19340 16031 19392 16040
rect 19340 15997 19349 16031
rect 19349 15997 19383 16031
rect 19383 15997 19392 16031
rect 19340 15988 19392 15997
rect 18880 15963 18932 15972
rect 18880 15929 18889 15963
rect 18889 15929 18923 15963
rect 18923 15929 18932 15963
rect 18880 15920 18932 15929
rect 19248 15920 19300 15972
rect 15752 15852 15804 15904
rect 18512 15852 18564 15904
rect 22468 16031 22520 16040
rect 22468 15997 22477 16031
rect 22477 15997 22511 16031
rect 22511 15997 22520 16031
rect 22468 15988 22520 15997
rect 24584 16056 24636 16108
rect 24952 16056 25004 16108
rect 32588 16192 32640 16244
rect 33968 16192 34020 16244
rect 34060 16192 34112 16244
rect 34520 16192 34572 16244
rect 29552 16124 29604 16176
rect 28908 16056 28960 16108
rect 32772 16056 32824 16108
rect 36268 16056 36320 16108
rect 40500 16124 40552 16176
rect 48136 16124 48188 16176
rect 39764 16099 39816 16108
rect 39764 16065 39798 16099
rect 39798 16065 39816 16099
rect 39764 16056 39816 16065
rect 56600 16192 56652 16244
rect 56140 16124 56192 16176
rect 56968 16167 57020 16176
rect 56968 16133 56977 16167
rect 56977 16133 57011 16167
rect 57011 16133 57020 16167
rect 56968 16124 57020 16133
rect 58072 16056 58124 16108
rect 27068 15988 27120 16040
rect 26148 15920 26200 15972
rect 20720 15895 20772 15904
rect 20720 15861 20729 15895
rect 20729 15861 20763 15895
rect 20763 15861 20772 15895
rect 20720 15852 20772 15861
rect 23480 15852 23532 15904
rect 24124 15852 24176 15904
rect 25964 15852 26016 15904
rect 31024 15988 31076 16040
rect 34244 16031 34296 16040
rect 34244 15997 34253 16031
rect 34253 15997 34287 16031
rect 34287 15997 34296 16031
rect 34244 15988 34296 15997
rect 34704 15920 34756 15972
rect 40868 15963 40920 15972
rect 40868 15929 40877 15963
rect 40877 15929 40911 15963
rect 40911 15929 40920 15963
rect 40868 15920 40920 15929
rect 33140 15852 33192 15904
rect 36820 15895 36872 15904
rect 36820 15861 36829 15895
rect 36829 15861 36863 15895
rect 36863 15861 36872 15895
rect 36820 15852 36872 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 23296 15648 23348 15700
rect 21732 15580 21784 15632
rect 22560 15580 22612 15632
rect 25320 15648 25372 15700
rect 29460 15648 29512 15700
rect 48136 15691 48188 15700
rect 34704 15580 34756 15632
rect 11244 15512 11296 15564
rect 19340 15512 19392 15564
rect 21180 15512 21232 15564
rect 22468 15512 22520 15564
rect 26424 15512 26476 15564
rect 34796 15512 34848 15564
rect 36728 15580 36780 15632
rect 48136 15657 48145 15691
rect 48145 15657 48179 15691
rect 48179 15657 48188 15691
rect 48136 15648 48188 15657
rect 14004 15444 14056 15496
rect 15476 15444 15528 15496
rect 17684 15444 17736 15496
rect 19524 15444 19576 15496
rect 19984 15444 20036 15496
rect 20720 15444 20772 15496
rect 23572 15487 23624 15496
rect 23572 15453 23581 15487
rect 23581 15453 23615 15487
rect 23615 15453 23624 15487
rect 23572 15444 23624 15453
rect 26884 15487 26936 15496
rect 26884 15453 26893 15487
rect 26893 15453 26927 15487
rect 26927 15453 26936 15487
rect 26884 15444 26936 15453
rect 29736 15487 29788 15496
rect 29736 15453 29745 15487
rect 29745 15453 29779 15487
rect 29779 15453 29788 15487
rect 29736 15444 29788 15453
rect 29920 15444 29972 15496
rect 39948 15444 40000 15496
rect 1860 15419 1912 15428
rect 1860 15385 1869 15419
rect 1869 15385 1903 15419
rect 1903 15385 1912 15419
rect 1860 15376 1912 15385
rect 18512 15419 18564 15428
rect 18512 15385 18521 15419
rect 18521 15385 18555 15419
rect 18555 15385 18564 15419
rect 18512 15376 18564 15385
rect 23848 15376 23900 15428
rect 25688 15376 25740 15428
rect 29276 15376 29328 15428
rect 30104 15376 30156 15428
rect 35808 15376 35860 15428
rect 56048 15444 56100 15496
rect 57980 15487 58032 15496
rect 57980 15453 57989 15487
rect 57989 15453 58023 15487
rect 58023 15453 58032 15487
rect 57980 15444 58032 15453
rect 46848 15419 46900 15428
rect 46848 15385 46857 15419
rect 46857 15385 46891 15419
rect 46891 15385 46900 15419
rect 46848 15376 46900 15385
rect 57244 15419 57296 15428
rect 57244 15385 57253 15419
rect 57253 15385 57287 15419
rect 57287 15385 57296 15419
rect 57244 15376 57296 15385
rect 15108 15308 15160 15360
rect 16672 15308 16724 15360
rect 20812 15308 20864 15360
rect 21456 15351 21508 15360
rect 21456 15317 21465 15351
rect 21465 15317 21499 15351
rect 21499 15317 21508 15351
rect 21456 15308 21508 15317
rect 23204 15351 23256 15360
rect 23204 15317 23213 15351
rect 23213 15317 23247 15351
rect 23247 15317 23256 15351
rect 23204 15308 23256 15317
rect 23296 15351 23348 15360
rect 23296 15317 23305 15351
rect 23305 15317 23339 15351
rect 23339 15317 23348 15351
rect 23296 15308 23348 15317
rect 26884 15308 26936 15360
rect 29092 15351 29144 15360
rect 29092 15317 29101 15351
rect 29101 15317 29135 15351
rect 29135 15317 29144 15351
rect 29092 15308 29144 15317
rect 34980 15308 35032 15360
rect 35348 15351 35400 15360
rect 35348 15317 35357 15351
rect 35357 15317 35391 15351
rect 35391 15317 35400 15351
rect 35348 15308 35400 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 14924 15104 14976 15156
rect 19340 15104 19392 15156
rect 32404 15104 32456 15156
rect 18512 15036 18564 15088
rect 16764 14968 16816 15020
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 13820 14900 13872 14952
rect 14648 14943 14700 14952
rect 14648 14909 14657 14943
rect 14657 14909 14691 14943
rect 14691 14909 14700 14943
rect 14648 14900 14700 14909
rect 14924 14943 14976 14952
rect 14924 14909 14933 14943
rect 14933 14909 14967 14943
rect 14967 14909 14976 14943
rect 14924 14900 14976 14909
rect 17224 14900 17276 14952
rect 19984 15036 20036 15088
rect 21456 15036 21508 15088
rect 24124 15036 24176 15088
rect 19340 14968 19392 15020
rect 19432 14900 19484 14952
rect 22008 14900 22060 14952
rect 22468 14943 22520 14952
rect 22468 14909 22477 14943
rect 22477 14909 22511 14943
rect 22511 14909 22520 14943
rect 22468 14900 22520 14909
rect 26976 15036 27028 15088
rect 30196 15036 30248 15088
rect 26332 14968 26384 15020
rect 27160 15011 27212 15020
rect 27160 14977 27169 15011
rect 27169 14977 27203 15011
rect 27203 14977 27212 15011
rect 27160 14968 27212 14977
rect 29828 14968 29880 15020
rect 30288 15011 30340 15020
rect 30288 14977 30297 15011
rect 30297 14977 30331 15011
rect 30331 14977 30340 15011
rect 30288 14968 30340 14977
rect 31116 14968 31168 15020
rect 33140 15011 33192 15020
rect 33140 14977 33174 15011
rect 33174 14977 33192 15011
rect 33140 14968 33192 14977
rect 34796 14968 34848 15020
rect 34980 15011 35032 15020
rect 34980 14977 35014 15011
rect 35014 14977 35032 15011
rect 34980 14968 35032 14977
rect 13176 14832 13228 14884
rect 18144 14832 18196 14884
rect 18420 14875 18472 14884
rect 18420 14841 18429 14875
rect 18429 14841 18463 14875
rect 18463 14841 18472 14875
rect 18420 14832 18472 14841
rect 13820 14764 13872 14816
rect 14832 14764 14884 14816
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 16580 14764 16632 14816
rect 19156 14764 19208 14816
rect 21088 14764 21140 14816
rect 21364 14807 21416 14816
rect 21364 14773 21373 14807
rect 21373 14773 21407 14807
rect 21407 14773 21416 14807
rect 21364 14764 21416 14773
rect 21456 14764 21508 14816
rect 24768 14900 24820 14952
rect 24952 14832 25004 14884
rect 24676 14764 24728 14816
rect 29736 14764 29788 14816
rect 32496 14764 32548 14816
rect 33784 14764 33836 14816
rect 34244 14807 34296 14816
rect 34244 14773 34253 14807
rect 34253 14773 34287 14807
rect 34287 14773 34296 14807
rect 34244 14764 34296 14773
rect 35348 14764 35400 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 15476 14603 15528 14612
rect 15476 14569 15485 14603
rect 15485 14569 15519 14603
rect 15519 14569 15528 14603
rect 15476 14560 15528 14569
rect 18420 14560 18472 14612
rect 23020 14560 23072 14612
rect 30656 14560 30708 14612
rect 31116 14560 31168 14612
rect 31484 14560 31536 14612
rect 36728 14560 36780 14612
rect 58072 14603 58124 14612
rect 58072 14569 58081 14603
rect 58081 14569 58115 14603
rect 58115 14569 58124 14603
rect 58072 14560 58124 14569
rect 21824 14492 21876 14544
rect 15384 14424 15436 14476
rect 13912 14356 13964 14408
rect 15844 14356 15896 14408
rect 16028 14399 16080 14408
rect 16028 14365 16037 14399
rect 16037 14365 16071 14399
rect 16071 14365 16080 14399
rect 16028 14356 16080 14365
rect 19432 14356 19484 14408
rect 20352 14356 20404 14408
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 23940 14356 23992 14408
rect 24768 14399 24820 14408
rect 24768 14365 24777 14399
rect 24777 14365 24811 14399
rect 24811 14365 24820 14399
rect 24768 14356 24820 14365
rect 1860 14331 1912 14340
rect 1860 14297 1869 14331
rect 1869 14297 1903 14331
rect 1903 14297 1912 14331
rect 1860 14288 1912 14297
rect 29276 14424 29328 14476
rect 26424 14356 26476 14408
rect 27068 14356 27120 14408
rect 29092 14399 29144 14408
rect 29092 14365 29101 14399
rect 29101 14365 29135 14399
rect 29135 14365 29144 14399
rect 29092 14356 29144 14365
rect 29184 14356 29236 14408
rect 30012 14356 30064 14408
rect 34428 14492 34480 14544
rect 30196 14424 30248 14476
rect 30932 14424 30984 14476
rect 31300 14424 31352 14476
rect 25412 14288 25464 14340
rect 29736 14288 29788 14340
rect 31024 14356 31076 14408
rect 31484 14399 31536 14408
rect 31484 14365 31493 14399
rect 31493 14365 31527 14399
rect 31527 14365 31536 14399
rect 31484 14356 31536 14365
rect 32496 14399 32548 14408
rect 25136 14263 25188 14272
rect 25136 14229 25145 14263
rect 25145 14229 25179 14263
rect 25179 14229 25188 14263
rect 25136 14220 25188 14229
rect 27160 14220 27212 14272
rect 27344 14220 27396 14272
rect 31760 14288 31812 14340
rect 31668 14220 31720 14272
rect 32496 14365 32505 14399
rect 32505 14365 32539 14399
rect 32539 14365 32548 14399
rect 32496 14356 32548 14365
rect 57980 14399 58032 14408
rect 57980 14365 57989 14399
rect 57989 14365 58023 14399
rect 58023 14365 58032 14399
rect 57980 14356 58032 14365
rect 33232 14288 33284 14340
rect 34152 14288 34204 14340
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 14924 14016 14976 14068
rect 15844 14016 15896 14068
rect 20352 14059 20404 14068
rect 20352 14025 20361 14059
rect 20361 14025 20395 14059
rect 20395 14025 20404 14059
rect 20352 14016 20404 14025
rect 22468 14016 22520 14068
rect 26884 14016 26936 14068
rect 28632 14016 28684 14068
rect 15936 13880 15988 13932
rect 14648 13812 14700 13864
rect 19156 13923 19208 13932
rect 19156 13889 19165 13923
rect 19165 13889 19199 13923
rect 19199 13889 19208 13923
rect 19156 13880 19208 13889
rect 19432 13880 19484 13932
rect 19616 13880 19668 13932
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 22008 13880 22060 13889
rect 22284 13923 22336 13932
rect 22284 13889 22318 13923
rect 22318 13889 22336 13923
rect 22284 13880 22336 13889
rect 23480 13880 23532 13932
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 18512 13855 18564 13864
rect 18512 13821 18521 13855
rect 18521 13821 18555 13855
rect 18555 13821 18564 13855
rect 18512 13812 18564 13821
rect 23664 13812 23716 13864
rect 27252 13948 27304 14000
rect 28908 13948 28960 14000
rect 30840 14016 30892 14068
rect 32312 14016 32364 14068
rect 39948 14016 40000 14068
rect 27436 13923 27488 13932
rect 27436 13889 27470 13923
rect 27470 13889 27488 13923
rect 27436 13880 27488 13889
rect 17868 13744 17920 13796
rect 21824 13744 21876 13796
rect 17592 13676 17644 13728
rect 21456 13676 21508 13728
rect 28724 13812 28776 13864
rect 30012 13812 30064 13864
rect 30748 13855 30800 13864
rect 30748 13821 30757 13855
rect 30757 13821 30791 13855
rect 30791 13821 30800 13855
rect 30748 13812 30800 13821
rect 30932 13923 30984 13932
rect 30932 13889 30941 13923
rect 30941 13889 30975 13923
rect 30975 13889 30984 13923
rect 34152 13948 34204 14000
rect 30932 13880 30984 13889
rect 32128 13880 32180 13932
rect 32404 13880 32456 13932
rect 34428 13880 34480 13932
rect 37096 13880 37148 13932
rect 50712 13880 50764 13932
rect 58256 13880 58308 13932
rect 30196 13744 30248 13796
rect 31116 13744 31168 13796
rect 28080 13676 28132 13728
rect 29000 13719 29052 13728
rect 29000 13685 29009 13719
rect 29009 13685 29043 13719
rect 29043 13685 29052 13719
rect 29000 13676 29052 13685
rect 34244 13812 34296 13864
rect 57336 13855 57388 13864
rect 57336 13821 57345 13855
rect 57345 13821 57379 13855
rect 57379 13821 57388 13855
rect 57336 13812 57388 13821
rect 31668 13744 31720 13796
rect 31852 13676 31904 13728
rect 44824 13744 44876 13796
rect 34152 13719 34204 13728
rect 34152 13685 34161 13719
rect 34161 13685 34195 13719
rect 34195 13685 34204 13719
rect 34152 13676 34204 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 17224 13472 17276 13524
rect 22100 13472 22152 13524
rect 22284 13515 22336 13524
rect 22284 13481 22293 13515
rect 22293 13481 22327 13515
rect 22327 13481 22336 13515
rect 22284 13472 22336 13481
rect 23848 13515 23900 13524
rect 23848 13481 23857 13515
rect 23857 13481 23891 13515
rect 23891 13481 23900 13515
rect 23848 13472 23900 13481
rect 34244 13515 34296 13524
rect 18880 13404 18932 13456
rect 31116 13404 31168 13456
rect 32220 13404 32272 13456
rect 34244 13481 34253 13515
rect 34253 13481 34287 13515
rect 34287 13481 34296 13515
rect 34244 13472 34296 13481
rect 58256 13515 58308 13524
rect 58256 13481 58265 13515
rect 58265 13481 58299 13515
rect 58299 13481 58308 13515
rect 58256 13472 58308 13481
rect 39304 13404 39356 13456
rect 14648 13336 14700 13388
rect 19340 13336 19392 13388
rect 21824 13336 21876 13388
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 16580 13311 16632 13320
rect 16580 13277 16589 13311
rect 16589 13277 16623 13311
rect 16623 13277 16632 13311
rect 16580 13268 16632 13277
rect 18788 13268 18840 13320
rect 21088 13311 21140 13320
rect 21088 13277 21097 13311
rect 21097 13277 21131 13311
rect 21131 13277 21140 13311
rect 21088 13268 21140 13277
rect 24768 13336 24820 13388
rect 25688 13379 25740 13388
rect 25688 13345 25697 13379
rect 25697 13345 25731 13379
rect 25731 13345 25740 13379
rect 25688 13336 25740 13345
rect 27252 13336 27304 13388
rect 17224 13200 17276 13252
rect 17868 13200 17920 13252
rect 19984 13243 20036 13252
rect 18972 13132 19024 13184
rect 19984 13209 19993 13243
rect 19993 13209 20027 13243
rect 20027 13209 20036 13243
rect 19984 13200 20036 13209
rect 19892 13132 19944 13184
rect 20628 13200 20680 13252
rect 25136 13268 25188 13320
rect 29000 13268 29052 13320
rect 30288 13268 30340 13320
rect 56876 13379 56928 13388
rect 56876 13345 56885 13379
rect 56885 13345 56919 13379
rect 56919 13345 56928 13379
rect 56876 13336 56928 13345
rect 31852 13311 31904 13320
rect 31852 13277 31861 13311
rect 31861 13277 31895 13311
rect 31895 13277 31904 13311
rect 31852 13268 31904 13277
rect 31944 13311 31996 13320
rect 31944 13277 31953 13311
rect 31953 13277 31987 13311
rect 31987 13277 31996 13311
rect 31944 13268 31996 13277
rect 25044 13200 25096 13252
rect 30840 13200 30892 13252
rect 31760 13200 31812 13252
rect 32220 13311 32272 13320
rect 32220 13277 32229 13311
rect 32229 13277 32263 13311
rect 32263 13277 32272 13311
rect 32220 13268 32272 13277
rect 33692 13200 33744 13252
rect 21456 13132 21508 13184
rect 28724 13175 28776 13184
rect 28724 13141 28733 13175
rect 28733 13141 28767 13175
rect 28767 13141 28776 13175
rect 28724 13132 28776 13141
rect 31116 13175 31168 13184
rect 31116 13141 31125 13175
rect 31125 13141 31159 13175
rect 31159 13141 31168 13175
rect 31116 13132 31168 13141
rect 46204 13200 46256 13252
rect 56784 13200 56836 13252
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 1584 12928 1636 12980
rect 12348 12792 12400 12844
rect 14648 12835 14700 12844
rect 14648 12801 14657 12835
rect 14657 12801 14691 12835
rect 14691 12801 14700 12835
rect 14648 12792 14700 12801
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 15108 12724 15160 12776
rect 18144 12928 18196 12980
rect 18972 12928 19024 12980
rect 20904 12903 20956 12912
rect 20904 12869 20913 12903
rect 20913 12869 20947 12903
rect 20947 12869 20956 12903
rect 20904 12860 20956 12869
rect 17500 12835 17552 12844
rect 17500 12801 17509 12835
rect 17509 12801 17543 12835
rect 17543 12801 17552 12835
rect 17500 12792 17552 12801
rect 20720 12835 20772 12844
rect 20720 12801 20729 12835
rect 20729 12801 20763 12835
rect 20763 12801 20772 12835
rect 20720 12792 20772 12801
rect 21640 12724 21692 12776
rect 22284 12928 22336 12980
rect 22100 12860 22152 12912
rect 25872 12928 25924 12980
rect 26240 12928 26292 12980
rect 30840 12971 30892 12980
rect 30840 12937 30849 12971
rect 30849 12937 30883 12971
rect 30883 12937 30892 12971
rect 30840 12928 30892 12937
rect 31208 12971 31260 12980
rect 31208 12937 31217 12971
rect 31217 12937 31251 12971
rect 31251 12937 31260 12971
rect 31208 12928 31260 12937
rect 33692 12971 33744 12980
rect 33692 12937 33701 12971
rect 33701 12937 33735 12971
rect 33735 12937 33744 12971
rect 33692 12928 33744 12937
rect 46204 12928 46256 12980
rect 22652 12792 22704 12844
rect 23940 12860 23992 12912
rect 23756 12792 23808 12844
rect 24124 12792 24176 12844
rect 26148 12835 26200 12844
rect 22560 12767 22612 12776
rect 21548 12656 21600 12708
rect 22560 12733 22569 12767
rect 22569 12733 22603 12767
rect 22603 12733 22612 12767
rect 22560 12724 22612 12733
rect 23204 12724 23256 12776
rect 24860 12767 24912 12776
rect 24860 12733 24869 12767
rect 24869 12733 24903 12767
rect 24903 12733 24912 12767
rect 24860 12724 24912 12733
rect 26148 12801 26157 12835
rect 26157 12801 26191 12835
rect 26191 12801 26200 12835
rect 26148 12792 26200 12801
rect 29092 12860 29144 12912
rect 26516 12792 26568 12844
rect 27068 12792 27120 12844
rect 27344 12835 27396 12844
rect 27344 12801 27353 12835
rect 27353 12801 27387 12835
rect 27387 12801 27396 12835
rect 27344 12792 27396 12801
rect 28080 12835 28132 12844
rect 28080 12801 28089 12835
rect 28089 12801 28123 12835
rect 28123 12801 28132 12835
rect 28080 12792 28132 12801
rect 33416 12860 33468 12912
rect 31208 12792 31260 12844
rect 36544 12860 36596 12912
rect 37188 12860 37240 12912
rect 46848 12860 46900 12912
rect 30196 12724 30248 12776
rect 31116 12724 31168 12776
rect 16028 12631 16080 12640
rect 16028 12597 16037 12631
rect 16037 12597 16071 12631
rect 16071 12597 16080 12631
rect 16028 12588 16080 12597
rect 20444 12631 20496 12640
rect 20444 12597 20453 12631
rect 20453 12597 20487 12631
rect 20487 12597 20496 12631
rect 20444 12588 20496 12597
rect 22468 12656 22520 12708
rect 26332 12656 26384 12708
rect 29000 12656 29052 12708
rect 32588 12724 32640 12776
rect 34152 12835 34204 12844
rect 34152 12801 34161 12835
rect 34161 12801 34195 12835
rect 34195 12801 34204 12835
rect 34152 12792 34204 12801
rect 31484 12656 31536 12708
rect 56600 12792 56652 12844
rect 58256 12835 58308 12844
rect 56416 12724 56468 12776
rect 57888 12724 57940 12776
rect 58256 12801 58265 12835
rect 58265 12801 58299 12835
rect 58299 12801 58308 12835
rect 58256 12792 58308 12801
rect 56784 12699 56836 12708
rect 56784 12665 56793 12699
rect 56793 12665 56827 12699
rect 56827 12665 56836 12699
rect 56784 12656 56836 12665
rect 23112 12588 23164 12640
rect 30656 12588 30708 12640
rect 31668 12588 31720 12640
rect 32772 12588 32824 12640
rect 37464 12588 37516 12640
rect 40776 12588 40828 12640
rect 43260 12588 43312 12640
rect 56876 12588 56928 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 12348 12384 12400 12436
rect 13820 12384 13872 12436
rect 16672 12384 16724 12436
rect 17132 12384 17184 12436
rect 19432 12384 19484 12436
rect 21824 12384 21876 12436
rect 31944 12384 31996 12436
rect 19892 12316 19944 12368
rect 20996 12316 21048 12368
rect 30196 12316 30248 12368
rect 13820 12248 13872 12300
rect 17040 12248 17092 12300
rect 17132 12248 17184 12300
rect 27160 12248 27212 12300
rect 30288 12291 30340 12300
rect 30288 12257 30297 12291
rect 30297 12257 30331 12291
rect 30331 12257 30340 12291
rect 30288 12248 30340 12257
rect 12992 12180 13044 12232
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 1860 12155 1912 12164
rect 1860 12121 1869 12155
rect 1869 12121 1903 12155
rect 1903 12121 1912 12155
rect 1860 12112 1912 12121
rect 16120 12180 16172 12232
rect 16672 12180 16724 12232
rect 18420 12180 18472 12232
rect 25504 12180 25556 12232
rect 26056 12223 26108 12232
rect 26056 12189 26065 12223
rect 26065 12189 26099 12223
rect 26099 12189 26108 12223
rect 26056 12180 26108 12189
rect 30104 12223 30156 12232
rect 30104 12189 30113 12223
rect 30113 12189 30147 12223
rect 30147 12189 30156 12223
rect 30104 12180 30156 12189
rect 17960 12112 18012 12164
rect 20444 12155 20496 12164
rect 20444 12121 20453 12155
rect 20453 12121 20487 12155
rect 20487 12121 20496 12155
rect 20444 12112 20496 12121
rect 20812 12112 20864 12164
rect 20996 12112 21048 12164
rect 22192 12112 22244 12164
rect 23204 12112 23256 12164
rect 28172 12112 28224 12164
rect 29092 12112 29144 12164
rect 33876 12180 33928 12232
rect 40040 12180 40092 12232
rect 57980 12223 58032 12232
rect 16120 12087 16172 12096
rect 16120 12053 16129 12087
rect 16129 12053 16163 12087
rect 16163 12053 16172 12087
rect 16120 12044 16172 12053
rect 16488 12044 16540 12096
rect 22284 12044 22336 12096
rect 22376 12044 22428 12096
rect 23020 12044 23072 12096
rect 23940 12044 23992 12096
rect 25044 12087 25096 12096
rect 25044 12053 25053 12087
rect 25053 12053 25087 12087
rect 25087 12053 25096 12087
rect 25044 12044 25096 12053
rect 27896 12044 27948 12096
rect 28448 12044 28500 12096
rect 29736 12087 29788 12096
rect 29736 12053 29745 12087
rect 29745 12053 29779 12087
rect 29779 12053 29788 12087
rect 29736 12044 29788 12053
rect 30196 12087 30248 12096
rect 30196 12053 30205 12087
rect 30205 12053 30239 12087
rect 30239 12053 30248 12087
rect 30196 12044 30248 12053
rect 30288 12044 30340 12096
rect 38292 12112 38344 12164
rect 57244 12155 57296 12164
rect 57244 12121 57253 12155
rect 57253 12121 57287 12155
rect 57287 12121 57296 12155
rect 57244 12112 57296 12121
rect 57980 12189 57989 12223
rect 57989 12189 58023 12223
rect 58023 12189 58032 12223
rect 57980 12180 58032 12189
rect 58256 12112 58308 12164
rect 32680 12044 32732 12096
rect 35440 12044 35492 12096
rect 37188 12044 37240 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 12992 11883 13044 11892
rect 12992 11849 13001 11883
rect 13001 11849 13035 11883
rect 13035 11849 13044 11883
rect 12992 11840 13044 11849
rect 15936 11883 15988 11892
rect 15936 11849 15945 11883
rect 15945 11849 15979 11883
rect 15979 11849 15988 11883
rect 15936 11840 15988 11849
rect 16028 11840 16080 11892
rect 16488 11840 16540 11892
rect 17040 11883 17092 11892
rect 17040 11849 17049 11883
rect 17049 11849 17083 11883
rect 17083 11849 17092 11883
rect 17040 11840 17092 11849
rect 17500 11840 17552 11892
rect 17776 11840 17828 11892
rect 19064 11840 19116 11892
rect 19432 11840 19484 11892
rect 11060 11704 11112 11756
rect 13268 11772 13320 11824
rect 17408 11772 17460 11824
rect 13820 11704 13872 11756
rect 15384 11704 15436 11756
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 19340 11772 19392 11824
rect 1768 11679 1820 11688
rect 1768 11645 1777 11679
rect 1777 11645 1811 11679
rect 1811 11645 1820 11679
rect 1768 11636 1820 11645
rect 13452 11679 13504 11688
rect 13452 11645 13461 11679
rect 13461 11645 13495 11679
rect 13495 11645 13504 11679
rect 18788 11704 18840 11756
rect 20812 11704 20864 11756
rect 13452 11636 13504 11645
rect 17960 11679 18012 11688
rect 17684 11568 17736 11620
rect 17960 11645 17969 11679
rect 17969 11645 18003 11679
rect 18003 11645 18012 11679
rect 17960 11636 18012 11645
rect 18604 11679 18656 11688
rect 18144 11568 18196 11620
rect 18604 11645 18613 11679
rect 18613 11645 18647 11679
rect 18647 11645 18656 11679
rect 19800 11679 19852 11688
rect 18604 11636 18656 11645
rect 19800 11645 19809 11679
rect 19809 11645 19843 11679
rect 19843 11645 19852 11679
rect 19800 11636 19852 11645
rect 21732 11840 21784 11892
rect 23756 11883 23808 11892
rect 23756 11849 23765 11883
rect 23765 11849 23799 11883
rect 23799 11849 23808 11883
rect 23756 11840 23808 11849
rect 25504 11883 25556 11892
rect 25504 11849 25513 11883
rect 25513 11849 25547 11883
rect 25547 11849 25556 11883
rect 25504 11840 25556 11849
rect 26056 11840 26108 11892
rect 32864 11840 32916 11892
rect 34152 11840 34204 11892
rect 22284 11772 22336 11824
rect 22100 11704 22152 11756
rect 23112 11747 23164 11756
rect 23112 11713 23121 11747
rect 23121 11713 23155 11747
rect 23155 11713 23164 11747
rect 23112 11704 23164 11713
rect 23664 11747 23716 11756
rect 23664 11713 23673 11747
rect 23673 11713 23707 11747
rect 23707 11713 23716 11747
rect 23664 11704 23716 11713
rect 23848 11747 23900 11756
rect 23848 11713 23857 11747
rect 23857 11713 23891 11747
rect 23891 11713 23900 11747
rect 23848 11704 23900 11713
rect 27252 11704 27304 11756
rect 29736 11772 29788 11824
rect 29828 11772 29880 11824
rect 30288 11772 30340 11824
rect 34336 11772 34388 11824
rect 28172 11704 28224 11756
rect 29276 11747 29328 11756
rect 29276 11713 29285 11747
rect 29285 11713 29319 11747
rect 29319 11713 29328 11747
rect 29276 11704 29328 11713
rect 30104 11704 30156 11756
rect 33692 11747 33744 11756
rect 33692 11713 33701 11747
rect 33701 11713 33735 11747
rect 33735 11713 33744 11747
rect 33692 11704 33744 11713
rect 33876 11747 33928 11756
rect 33876 11713 33883 11747
rect 33883 11713 33928 11747
rect 33876 11704 33928 11713
rect 33968 11747 34020 11756
rect 33968 11713 33977 11747
rect 33977 11713 34011 11747
rect 34011 11713 34020 11747
rect 34152 11747 34204 11756
rect 33968 11704 34020 11713
rect 34152 11713 34166 11747
rect 34166 11713 34200 11747
rect 34200 11713 34204 11747
rect 34152 11704 34204 11713
rect 35716 11840 35768 11892
rect 34612 11772 34664 11824
rect 47860 11772 47912 11824
rect 36084 11704 36136 11756
rect 37924 11704 37976 11756
rect 42708 11704 42760 11756
rect 43444 11704 43496 11756
rect 47676 11704 47728 11756
rect 51448 11704 51500 11756
rect 57152 11747 57204 11756
rect 57152 11713 57161 11747
rect 57161 11713 57195 11747
rect 57195 11713 57204 11747
rect 57152 11704 57204 11713
rect 18328 11568 18380 11620
rect 19984 11568 20036 11620
rect 19064 11543 19116 11552
rect 19064 11509 19073 11543
rect 19073 11509 19107 11543
rect 19107 11509 19116 11543
rect 21824 11568 21876 11620
rect 23020 11679 23072 11688
rect 23020 11645 23029 11679
rect 23029 11645 23063 11679
rect 23063 11645 23072 11679
rect 23020 11636 23072 11645
rect 34060 11636 34112 11688
rect 38384 11679 38436 11688
rect 25596 11568 25648 11620
rect 28448 11568 28500 11620
rect 33968 11568 34020 11620
rect 34612 11568 34664 11620
rect 38384 11645 38393 11679
rect 38393 11645 38427 11679
rect 38427 11645 38436 11679
rect 38384 11636 38436 11645
rect 19064 11500 19116 11509
rect 21732 11500 21784 11552
rect 30196 11500 30248 11552
rect 34336 11543 34388 11552
rect 34336 11509 34345 11543
rect 34345 11509 34379 11543
rect 34379 11509 34388 11543
rect 34796 11543 34848 11552
rect 34336 11500 34388 11509
rect 34796 11509 34805 11543
rect 34805 11509 34839 11543
rect 34839 11509 34848 11543
rect 34796 11500 34848 11509
rect 57244 11543 57296 11552
rect 57244 11509 57253 11543
rect 57253 11509 57287 11543
rect 57287 11509 57296 11543
rect 57244 11500 57296 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 13544 11296 13596 11348
rect 17684 11296 17736 11348
rect 9128 11228 9180 11280
rect 16212 11228 16264 11280
rect 19432 11228 19484 11280
rect 20444 11296 20496 11348
rect 20628 11296 20680 11348
rect 20812 11339 20864 11348
rect 20812 11305 20821 11339
rect 20821 11305 20855 11339
rect 20855 11305 20864 11339
rect 20812 11296 20864 11305
rect 21272 11339 21324 11348
rect 21272 11305 21281 11339
rect 21281 11305 21315 11339
rect 21315 11305 21324 11339
rect 21272 11296 21324 11305
rect 22560 11296 22612 11348
rect 23848 11296 23900 11348
rect 24584 11339 24636 11348
rect 24584 11305 24593 11339
rect 24593 11305 24627 11339
rect 24627 11305 24636 11339
rect 24584 11296 24636 11305
rect 25504 11296 25556 11348
rect 21456 11228 21508 11280
rect 12808 11160 12860 11212
rect 17132 11160 17184 11212
rect 18144 11160 18196 11212
rect 19156 11160 19208 11212
rect 14832 11092 14884 11144
rect 16028 11092 16080 11144
rect 18604 11092 18656 11144
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 20628 11092 20680 11144
rect 17500 11024 17552 11076
rect 20352 11024 20404 11076
rect 20904 11092 20956 11144
rect 21456 11092 21508 11144
rect 26424 11160 26476 11212
rect 33232 11296 33284 11348
rect 33692 11296 33744 11348
rect 34060 11296 34112 11348
rect 58256 11339 58308 11348
rect 58256 11305 58265 11339
rect 58265 11305 58299 11339
rect 58299 11305 58308 11339
rect 58256 11296 58308 11305
rect 32588 11228 32640 11280
rect 22560 11092 22612 11144
rect 23296 11092 23348 11144
rect 23388 11092 23440 11144
rect 24216 11092 24268 11144
rect 24676 11092 24728 11144
rect 25596 11135 25648 11144
rect 20996 11024 21048 11076
rect 25596 11101 25605 11135
rect 25605 11101 25639 11135
rect 25639 11101 25648 11135
rect 25596 11092 25648 11101
rect 28448 11092 28500 11144
rect 29000 11160 29052 11212
rect 34060 11160 34112 11212
rect 34612 11228 34664 11280
rect 34796 11160 34848 11212
rect 33232 11092 33284 11144
rect 34888 11135 34940 11144
rect 28264 11024 28316 11076
rect 29460 11024 29512 11076
rect 32404 11067 32456 11076
rect 32404 11033 32413 11067
rect 32413 11033 32447 11067
rect 32447 11033 32456 11067
rect 32404 11024 32456 11033
rect 32588 11067 32640 11076
rect 32588 11033 32597 11067
rect 32597 11033 32631 11067
rect 32631 11033 32640 11067
rect 32588 11024 32640 11033
rect 33784 11024 33836 11076
rect 34888 11101 34897 11135
rect 34897 11101 34931 11135
rect 34931 11101 34940 11135
rect 34888 11092 34940 11101
rect 36544 11160 36596 11212
rect 37004 11160 37056 11212
rect 37924 11160 37976 11212
rect 56876 11203 56928 11212
rect 56876 11169 56885 11203
rect 56885 11169 56919 11203
rect 56919 11169 56928 11203
rect 56876 11160 56928 11169
rect 36636 11092 36688 11144
rect 34152 11024 34204 11076
rect 34612 11024 34664 11076
rect 35900 11024 35952 11076
rect 39120 11092 39172 11144
rect 40408 11024 40460 11076
rect 56784 11024 56836 11076
rect 18052 10999 18104 11008
rect 18052 10965 18061 10999
rect 18061 10965 18095 10999
rect 18095 10965 18104 10999
rect 18052 10956 18104 10965
rect 19984 10956 20036 11008
rect 25780 10956 25832 11008
rect 25872 10956 25924 11008
rect 28356 10999 28408 11008
rect 28356 10965 28365 10999
rect 28365 10965 28399 10999
rect 28399 10965 28408 10999
rect 28356 10956 28408 10965
rect 29092 10956 29144 11008
rect 32772 10999 32824 11008
rect 32772 10965 32781 10999
rect 32781 10965 32815 10999
rect 32815 10965 32824 10999
rect 32772 10956 32824 10965
rect 33876 10956 33928 11008
rect 36452 10956 36504 11008
rect 40132 10956 40184 11008
rect 41696 10956 41748 11008
rect 49240 10956 49292 11008
rect 51264 10956 51316 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 11060 10752 11112 10804
rect 21456 10795 21508 10804
rect 17132 10684 17184 10736
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 14004 10616 14056 10668
rect 1768 10591 1820 10600
rect 1768 10557 1777 10591
rect 1777 10557 1811 10591
rect 1811 10557 1820 10591
rect 1768 10548 1820 10557
rect 12992 10548 13044 10600
rect 13360 10591 13412 10600
rect 13360 10557 13369 10591
rect 13369 10557 13403 10591
rect 13403 10557 13412 10591
rect 13360 10548 13412 10557
rect 6000 10480 6052 10532
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 15200 10591 15252 10600
rect 15200 10557 15209 10591
rect 15209 10557 15243 10591
rect 15243 10557 15252 10591
rect 17776 10591 17828 10600
rect 15200 10548 15252 10557
rect 17776 10557 17785 10591
rect 17785 10557 17819 10591
rect 17819 10557 17828 10591
rect 17776 10548 17828 10557
rect 18512 10684 18564 10736
rect 18880 10684 18932 10736
rect 20628 10684 20680 10736
rect 21456 10761 21465 10795
rect 21465 10761 21499 10795
rect 21499 10761 21508 10795
rect 21456 10752 21508 10761
rect 21640 10752 21692 10804
rect 21916 10752 21968 10804
rect 21272 10616 21324 10668
rect 18512 10548 18564 10600
rect 21640 10616 21692 10668
rect 22284 10616 22336 10668
rect 22836 10616 22888 10668
rect 24584 10684 24636 10736
rect 23940 10659 23992 10668
rect 23940 10625 23974 10659
rect 23974 10625 23992 10659
rect 23940 10616 23992 10625
rect 17132 10480 17184 10532
rect 18052 10480 18104 10532
rect 21456 10548 21508 10600
rect 22008 10548 22060 10600
rect 22192 10548 22244 10600
rect 22652 10591 22704 10600
rect 22652 10557 22661 10591
rect 22661 10557 22695 10591
rect 22695 10557 22704 10591
rect 22652 10548 22704 10557
rect 28356 10616 28408 10668
rect 27436 10591 27488 10600
rect 21548 10480 21600 10532
rect 27436 10557 27445 10591
rect 27445 10557 27479 10591
rect 27479 10557 27488 10591
rect 27436 10548 27488 10557
rect 28540 10752 28592 10804
rect 28632 10684 28684 10736
rect 33784 10684 33836 10736
rect 29276 10659 29328 10668
rect 29276 10625 29285 10659
rect 29285 10625 29319 10659
rect 29319 10625 29328 10659
rect 29276 10616 29328 10625
rect 29460 10659 29512 10668
rect 29460 10625 29469 10659
rect 29469 10625 29503 10659
rect 29503 10625 29512 10659
rect 29460 10616 29512 10625
rect 30932 10616 30984 10668
rect 34888 10684 34940 10736
rect 33968 10616 34020 10668
rect 21272 10412 21324 10464
rect 26976 10480 27028 10532
rect 28172 10480 28224 10532
rect 32404 10480 32456 10532
rect 47676 10752 47728 10804
rect 35992 10727 36044 10736
rect 35992 10693 36001 10727
rect 36001 10693 36035 10727
rect 36035 10693 36044 10727
rect 35992 10684 36044 10693
rect 56600 10684 56652 10736
rect 57152 10752 57204 10804
rect 35900 10659 35952 10668
rect 35900 10625 35909 10659
rect 35909 10625 35943 10659
rect 35943 10625 35952 10659
rect 35900 10616 35952 10625
rect 36084 10659 36136 10668
rect 36084 10625 36093 10659
rect 36093 10625 36127 10659
rect 36127 10625 36136 10659
rect 36084 10616 36136 10625
rect 37740 10659 37792 10668
rect 37740 10625 37774 10659
rect 37774 10625 37792 10659
rect 37740 10616 37792 10625
rect 35072 10548 35124 10600
rect 56600 10548 56652 10600
rect 57888 10616 57940 10668
rect 58256 10659 58308 10668
rect 58256 10625 58265 10659
rect 58265 10625 58299 10659
rect 58299 10625 58308 10659
rect 58256 10616 58308 10625
rect 36820 10480 36872 10532
rect 56784 10523 56836 10532
rect 56784 10489 56793 10523
rect 56793 10489 56827 10523
rect 56827 10489 56836 10523
rect 56784 10480 56836 10489
rect 23848 10412 23900 10464
rect 25044 10455 25096 10464
rect 25044 10421 25053 10455
rect 25053 10421 25087 10455
rect 25087 10421 25096 10455
rect 25044 10412 25096 10421
rect 26608 10455 26660 10464
rect 26608 10421 26617 10455
rect 26617 10421 26651 10455
rect 26651 10421 26660 10455
rect 26608 10412 26660 10421
rect 26792 10412 26844 10464
rect 29092 10412 29144 10464
rect 29368 10455 29420 10464
rect 29368 10421 29377 10455
rect 29377 10421 29411 10455
rect 29411 10421 29420 10455
rect 29368 10412 29420 10421
rect 29736 10412 29788 10464
rect 32312 10412 32364 10464
rect 33232 10412 33284 10464
rect 36268 10455 36320 10464
rect 36268 10421 36277 10455
rect 36277 10421 36311 10455
rect 36311 10421 36320 10455
rect 36268 10412 36320 10421
rect 38844 10455 38896 10464
rect 38844 10421 38853 10455
rect 38853 10421 38887 10455
rect 38887 10421 38896 10455
rect 38844 10412 38896 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 13452 10208 13504 10260
rect 17776 10208 17828 10260
rect 21548 10208 21600 10260
rect 22008 10208 22060 10260
rect 22652 10208 22704 10260
rect 25780 10251 25832 10260
rect 8944 10140 8996 10192
rect 8392 10072 8444 10124
rect 14924 10140 14976 10192
rect 20076 10140 20128 10192
rect 21916 10183 21968 10192
rect 21916 10149 21925 10183
rect 21925 10149 21959 10183
rect 21959 10149 21968 10183
rect 21916 10140 21968 10149
rect 25780 10217 25789 10251
rect 25789 10217 25823 10251
rect 25823 10217 25832 10251
rect 25780 10208 25832 10217
rect 28632 10208 28684 10260
rect 22468 10072 22520 10124
rect 12900 10004 12952 10056
rect 12992 10004 13044 10056
rect 1860 9979 1912 9988
rect 1860 9945 1869 9979
rect 1869 9945 1903 9979
rect 1903 9945 1912 9979
rect 1860 9936 1912 9945
rect 14004 9936 14056 9988
rect 20628 10004 20680 10056
rect 21272 10004 21324 10056
rect 21640 10004 21692 10056
rect 21732 9936 21784 9988
rect 22100 10004 22152 10056
rect 23664 10047 23716 10056
rect 23664 10013 23673 10047
rect 23673 10013 23707 10047
rect 23707 10013 23716 10047
rect 23664 10004 23716 10013
rect 23756 10047 23808 10056
rect 23756 10013 23765 10047
rect 23765 10013 23799 10047
rect 23799 10013 23808 10047
rect 23756 10004 23808 10013
rect 24216 10004 24268 10056
rect 25872 10004 25924 10056
rect 27620 10004 27672 10056
rect 30472 10208 30524 10260
rect 31668 10208 31720 10260
rect 29184 10140 29236 10192
rect 29736 10047 29788 10056
rect 29736 10013 29745 10047
rect 29745 10013 29779 10047
rect 29779 10013 29788 10047
rect 30748 10140 30800 10192
rect 30472 10072 30524 10124
rect 30932 10115 30984 10124
rect 30932 10081 30941 10115
rect 30941 10081 30975 10115
rect 30975 10081 30984 10115
rect 30932 10072 30984 10081
rect 29736 10004 29788 10013
rect 26424 9868 26476 9920
rect 26608 9936 26660 9988
rect 29644 9936 29696 9988
rect 28540 9868 28592 9920
rect 29092 9911 29144 9920
rect 29092 9877 29101 9911
rect 29101 9877 29135 9911
rect 29135 9877 29144 9911
rect 29092 9868 29144 9877
rect 29460 9868 29512 9920
rect 30380 10004 30432 10056
rect 31668 10072 31720 10124
rect 37740 10208 37792 10260
rect 38844 10140 38896 10192
rect 38384 10115 38436 10124
rect 38384 10081 38393 10115
rect 38393 10081 38427 10115
rect 38427 10081 38436 10115
rect 58164 10115 58216 10124
rect 38384 10072 38436 10081
rect 31208 10047 31260 10056
rect 31208 10013 31217 10047
rect 31217 10013 31251 10047
rect 31251 10013 31260 10047
rect 31208 10004 31260 10013
rect 35900 10004 35952 10056
rect 36360 10004 36412 10056
rect 38660 10004 38712 10056
rect 34888 9936 34940 9988
rect 58164 10081 58173 10115
rect 58173 10081 58207 10115
rect 58207 10081 58216 10115
rect 58164 10072 58216 10081
rect 42156 10004 42208 10056
rect 53840 10004 53892 10056
rect 39948 9936 40000 9988
rect 31300 9868 31352 9920
rect 32036 9868 32088 9920
rect 32956 9868 33008 9920
rect 45100 9936 45152 9988
rect 57060 9979 57112 9988
rect 57060 9945 57069 9979
rect 57069 9945 57103 9979
rect 57103 9945 57112 9979
rect 57060 9936 57112 9945
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 10508 9664 10560 9716
rect 23572 9664 23624 9716
rect 23664 9664 23716 9716
rect 14004 9639 14056 9648
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 12164 9460 12216 9512
rect 14004 9605 14013 9639
rect 14013 9605 14047 9639
rect 14047 9605 14056 9639
rect 14004 9596 14056 9605
rect 25780 9664 25832 9716
rect 25872 9596 25924 9648
rect 27436 9664 27488 9716
rect 30380 9664 30432 9716
rect 31208 9664 31260 9716
rect 31392 9664 31444 9716
rect 44824 9664 44876 9716
rect 25688 9528 25740 9580
rect 27416 9571 27468 9580
rect 27416 9537 27425 9571
rect 27425 9537 27459 9571
rect 27459 9537 27468 9571
rect 27416 9528 27468 9537
rect 29368 9596 29420 9648
rect 29552 9596 29604 9648
rect 30012 9596 30064 9648
rect 33876 9596 33928 9648
rect 34888 9596 34940 9648
rect 13360 9460 13412 9512
rect 15200 9460 15252 9512
rect 18144 9460 18196 9512
rect 12532 9392 12584 9444
rect 12716 9435 12768 9444
rect 12716 9401 12725 9435
rect 12725 9401 12759 9435
rect 12759 9401 12768 9435
rect 12716 9392 12768 9401
rect 12992 9392 13044 9444
rect 15752 9392 15804 9444
rect 20628 9460 20680 9512
rect 27068 9460 27120 9512
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 20812 9392 20864 9444
rect 23112 9392 23164 9444
rect 26700 9392 26752 9444
rect 27620 9392 27672 9444
rect 27712 9392 27764 9444
rect 28172 9528 28224 9580
rect 29460 9528 29512 9580
rect 30104 9571 30156 9580
rect 30104 9537 30113 9571
rect 30113 9537 30147 9571
rect 30147 9537 30156 9571
rect 30104 9528 30156 9537
rect 30196 9528 30248 9580
rect 31116 9571 31168 9580
rect 31116 9537 31125 9571
rect 31125 9537 31159 9571
rect 31159 9537 31168 9571
rect 31116 9528 31168 9537
rect 31208 9577 31260 9586
rect 31208 9543 31217 9577
rect 31217 9543 31251 9577
rect 31251 9543 31260 9577
rect 31208 9534 31260 9543
rect 31484 9528 31536 9580
rect 34336 9528 34388 9580
rect 35072 9571 35124 9580
rect 35072 9537 35081 9571
rect 35081 9537 35115 9571
rect 35115 9537 35124 9571
rect 35072 9528 35124 9537
rect 35716 9528 35768 9580
rect 30288 9503 30340 9512
rect 30288 9469 30297 9503
rect 30297 9469 30331 9503
rect 30331 9469 30340 9503
rect 30288 9460 30340 9469
rect 34520 9460 34572 9512
rect 30104 9392 30156 9444
rect 32036 9392 32088 9444
rect 32588 9392 32640 9444
rect 28080 9324 28132 9376
rect 28172 9367 28224 9376
rect 28172 9333 28181 9367
rect 28181 9333 28215 9367
rect 28215 9333 28224 9367
rect 28172 9324 28224 9333
rect 29552 9324 29604 9376
rect 57244 9596 57296 9648
rect 37556 9528 37608 9580
rect 37648 9460 37700 9512
rect 38292 9528 38344 9580
rect 38660 9528 38712 9580
rect 39948 9528 40000 9580
rect 40500 9571 40552 9580
rect 40500 9537 40509 9571
rect 40509 9537 40543 9571
rect 40543 9537 40552 9571
rect 40500 9528 40552 9537
rect 41052 9528 41104 9580
rect 39672 9460 39724 9512
rect 40132 9460 40184 9512
rect 40316 9460 40368 9512
rect 36636 9392 36688 9444
rect 39948 9392 40000 9444
rect 40500 9392 40552 9444
rect 41604 9392 41656 9444
rect 56324 9528 56376 9580
rect 57428 9596 57480 9648
rect 57888 9596 57940 9648
rect 57520 9571 57572 9580
rect 57520 9537 57529 9571
rect 57529 9537 57563 9571
rect 57563 9537 57572 9571
rect 57520 9528 57572 9537
rect 50068 9460 50120 9512
rect 50804 9460 50856 9512
rect 37280 9324 37332 9376
rect 37832 9324 37884 9376
rect 38016 9367 38068 9376
rect 38016 9333 38025 9367
rect 38025 9333 38059 9367
rect 38059 9333 38068 9367
rect 38016 9324 38068 9333
rect 40316 9324 40368 9376
rect 53840 9324 53892 9376
rect 58256 9324 58308 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 18236 9120 18288 9172
rect 20812 9163 20864 9172
rect 19432 9052 19484 9104
rect 20812 9129 20821 9163
rect 20821 9129 20855 9163
rect 20855 9129 20864 9163
rect 20812 9120 20864 9129
rect 27804 9120 27856 9172
rect 28080 9120 28132 9172
rect 30380 9120 30432 9172
rect 30472 9120 30524 9172
rect 31668 9120 31720 9172
rect 31852 9120 31904 9172
rect 37280 9120 37332 9172
rect 37464 9120 37516 9172
rect 37832 9120 37884 9172
rect 38108 9120 38160 9172
rect 38292 9120 38344 9172
rect 39764 9120 39816 9172
rect 39948 9120 40000 9172
rect 11796 8916 11848 8968
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 23664 8984 23716 9036
rect 24584 9027 24636 9036
rect 24584 8993 24593 9027
rect 24593 8993 24627 9027
rect 24627 8993 24636 9027
rect 24584 8984 24636 8993
rect 23572 8959 23624 8968
rect 23572 8925 23581 8959
rect 23581 8925 23615 8959
rect 23615 8925 23624 8959
rect 23572 8916 23624 8925
rect 34612 9052 34664 9104
rect 1860 8891 1912 8900
rect 1860 8857 1869 8891
rect 1869 8857 1903 8891
rect 1903 8857 1912 8891
rect 1860 8848 1912 8857
rect 16488 8848 16540 8900
rect 30472 8916 30524 8968
rect 25872 8848 25924 8900
rect 29736 8848 29788 8900
rect 31300 8916 31352 8968
rect 31668 8916 31720 8968
rect 32036 8959 32088 8968
rect 31484 8848 31536 8900
rect 31760 8848 31812 8900
rect 32036 8925 32045 8959
rect 32045 8925 32079 8959
rect 32079 8925 32088 8959
rect 32036 8916 32088 8925
rect 32128 8959 32180 8968
rect 32128 8925 32137 8959
rect 32137 8925 32171 8959
rect 32171 8925 32180 8959
rect 32128 8916 32180 8925
rect 32404 8848 32456 8900
rect 17960 8780 18012 8832
rect 19984 8780 20036 8832
rect 25964 8823 26016 8832
rect 25964 8789 25973 8823
rect 25973 8789 26007 8823
rect 26007 8789 26016 8823
rect 25964 8780 26016 8789
rect 31208 8780 31260 8832
rect 31944 8780 31996 8832
rect 34796 8916 34848 8968
rect 36268 8984 36320 9036
rect 36452 9052 36504 9104
rect 39396 9052 39448 9104
rect 40132 9052 40184 9104
rect 41052 9120 41104 9172
rect 58348 9120 58400 9172
rect 41052 9027 41104 9036
rect 32864 8848 32916 8900
rect 34888 8848 34940 8900
rect 35532 8959 35584 8968
rect 35532 8925 35541 8959
rect 35541 8925 35575 8959
rect 35575 8925 35584 8959
rect 37280 8959 37332 8968
rect 35532 8916 35584 8925
rect 37280 8925 37289 8959
rect 37289 8925 37323 8959
rect 37323 8925 37332 8959
rect 37280 8916 37332 8925
rect 38568 8916 38620 8968
rect 38752 8916 38804 8968
rect 40316 8959 40368 8968
rect 40316 8925 40325 8959
rect 40325 8925 40359 8959
rect 40359 8925 40368 8959
rect 40316 8916 40368 8925
rect 40500 8916 40552 8968
rect 41052 8993 41061 9027
rect 41061 8993 41095 9027
rect 41095 8993 41104 9027
rect 41052 8984 41104 8993
rect 43352 8984 43404 9036
rect 56876 9027 56928 9036
rect 56876 8993 56885 9027
rect 56885 8993 56919 9027
rect 56919 8993 56928 9027
rect 56876 8984 56928 8993
rect 37096 8848 37148 8900
rect 38108 8848 38160 8900
rect 38200 8848 38252 8900
rect 40224 8891 40276 8900
rect 34428 8780 34480 8832
rect 37832 8780 37884 8832
rect 38752 8780 38804 8832
rect 39028 8823 39080 8832
rect 39028 8789 39053 8823
rect 39053 8789 39080 8823
rect 39212 8823 39264 8832
rect 39028 8780 39080 8789
rect 39212 8789 39221 8823
rect 39221 8789 39255 8823
rect 39255 8789 39264 8823
rect 39212 8780 39264 8789
rect 40224 8857 40233 8891
rect 40233 8857 40267 8891
rect 40267 8857 40276 8891
rect 40224 8848 40276 8857
rect 40316 8780 40368 8832
rect 41052 8780 41104 8832
rect 50068 8916 50120 8968
rect 58072 8848 58124 8900
rect 43352 8780 43404 8832
rect 56600 8780 56652 8832
rect 57520 8780 57572 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 13084 8508 13136 8560
rect 18328 8508 18380 8560
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 12164 8415 12216 8424
rect 12164 8381 12173 8415
rect 12173 8381 12207 8415
rect 12207 8381 12216 8415
rect 12164 8372 12216 8381
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 12532 8372 12584 8424
rect 18144 8440 18196 8492
rect 19432 8508 19484 8560
rect 19984 8576 20036 8628
rect 25872 8619 25924 8628
rect 25872 8585 25881 8619
rect 25881 8585 25915 8619
rect 25915 8585 25924 8619
rect 25872 8576 25924 8585
rect 26516 8576 26568 8628
rect 29736 8619 29788 8628
rect 25964 8508 26016 8560
rect 13268 8415 13320 8424
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 17960 8372 18012 8424
rect 18604 8372 18656 8424
rect 18972 8372 19024 8424
rect 24768 8440 24820 8492
rect 29736 8585 29745 8619
rect 29745 8585 29779 8619
rect 29779 8585 29788 8619
rect 29736 8576 29788 8585
rect 30748 8576 30800 8628
rect 31576 8576 31628 8628
rect 40224 8576 40276 8628
rect 56324 8619 56376 8628
rect 56324 8585 56333 8619
rect 56333 8585 56367 8619
rect 56367 8585 56376 8619
rect 56324 8576 56376 8585
rect 57152 8576 57204 8628
rect 58256 8619 58308 8628
rect 13912 8304 13964 8356
rect 20444 8372 20496 8424
rect 11980 8236 12032 8288
rect 19064 8236 19116 8288
rect 19708 8236 19760 8288
rect 21824 8372 21876 8424
rect 23020 8372 23072 8424
rect 24216 8372 24268 8424
rect 28080 8440 28132 8492
rect 30012 8508 30064 8560
rect 32128 8508 32180 8560
rect 32404 8508 32456 8560
rect 34612 8551 34664 8560
rect 29460 8440 29512 8492
rect 30472 8483 30524 8492
rect 26424 8415 26476 8424
rect 26424 8381 26433 8415
rect 26433 8381 26467 8415
rect 26467 8381 26476 8415
rect 26424 8372 26476 8381
rect 30472 8449 30481 8483
rect 30481 8449 30515 8483
rect 30515 8449 30524 8483
rect 30472 8440 30524 8449
rect 30748 8483 30800 8492
rect 30748 8449 30757 8483
rect 30757 8449 30791 8483
rect 30791 8449 30800 8483
rect 30748 8440 30800 8449
rect 31300 8440 31352 8492
rect 31576 8483 31628 8492
rect 31576 8449 31585 8483
rect 31585 8449 31619 8483
rect 31619 8449 31628 8483
rect 31576 8440 31628 8449
rect 32312 8440 32364 8492
rect 32772 8483 32824 8492
rect 32772 8449 32781 8483
rect 32781 8449 32815 8483
rect 32815 8449 32824 8483
rect 32772 8440 32824 8449
rect 34612 8517 34621 8551
rect 34621 8517 34655 8551
rect 34655 8517 34664 8551
rect 34612 8508 34664 8517
rect 34704 8551 34756 8560
rect 34704 8517 34713 8551
rect 34713 8517 34747 8551
rect 34747 8517 34756 8551
rect 34704 8508 34756 8517
rect 25504 8304 25556 8356
rect 30380 8372 30432 8424
rect 31668 8415 31720 8424
rect 31668 8381 31677 8415
rect 31677 8381 31711 8415
rect 31711 8381 31720 8415
rect 31668 8372 31720 8381
rect 33324 8372 33376 8424
rect 33692 8415 33744 8424
rect 33692 8381 33701 8415
rect 33701 8381 33735 8415
rect 33735 8381 33744 8415
rect 33692 8372 33744 8381
rect 33968 8372 34020 8424
rect 34428 8483 34480 8492
rect 34428 8449 34438 8483
rect 34438 8449 34472 8483
rect 34472 8449 34480 8483
rect 34428 8440 34480 8449
rect 34888 8440 34940 8492
rect 39212 8508 39264 8560
rect 39396 8508 39448 8560
rect 41604 8508 41656 8560
rect 57336 8551 57388 8560
rect 57336 8517 57345 8551
rect 57345 8517 57379 8551
rect 57379 8517 57388 8551
rect 57336 8508 57388 8517
rect 58256 8585 58265 8619
rect 58265 8585 58299 8619
rect 58299 8585 58308 8619
rect 58256 8576 58308 8585
rect 35532 8372 35584 8424
rect 29184 8347 29236 8356
rect 29184 8313 29193 8347
rect 29193 8313 29227 8347
rect 29227 8313 29236 8347
rect 29184 8304 29236 8313
rect 26792 8236 26844 8288
rect 28356 8279 28408 8288
rect 28356 8245 28365 8279
rect 28365 8245 28399 8279
rect 28399 8245 28408 8279
rect 28356 8236 28408 8245
rect 33416 8304 33468 8356
rect 37740 8440 37792 8492
rect 38108 8440 38160 8492
rect 37464 8372 37516 8424
rect 38660 8483 38712 8492
rect 38660 8449 38669 8483
rect 38669 8449 38703 8483
rect 38703 8449 38712 8483
rect 38660 8440 38712 8449
rect 40132 8440 40184 8492
rect 40316 8440 40368 8492
rect 56232 8483 56284 8492
rect 39212 8372 39264 8424
rect 31392 8236 31444 8288
rect 32312 8236 32364 8288
rect 38936 8304 38988 8356
rect 37648 8279 37700 8288
rect 37648 8245 37657 8279
rect 37657 8245 37691 8279
rect 37691 8245 37700 8279
rect 37648 8236 37700 8245
rect 38108 8236 38160 8288
rect 40500 8372 40552 8424
rect 56232 8449 56241 8483
rect 56241 8449 56275 8483
rect 56275 8449 56284 8483
rect 56232 8440 56284 8449
rect 57520 8440 57572 8492
rect 58348 8483 58400 8492
rect 58348 8449 58357 8483
rect 58357 8449 58391 8483
rect 58391 8449 58400 8483
rect 58348 8440 58400 8449
rect 58532 8372 58584 8424
rect 58072 8347 58124 8356
rect 58072 8313 58081 8347
rect 58081 8313 58115 8347
rect 58115 8313 58124 8347
rect 58072 8304 58124 8313
rect 56140 8236 56192 8288
rect 57152 8236 57204 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 12256 8032 12308 8084
rect 16948 8032 17000 8084
rect 17132 8075 17184 8084
rect 17132 8041 17141 8075
rect 17141 8041 17175 8075
rect 17175 8041 17184 8075
rect 17132 8032 17184 8041
rect 17408 8032 17460 8084
rect 11152 7964 11204 8016
rect 16856 7964 16908 8016
rect 19156 7964 19208 8016
rect 2688 7896 2740 7948
rect 11796 7828 11848 7880
rect 19432 7896 19484 7948
rect 20720 8032 20772 8084
rect 21456 8032 21508 8084
rect 32036 8032 32088 8084
rect 32128 8032 32180 8084
rect 36636 8032 36688 8084
rect 38016 8032 38068 8084
rect 38752 8032 38804 8084
rect 38936 8032 38988 8084
rect 40132 8075 40184 8084
rect 40132 8041 40141 8075
rect 40141 8041 40175 8075
rect 40175 8041 40184 8075
rect 40132 8032 40184 8041
rect 27160 7964 27212 8016
rect 27528 7964 27580 8016
rect 1860 7803 1912 7812
rect 1860 7769 1869 7803
rect 1869 7769 1903 7803
rect 1903 7769 1912 7803
rect 1860 7760 1912 7769
rect 12164 7760 12216 7812
rect 24676 7828 24728 7880
rect 30472 7896 30524 7948
rect 31024 7939 31076 7948
rect 31024 7905 31033 7939
rect 31033 7905 31067 7939
rect 31067 7905 31076 7939
rect 31024 7896 31076 7905
rect 31208 7939 31260 7948
rect 31208 7905 31217 7939
rect 31217 7905 31251 7939
rect 31251 7905 31260 7939
rect 31208 7896 31260 7905
rect 31484 7896 31536 7948
rect 32128 7939 32180 7948
rect 30748 7828 30800 7880
rect 30840 7828 30892 7880
rect 19616 7760 19668 7812
rect 19984 7760 20036 7812
rect 20352 7760 20404 7812
rect 20536 7760 20588 7812
rect 23664 7803 23716 7812
rect 23664 7769 23673 7803
rect 23673 7769 23707 7803
rect 23707 7769 23716 7803
rect 23664 7760 23716 7769
rect 18236 7692 18288 7744
rect 18328 7692 18380 7744
rect 20904 7735 20956 7744
rect 20904 7701 20913 7735
rect 20913 7701 20947 7735
rect 20947 7701 20956 7735
rect 20904 7692 20956 7701
rect 24860 7692 24912 7744
rect 25780 7760 25832 7812
rect 26424 7760 26476 7812
rect 28724 7760 28776 7812
rect 31576 7828 31628 7880
rect 31760 7871 31812 7880
rect 31760 7837 31769 7871
rect 31769 7837 31803 7871
rect 31803 7837 31812 7871
rect 32128 7905 32137 7939
rect 32137 7905 32171 7939
rect 32171 7905 32180 7939
rect 32128 7896 32180 7905
rect 32404 7896 32456 7948
rect 37280 7964 37332 8016
rect 33324 7896 33376 7948
rect 31760 7828 31812 7837
rect 34152 7896 34204 7948
rect 35348 7896 35400 7948
rect 36084 7896 36136 7948
rect 38200 7896 38252 7948
rect 38384 7896 38436 7948
rect 38844 7896 38896 7948
rect 39764 7896 39816 7948
rect 26148 7692 26200 7744
rect 28080 7692 28132 7744
rect 29460 7692 29512 7744
rect 33600 7760 33652 7812
rect 34980 7760 35032 7812
rect 37372 7828 37424 7880
rect 37740 7828 37792 7880
rect 38108 7828 38160 7880
rect 55312 7828 55364 7880
rect 57244 8032 57296 8084
rect 56876 7939 56928 7948
rect 39764 7760 39816 7812
rect 40132 7760 40184 7812
rect 50160 7760 50212 7812
rect 56140 7803 56192 7812
rect 56140 7769 56149 7803
rect 56149 7769 56183 7803
rect 56183 7769 56192 7803
rect 56140 7760 56192 7769
rect 56416 7871 56468 7880
rect 56416 7837 56425 7871
rect 56425 7837 56459 7871
rect 56459 7837 56468 7871
rect 56876 7905 56885 7939
rect 56885 7905 56919 7939
rect 56919 7905 56928 7939
rect 56876 7896 56928 7905
rect 56416 7828 56468 7837
rect 31668 7692 31720 7744
rect 36912 7692 36964 7744
rect 38016 7692 38068 7744
rect 56508 7692 56560 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 11796 7531 11848 7540
rect 11796 7497 11805 7531
rect 11805 7497 11839 7531
rect 11839 7497 11848 7531
rect 11796 7488 11848 7497
rect 13268 7531 13320 7540
rect 13268 7497 13277 7531
rect 13277 7497 13311 7531
rect 13311 7497 13320 7531
rect 13268 7488 13320 7497
rect 17960 7488 18012 7540
rect 19432 7488 19484 7540
rect 23756 7488 23808 7540
rect 24676 7531 24728 7540
rect 24676 7497 24685 7531
rect 24685 7497 24719 7531
rect 24719 7497 24728 7531
rect 24676 7488 24728 7497
rect 24768 7488 24820 7540
rect 30932 7488 30984 7540
rect 32404 7531 32456 7540
rect 32404 7497 32413 7531
rect 32413 7497 32447 7531
rect 32447 7497 32456 7531
rect 32404 7488 32456 7497
rect 34980 7531 35032 7540
rect 7656 7420 7708 7472
rect 11060 7352 11112 7404
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 11980 7352 12032 7361
rect 13268 7352 13320 7404
rect 20352 7395 20404 7404
rect 20352 7361 20361 7395
rect 20361 7361 20395 7395
rect 20395 7361 20404 7395
rect 20352 7352 20404 7361
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 12256 7327 12308 7336
rect 12256 7293 12265 7327
rect 12265 7293 12299 7327
rect 12299 7293 12308 7327
rect 12256 7284 12308 7293
rect 18512 7327 18564 7336
rect 18512 7293 18521 7327
rect 18521 7293 18555 7327
rect 18555 7293 18564 7327
rect 18512 7284 18564 7293
rect 13084 7259 13136 7268
rect 13084 7225 13093 7259
rect 13093 7225 13127 7259
rect 13127 7225 13136 7259
rect 13084 7216 13136 7225
rect 18696 7216 18748 7268
rect 18880 7216 18932 7268
rect 19800 7216 19852 7268
rect 19984 7259 20036 7268
rect 19984 7225 19993 7259
rect 19993 7225 20027 7259
rect 20027 7225 20036 7259
rect 19984 7216 20036 7225
rect 20904 7352 20956 7404
rect 29920 7463 29972 7472
rect 29920 7429 29929 7463
rect 29929 7429 29963 7463
rect 29963 7429 29972 7463
rect 29920 7420 29972 7429
rect 34980 7497 34989 7531
rect 34989 7497 35023 7531
rect 35023 7497 35032 7531
rect 34980 7488 35032 7497
rect 35164 7488 35216 7540
rect 36084 7488 36136 7540
rect 36912 7488 36964 7540
rect 25504 7352 25556 7404
rect 27160 7395 27212 7404
rect 27160 7361 27169 7395
rect 27169 7361 27203 7395
rect 27203 7361 27212 7395
rect 27160 7352 27212 7361
rect 28080 7352 28132 7404
rect 32312 7395 32364 7404
rect 32312 7361 32321 7395
rect 32321 7361 32355 7395
rect 32355 7361 32364 7395
rect 32312 7352 32364 7361
rect 32404 7352 32456 7404
rect 38660 7420 38712 7472
rect 33232 7352 33284 7404
rect 33416 7352 33468 7404
rect 34152 7395 34204 7404
rect 34152 7361 34161 7395
rect 34161 7361 34195 7395
rect 34195 7361 34204 7395
rect 34152 7352 34204 7361
rect 34612 7352 34664 7404
rect 20628 7327 20680 7336
rect 20628 7293 20637 7327
rect 20637 7293 20671 7327
rect 20671 7293 20680 7327
rect 20628 7284 20680 7293
rect 23204 7284 23256 7336
rect 28540 7284 28592 7336
rect 28632 7284 28684 7336
rect 33784 7284 33836 7336
rect 21364 7216 21416 7268
rect 20536 7148 20588 7200
rect 30840 7148 30892 7200
rect 31208 7148 31260 7200
rect 32588 7148 32640 7200
rect 34520 7284 34572 7336
rect 35440 7395 35492 7404
rect 35440 7361 35449 7395
rect 35449 7361 35483 7395
rect 35483 7361 35492 7395
rect 35440 7352 35492 7361
rect 35900 7352 35952 7404
rect 37556 7395 37608 7404
rect 37556 7361 37565 7395
rect 37565 7361 37599 7395
rect 37599 7361 37608 7395
rect 37556 7352 37608 7361
rect 38292 7352 38344 7404
rect 38752 7395 38804 7404
rect 38752 7361 38761 7395
rect 38761 7361 38795 7395
rect 38795 7361 38804 7395
rect 38752 7352 38804 7361
rect 35532 7284 35584 7336
rect 37740 7284 37792 7336
rect 38844 7327 38896 7336
rect 38844 7293 38853 7327
rect 38853 7293 38887 7327
rect 38887 7293 38896 7327
rect 38844 7284 38896 7293
rect 39212 7352 39264 7404
rect 39764 7463 39816 7472
rect 39764 7429 39773 7463
rect 39773 7429 39807 7463
rect 39807 7429 39816 7463
rect 39764 7420 39816 7429
rect 39672 7395 39724 7404
rect 39672 7361 39681 7395
rect 39681 7361 39715 7395
rect 39715 7361 39724 7395
rect 50160 7420 50212 7472
rect 39672 7352 39724 7361
rect 53564 7352 53616 7404
rect 56508 7352 56560 7404
rect 57244 7420 57296 7472
rect 57428 7420 57480 7472
rect 57612 7420 57664 7472
rect 57152 7352 57204 7404
rect 39948 7284 40000 7336
rect 56232 7284 56284 7336
rect 56416 7327 56468 7336
rect 56416 7293 56425 7327
rect 56425 7293 56459 7327
rect 56459 7293 56468 7327
rect 56416 7284 56468 7293
rect 34704 7216 34756 7268
rect 35164 7216 35216 7268
rect 39212 7259 39264 7268
rect 39212 7225 39221 7259
rect 39221 7225 39255 7259
rect 39255 7225 39264 7259
rect 39212 7216 39264 7225
rect 33876 7148 33928 7200
rect 34612 7191 34664 7200
rect 34612 7157 34621 7191
rect 34621 7157 34655 7191
rect 34655 7157 34664 7191
rect 34612 7148 34664 7157
rect 35256 7148 35308 7200
rect 35532 7148 35584 7200
rect 37188 7148 37240 7200
rect 38384 7191 38436 7200
rect 38384 7157 38393 7191
rect 38393 7157 38427 7191
rect 38427 7157 38436 7191
rect 38384 7148 38436 7157
rect 38660 7148 38712 7200
rect 38844 7148 38896 7200
rect 55404 7216 55456 7268
rect 47124 7148 47176 7200
rect 56600 7148 56652 7200
rect 57520 7148 57572 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 16856 6944 16908 6996
rect 20536 6944 20588 6996
rect 11060 6851 11112 6860
rect 11060 6817 11069 6851
rect 11069 6817 11103 6851
rect 11103 6817 11112 6851
rect 11060 6808 11112 6817
rect 11244 6851 11296 6860
rect 11244 6817 11253 6851
rect 11253 6817 11287 6851
rect 11287 6817 11296 6851
rect 11244 6808 11296 6817
rect 13544 6808 13596 6860
rect 13820 6808 13872 6860
rect 14004 6808 14056 6860
rect 19248 6876 19300 6928
rect 15292 6808 15344 6860
rect 18236 6808 18288 6860
rect 20168 6851 20220 6860
rect 20168 6817 20177 6851
rect 20177 6817 20211 6851
rect 20211 6817 20220 6851
rect 20168 6808 20220 6817
rect 20444 6876 20496 6928
rect 21364 6876 21416 6928
rect 22376 6919 22428 6928
rect 22376 6885 22385 6919
rect 22385 6885 22419 6919
rect 22419 6885 22428 6919
rect 22376 6876 22428 6885
rect 23572 6944 23624 6996
rect 26608 6944 26660 6996
rect 26792 6944 26844 6996
rect 38384 6944 38436 6996
rect 38660 6944 38712 6996
rect 47124 6944 47176 6996
rect 22836 6808 22888 6860
rect 9404 6783 9456 6792
rect 1860 6715 1912 6724
rect 1860 6681 1869 6715
rect 1869 6681 1903 6715
rect 1903 6681 1912 6715
rect 1860 6672 1912 6681
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 13268 6783 13320 6792
rect 11520 6740 11572 6749
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 9956 6672 10008 6724
rect 10140 6715 10192 6724
rect 10140 6681 10149 6715
rect 10149 6681 10183 6715
rect 10183 6681 10192 6715
rect 10140 6672 10192 6681
rect 11060 6672 11112 6724
rect 22100 6740 22152 6792
rect 20076 6672 20128 6724
rect 22560 6715 22612 6724
rect 22560 6681 22569 6715
rect 22569 6681 22603 6715
rect 22603 6681 22612 6715
rect 22560 6672 22612 6681
rect 17776 6604 17828 6656
rect 19984 6604 20036 6656
rect 22376 6604 22428 6656
rect 23020 6740 23072 6792
rect 23940 6876 23992 6928
rect 24032 6876 24084 6928
rect 24584 6851 24636 6860
rect 24584 6817 24593 6851
rect 24593 6817 24627 6851
rect 24627 6817 24636 6851
rect 24584 6808 24636 6817
rect 27620 6808 27672 6860
rect 28172 6808 28224 6860
rect 25136 6783 25188 6792
rect 25136 6749 25145 6783
rect 25145 6749 25179 6783
rect 25179 6749 25188 6783
rect 25136 6740 25188 6749
rect 28080 6740 28132 6792
rect 28632 6783 28684 6792
rect 28632 6749 28641 6783
rect 28641 6749 28675 6783
rect 28675 6749 28684 6783
rect 28632 6740 28684 6749
rect 29184 6808 29236 6860
rect 31484 6851 31536 6860
rect 31484 6817 31493 6851
rect 31493 6817 31527 6851
rect 31527 6817 31536 6851
rect 31484 6808 31536 6817
rect 31668 6808 31720 6860
rect 35900 6876 35952 6928
rect 37372 6876 37424 6928
rect 37556 6876 37608 6928
rect 39672 6876 39724 6928
rect 35440 6808 35492 6860
rect 36176 6808 36228 6860
rect 37188 6851 37240 6860
rect 37188 6817 37197 6851
rect 37197 6817 37231 6851
rect 37231 6817 37240 6851
rect 37188 6808 37240 6817
rect 37832 6851 37884 6860
rect 37832 6817 37841 6851
rect 37841 6817 37875 6851
rect 37875 6817 37884 6851
rect 37832 6808 37884 6817
rect 38016 6808 38068 6860
rect 39028 6851 39080 6860
rect 30380 6740 30432 6792
rect 30564 6740 30616 6792
rect 31208 6783 31260 6792
rect 24676 6672 24728 6724
rect 24584 6604 24636 6656
rect 25596 6672 25648 6724
rect 27160 6672 27212 6724
rect 31208 6749 31217 6783
rect 31217 6749 31251 6783
rect 31251 6749 31260 6783
rect 31208 6740 31260 6749
rect 31300 6749 31310 6758
rect 31310 6749 31344 6758
rect 31344 6749 31352 6758
rect 31300 6706 31352 6749
rect 32864 6783 32916 6792
rect 32864 6749 32873 6783
rect 32873 6749 32907 6783
rect 32907 6749 32916 6783
rect 32864 6740 32916 6749
rect 35624 6783 35676 6792
rect 35624 6749 35633 6783
rect 35633 6749 35667 6783
rect 35667 6749 35676 6783
rect 35624 6740 35676 6749
rect 24952 6647 25004 6656
rect 24952 6613 24961 6647
rect 24961 6613 24995 6647
rect 24995 6613 25004 6647
rect 24952 6604 25004 6613
rect 25136 6604 25188 6656
rect 31576 6672 31628 6724
rect 33968 6715 34020 6724
rect 33968 6681 33977 6715
rect 33977 6681 34011 6715
rect 34011 6681 34020 6715
rect 33968 6672 34020 6681
rect 27620 6604 27672 6656
rect 28908 6604 28960 6656
rect 31760 6604 31812 6656
rect 33048 6647 33100 6656
rect 33048 6613 33057 6647
rect 33057 6613 33091 6647
rect 33091 6613 33100 6647
rect 33048 6604 33100 6613
rect 34612 6672 34664 6724
rect 34704 6604 34756 6656
rect 36544 6647 36596 6656
rect 36544 6613 36553 6647
rect 36553 6613 36587 6647
rect 36587 6613 36596 6647
rect 36544 6604 36596 6613
rect 36820 6604 36872 6656
rect 37648 6672 37700 6724
rect 38292 6783 38344 6792
rect 38292 6749 38301 6783
rect 38301 6749 38335 6783
rect 38335 6749 38344 6783
rect 39028 6817 39037 6851
rect 39037 6817 39071 6851
rect 39071 6817 39080 6851
rect 39028 6808 39080 6817
rect 38292 6740 38344 6749
rect 38752 6740 38804 6792
rect 37004 6647 37056 6656
rect 37004 6613 37013 6647
rect 37013 6613 37047 6647
rect 37047 6613 37056 6647
rect 37004 6604 37056 6613
rect 38476 6604 38528 6656
rect 56692 6740 56744 6792
rect 57520 6740 57572 6792
rect 57520 6604 57572 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 11520 6400 11572 6452
rect 12256 6400 12308 6452
rect 17776 6400 17828 6452
rect 17868 6443 17920 6452
rect 17868 6409 17877 6443
rect 17877 6409 17911 6443
rect 17911 6409 17920 6443
rect 17868 6400 17920 6409
rect 11612 6332 11664 6384
rect 13268 6332 13320 6384
rect 18236 6375 18288 6384
rect 18236 6341 18245 6375
rect 18245 6341 18279 6375
rect 18279 6341 18288 6375
rect 18236 6332 18288 6341
rect 18512 6332 18564 6384
rect 9496 6264 9548 6316
rect 16948 6264 17000 6316
rect 19524 6400 19576 6452
rect 20076 6400 20128 6452
rect 23940 6400 23992 6452
rect 24768 6400 24820 6452
rect 24952 6443 25004 6452
rect 24952 6409 24961 6443
rect 24961 6409 24995 6443
rect 24995 6409 25004 6443
rect 24952 6400 25004 6409
rect 25320 6400 25372 6452
rect 25780 6443 25832 6452
rect 25780 6409 25789 6443
rect 25789 6409 25823 6443
rect 25823 6409 25832 6443
rect 25780 6400 25832 6409
rect 26148 6400 26200 6452
rect 27160 6443 27212 6452
rect 27160 6409 27169 6443
rect 27169 6409 27203 6443
rect 27203 6409 27212 6443
rect 27160 6400 27212 6409
rect 28264 6400 28316 6452
rect 19248 6332 19300 6384
rect 19984 6332 20036 6384
rect 1768 6239 1820 6248
rect 1768 6205 1777 6239
rect 1777 6205 1811 6239
rect 1811 6205 1820 6239
rect 1768 6196 1820 6205
rect 11060 6196 11112 6248
rect 12348 6196 12400 6248
rect 8852 6128 8904 6180
rect 11520 6128 11572 6180
rect 10140 6060 10192 6112
rect 15568 6196 15620 6248
rect 15660 6196 15712 6248
rect 18328 6239 18380 6248
rect 18328 6205 18337 6239
rect 18337 6205 18371 6239
rect 18371 6205 18380 6239
rect 18328 6196 18380 6205
rect 18604 6196 18656 6248
rect 14556 6128 14608 6180
rect 16120 6171 16172 6180
rect 16120 6137 16129 6171
rect 16129 6137 16163 6171
rect 16163 6137 16172 6171
rect 16120 6128 16172 6137
rect 19156 6264 19208 6316
rect 21640 6264 21692 6316
rect 22928 6264 22980 6316
rect 23664 6307 23716 6316
rect 23664 6273 23673 6307
rect 23673 6273 23707 6307
rect 23707 6273 23716 6307
rect 23664 6264 23716 6273
rect 25044 6332 25096 6384
rect 25596 6332 25648 6384
rect 29000 6400 29052 6452
rect 30012 6443 30064 6452
rect 30012 6409 30021 6443
rect 30021 6409 30055 6443
rect 30055 6409 30064 6443
rect 30012 6400 30064 6409
rect 31852 6400 31904 6452
rect 24860 6307 24912 6316
rect 24860 6273 24869 6307
rect 24869 6273 24903 6307
rect 24903 6273 24912 6307
rect 24860 6264 24912 6273
rect 25504 6264 25556 6316
rect 26056 6264 26108 6316
rect 27528 6264 27580 6316
rect 19064 6128 19116 6180
rect 22560 6128 22612 6180
rect 22836 6196 22888 6248
rect 23848 6128 23900 6180
rect 25688 6196 25740 6248
rect 25964 6196 26016 6248
rect 26424 6239 26476 6248
rect 26424 6205 26433 6239
rect 26433 6205 26467 6239
rect 26467 6205 26476 6239
rect 26424 6196 26476 6205
rect 27620 6239 27672 6248
rect 27620 6205 27629 6239
rect 27629 6205 27663 6239
rect 27663 6205 27672 6239
rect 27620 6196 27672 6205
rect 28080 6264 28132 6316
rect 28908 6239 28960 6248
rect 28908 6205 28917 6239
rect 28917 6205 28951 6239
rect 28951 6205 28960 6239
rect 28908 6196 28960 6205
rect 31208 6264 31260 6316
rect 31944 6264 31996 6316
rect 32680 6264 32732 6316
rect 33048 6375 33100 6384
rect 33048 6341 33082 6375
rect 33082 6341 33100 6375
rect 33048 6332 33100 6341
rect 35624 6332 35676 6384
rect 35808 6332 35860 6384
rect 57612 6400 57664 6452
rect 34796 6264 34848 6316
rect 37372 6332 37424 6384
rect 30932 6196 30984 6248
rect 57244 6264 57296 6316
rect 57520 6307 57572 6316
rect 57520 6273 57529 6307
rect 57529 6273 57563 6307
rect 57563 6273 57572 6307
rect 57520 6264 57572 6273
rect 38568 6196 38620 6248
rect 30104 6128 30156 6180
rect 31300 6128 31352 6180
rect 33784 6128 33836 6180
rect 37188 6128 37240 6180
rect 24032 6060 24084 6112
rect 24492 6103 24544 6112
rect 24492 6069 24501 6103
rect 24501 6069 24535 6103
rect 24535 6069 24544 6103
rect 24492 6060 24544 6069
rect 24584 6060 24636 6112
rect 33140 6060 33192 6112
rect 33416 6060 33468 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 13084 5856 13136 5908
rect 16120 5856 16172 5908
rect 12992 5788 13044 5840
rect 13544 5788 13596 5840
rect 22836 5856 22888 5908
rect 26332 5856 26384 5908
rect 31116 5856 31168 5908
rect 32864 5899 32916 5908
rect 32864 5865 32873 5899
rect 32873 5865 32907 5899
rect 32907 5865 32916 5899
rect 32864 5856 32916 5865
rect 18972 5788 19024 5840
rect 23572 5788 23624 5840
rect 23664 5788 23716 5840
rect 28172 5788 28224 5840
rect 29000 5788 29052 5840
rect 36820 5856 36872 5908
rect 18604 5720 18656 5772
rect 19432 5763 19484 5772
rect 19432 5729 19441 5763
rect 19441 5729 19475 5763
rect 19475 5729 19484 5763
rect 19432 5720 19484 5729
rect 17776 5652 17828 5704
rect 22008 5720 22060 5772
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 24676 5720 24728 5772
rect 25596 5763 25648 5772
rect 11704 5584 11756 5636
rect 12532 5584 12584 5636
rect 13360 5584 13412 5636
rect 14188 5584 14240 5636
rect 16580 5584 16632 5636
rect 22284 5652 22336 5704
rect 22652 5695 22704 5704
rect 22652 5661 22661 5695
rect 22661 5661 22695 5695
rect 22695 5661 22704 5695
rect 22652 5652 22704 5661
rect 24032 5695 24084 5704
rect 18972 5584 19024 5636
rect 21364 5584 21416 5636
rect 21824 5584 21876 5636
rect 22376 5584 22428 5636
rect 23020 5627 23072 5636
rect 14464 5559 14516 5568
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 14464 5516 14516 5525
rect 17132 5516 17184 5568
rect 18512 5559 18564 5568
rect 18512 5525 18521 5559
rect 18521 5525 18555 5559
rect 18555 5525 18564 5559
rect 18512 5516 18564 5525
rect 18604 5559 18656 5568
rect 18604 5525 18613 5559
rect 18613 5525 18647 5559
rect 18647 5525 18656 5559
rect 18604 5516 18656 5525
rect 18880 5516 18932 5568
rect 20260 5516 20312 5568
rect 20812 5559 20864 5568
rect 20812 5525 20821 5559
rect 20821 5525 20855 5559
rect 20855 5525 20864 5559
rect 20812 5516 20864 5525
rect 22744 5559 22796 5568
rect 22744 5525 22753 5559
rect 22753 5525 22787 5559
rect 22787 5525 22796 5559
rect 22744 5516 22796 5525
rect 23020 5593 23029 5627
rect 23029 5593 23063 5627
rect 23063 5593 23072 5627
rect 23020 5584 23072 5593
rect 23664 5627 23716 5636
rect 23664 5593 23673 5627
rect 23673 5593 23707 5627
rect 23707 5593 23716 5627
rect 23664 5584 23716 5593
rect 24032 5661 24041 5695
rect 24041 5661 24075 5695
rect 24075 5661 24084 5695
rect 24032 5652 24084 5661
rect 24400 5584 24452 5636
rect 24584 5627 24636 5636
rect 24584 5593 24593 5627
rect 24593 5593 24627 5627
rect 24627 5593 24636 5627
rect 24584 5584 24636 5593
rect 25228 5652 25280 5704
rect 25596 5729 25605 5763
rect 25605 5729 25639 5763
rect 25639 5729 25648 5763
rect 25596 5720 25648 5729
rect 25780 5695 25832 5704
rect 25780 5661 25789 5695
rect 25789 5661 25823 5695
rect 25823 5661 25832 5695
rect 25780 5652 25832 5661
rect 25964 5652 26016 5704
rect 27620 5652 27672 5704
rect 28632 5720 28684 5772
rect 34612 5788 34664 5840
rect 33784 5720 33836 5772
rect 34520 5720 34572 5772
rect 35348 5720 35400 5772
rect 28356 5695 28408 5704
rect 28356 5661 28370 5695
rect 28370 5661 28404 5695
rect 28404 5661 28408 5695
rect 28356 5652 28408 5661
rect 30288 5695 30340 5704
rect 30288 5661 30297 5695
rect 30297 5661 30331 5695
rect 30331 5661 30340 5695
rect 30288 5652 30340 5661
rect 30472 5695 30524 5704
rect 30472 5661 30481 5695
rect 30481 5661 30515 5695
rect 30515 5661 30524 5695
rect 30472 5652 30524 5661
rect 31668 5652 31720 5704
rect 32128 5652 32180 5704
rect 33232 5695 33284 5704
rect 33232 5661 33241 5695
rect 33241 5661 33275 5695
rect 33275 5661 33284 5695
rect 33232 5652 33284 5661
rect 25136 5627 25188 5636
rect 25136 5593 25145 5627
rect 25145 5593 25179 5627
rect 25179 5593 25188 5627
rect 25136 5584 25188 5593
rect 23940 5516 23992 5568
rect 25872 5559 25924 5568
rect 25872 5525 25881 5559
rect 25881 5525 25915 5559
rect 25915 5525 25924 5559
rect 25872 5516 25924 5525
rect 28908 5584 28960 5636
rect 33416 5584 33468 5636
rect 33600 5584 33652 5636
rect 35532 5584 35584 5636
rect 35900 5627 35952 5636
rect 35900 5593 35909 5627
rect 35909 5593 35943 5627
rect 35943 5593 35952 5627
rect 35900 5584 35952 5593
rect 36728 5627 36780 5636
rect 36728 5593 36762 5627
rect 36762 5593 36780 5627
rect 36728 5584 36780 5593
rect 28356 5516 28408 5568
rect 28816 5516 28868 5568
rect 30656 5559 30708 5568
rect 30656 5525 30665 5559
rect 30665 5525 30699 5559
rect 30699 5525 30708 5559
rect 30656 5516 30708 5525
rect 32680 5516 32732 5568
rect 34520 5516 34572 5568
rect 34796 5516 34848 5568
rect 57520 5652 57572 5704
rect 57980 5695 58032 5704
rect 57980 5661 57989 5695
rect 57989 5661 58023 5695
rect 58023 5661 58032 5695
rect 57980 5652 58032 5661
rect 57244 5627 57296 5636
rect 57244 5593 57253 5627
rect 57253 5593 57287 5627
rect 57287 5593 57296 5627
rect 57244 5584 57296 5593
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 12348 5355 12400 5364
rect 12348 5321 12357 5355
rect 12357 5321 12391 5355
rect 12391 5321 12400 5355
rect 12348 5312 12400 5321
rect 18328 5312 18380 5364
rect 11152 5287 11204 5296
rect 11152 5253 11161 5287
rect 11161 5253 11195 5287
rect 11195 5253 11204 5287
rect 11152 5244 11204 5253
rect 13820 5287 13872 5296
rect 13820 5253 13829 5287
rect 13829 5253 13863 5287
rect 13863 5253 13872 5287
rect 13820 5244 13872 5253
rect 29000 5312 29052 5364
rect 29460 5355 29512 5364
rect 29460 5321 29469 5355
rect 29469 5321 29503 5355
rect 29503 5321 29512 5355
rect 29460 5312 29512 5321
rect 30472 5312 30524 5364
rect 31944 5312 31996 5364
rect 32772 5312 32824 5364
rect 34060 5312 34112 5364
rect 34704 5312 34756 5364
rect 36728 5355 36780 5364
rect 9864 5176 9916 5228
rect 10048 5176 10100 5228
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 13636 5219 13688 5228
rect 1768 5151 1820 5160
rect 1768 5117 1777 5151
rect 1777 5117 1811 5151
rect 1811 5117 1820 5151
rect 1768 5108 1820 5117
rect 7932 5108 7984 5160
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 17684 5176 17736 5228
rect 10416 5083 10468 5092
rect 10416 5049 10425 5083
rect 10425 5049 10459 5083
rect 10459 5049 10468 5083
rect 10416 5040 10468 5049
rect 13268 5108 13320 5160
rect 16120 5108 16172 5160
rect 10692 5040 10744 5092
rect 12808 5040 12860 5092
rect 18328 5040 18380 5092
rect 18512 5108 18564 5160
rect 20812 5176 20864 5228
rect 20996 5219 21048 5228
rect 20996 5185 21005 5219
rect 21005 5185 21039 5219
rect 21039 5185 21048 5219
rect 20996 5176 21048 5185
rect 23112 5244 23164 5296
rect 25504 5244 25556 5296
rect 19064 5151 19116 5160
rect 19064 5117 19073 5151
rect 19073 5117 19107 5151
rect 19107 5117 19116 5151
rect 19064 5108 19116 5117
rect 21640 5108 21692 5160
rect 22008 5108 22060 5160
rect 23940 5176 23992 5228
rect 24492 5176 24544 5228
rect 25872 5244 25924 5296
rect 36728 5321 36737 5355
rect 36737 5321 36771 5355
rect 36771 5321 36780 5355
rect 36728 5312 36780 5321
rect 36820 5312 36872 5364
rect 39856 5355 39908 5364
rect 39856 5321 39865 5355
rect 39865 5321 39899 5355
rect 39899 5321 39908 5355
rect 39856 5312 39908 5321
rect 40960 5312 41012 5364
rect 42156 5312 42208 5364
rect 28080 5219 28132 5228
rect 28080 5185 28089 5219
rect 28089 5185 28123 5219
rect 28123 5185 28132 5219
rect 28080 5176 28132 5185
rect 28356 5219 28408 5228
rect 28356 5185 28365 5219
rect 28365 5185 28399 5219
rect 28399 5185 28408 5219
rect 28356 5176 28408 5185
rect 23296 5108 23348 5160
rect 26516 5108 26568 5160
rect 26608 5108 26660 5160
rect 30564 5176 30616 5228
rect 32404 5176 32456 5228
rect 33048 5176 33100 5228
rect 33692 5176 33744 5228
rect 34612 5219 34664 5228
rect 34612 5185 34621 5219
rect 34621 5185 34655 5219
rect 34655 5185 34664 5219
rect 34612 5176 34664 5185
rect 35532 5244 35584 5296
rect 35992 5176 36044 5228
rect 36544 5219 36596 5228
rect 36544 5185 36553 5219
rect 36553 5185 36587 5219
rect 36587 5185 36596 5219
rect 36544 5176 36596 5185
rect 37372 5244 37424 5296
rect 38568 5176 38620 5228
rect 38660 5176 38712 5228
rect 39120 5176 39172 5228
rect 40040 5176 40092 5228
rect 43168 5244 43220 5296
rect 55588 5312 55640 5364
rect 56140 5312 56192 5364
rect 43812 5219 43864 5228
rect 43812 5185 43821 5219
rect 43821 5185 43855 5219
rect 43855 5185 43864 5219
rect 43812 5176 43864 5185
rect 43996 5176 44048 5228
rect 56600 5176 56652 5228
rect 58072 5219 58124 5228
rect 58072 5185 58081 5219
rect 58081 5185 58115 5219
rect 58115 5185 58124 5219
rect 58072 5176 58124 5185
rect 29552 5108 29604 5160
rect 31116 5108 31168 5160
rect 32680 5108 32732 5160
rect 32864 5108 32916 5160
rect 33784 5108 33836 5160
rect 14740 5015 14792 5024
rect 14740 4981 14749 5015
rect 14749 4981 14783 5015
rect 14783 4981 14792 5015
rect 14740 4972 14792 4981
rect 17960 4972 18012 5024
rect 18052 4972 18104 5024
rect 22928 4972 22980 5024
rect 25044 5040 25096 5092
rect 29092 5040 29144 5092
rect 37004 5108 37056 5160
rect 37096 5108 37148 5160
rect 37280 5040 37332 5092
rect 39304 5040 39356 5092
rect 42064 5040 42116 5092
rect 24768 5015 24820 5024
rect 24768 4981 24777 5015
rect 24777 4981 24811 5015
rect 24811 4981 24820 5015
rect 24768 4972 24820 4981
rect 27252 4972 27304 5024
rect 32312 5015 32364 5024
rect 32312 4981 32321 5015
rect 32321 4981 32355 5015
rect 32355 4981 32364 5015
rect 32312 4972 32364 4981
rect 44732 5015 44784 5024
rect 44732 4981 44741 5015
rect 44741 4981 44775 5015
rect 44775 4981 44784 5015
rect 44732 4972 44784 4981
rect 58256 5015 58308 5024
rect 58256 4981 58265 5015
rect 58265 4981 58299 5015
rect 58299 4981 58308 5015
rect 58256 4972 58308 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 9956 4768 10008 4820
rect 6920 4700 6972 4752
rect 10692 4700 10744 4752
rect 11244 4768 11296 4820
rect 11612 4811 11664 4820
rect 11612 4777 11621 4811
rect 11621 4777 11655 4811
rect 11655 4777 11664 4811
rect 11612 4768 11664 4777
rect 11980 4768 12032 4820
rect 18604 4768 18656 4820
rect 20996 4811 21048 4820
rect 20996 4777 21005 4811
rect 21005 4777 21039 4811
rect 21039 4777 21048 4811
rect 20996 4768 21048 4777
rect 23020 4768 23072 4820
rect 16120 4700 16172 4752
rect 22284 4700 22336 4752
rect 30564 4768 30616 4820
rect 33600 4768 33652 4820
rect 41696 4811 41748 4820
rect 41696 4777 41705 4811
rect 41705 4777 41739 4811
rect 41739 4777 41748 4811
rect 41696 4768 41748 4777
rect 43628 4768 43680 4820
rect 47584 4811 47636 4820
rect 47584 4777 47593 4811
rect 47593 4777 47627 4811
rect 47627 4777 47636 4811
rect 47584 4768 47636 4777
rect 55404 4768 55456 4820
rect 8300 4564 8352 4616
rect 9588 4564 9640 4616
rect 11612 4632 11664 4684
rect 18052 4632 18104 4684
rect 1860 4539 1912 4548
rect 1860 4505 1869 4539
rect 1869 4505 1903 4539
rect 1903 4505 1912 4539
rect 1860 4496 1912 4505
rect 7288 4496 7340 4548
rect 8576 4496 8628 4548
rect 7564 4471 7616 4480
rect 7564 4437 7573 4471
rect 7573 4437 7607 4471
rect 7607 4437 7616 4471
rect 7564 4428 7616 4437
rect 8760 4428 8812 4480
rect 10324 4496 10376 4548
rect 11152 4564 11204 4616
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 12348 4564 12400 4616
rect 19064 4632 19116 4684
rect 20628 4632 20680 4684
rect 19800 4564 19852 4616
rect 22192 4632 22244 4684
rect 21272 4564 21324 4616
rect 24768 4700 24820 4752
rect 29092 4700 29144 4752
rect 22928 4675 22980 4684
rect 22928 4641 22937 4675
rect 22937 4641 22971 4675
rect 22971 4641 22980 4675
rect 22928 4632 22980 4641
rect 25044 4675 25096 4684
rect 12440 4496 12492 4548
rect 14924 4496 14976 4548
rect 15844 4496 15896 4548
rect 16948 4496 17000 4548
rect 22836 4607 22888 4616
rect 22836 4573 22845 4607
rect 22845 4573 22879 4607
rect 22879 4573 22888 4607
rect 22836 4564 22888 4573
rect 21732 4496 21784 4548
rect 25044 4641 25053 4675
rect 25053 4641 25087 4675
rect 25087 4641 25096 4675
rect 25044 4632 25096 4641
rect 24952 4607 25004 4616
rect 24952 4573 24961 4607
rect 24961 4573 24995 4607
rect 24995 4573 25004 4607
rect 24952 4564 25004 4573
rect 26424 4632 26476 4684
rect 26884 4632 26936 4684
rect 32128 4675 32180 4684
rect 27436 4564 27488 4616
rect 27620 4564 27672 4616
rect 28908 4564 28960 4616
rect 30104 4564 30156 4616
rect 10232 4428 10284 4480
rect 11244 4428 11296 4480
rect 12348 4428 12400 4480
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 18512 4471 18564 4480
rect 18512 4437 18521 4471
rect 18521 4437 18555 4471
rect 18555 4437 18564 4471
rect 18512 4428 18564 4437
rect 19340 4428 19392 4480
rect 19984 4471 20036 4480
rect 19984 4437 19993 4471
rect 19993 4437 20027 4471
rect 20027 4437 20036 4471
rect 19984 4428 20036 4437
rect 20628 4428 20680 4480
rect 25136 4496 25188 4548
rect 28448 4496 28500 4548
rect 28540 4496 28592 4548
rect 30012 4496 30064 4548
rect 24584 4471 24636 4480
rect 24584 4437 24593 4471
rect 24593 4437 24627 4471
rect 24627 4437 24636 4471
rect 24584 4428 24636 4437
rect 28264 4428 28316 4480
rect 29000 4428 29052 4480
rect 29092 4471 29144 4480
rect 29092 4437 29101 4471
rect 29101 4437 29135 4471
rect 29135 4437 29144 4471
rect 30932 4564 30984 4616
rect 30656 4496 30708 4548
rect 32128 4641 32137 4675
rect 32137 4641 32171 4675
rect 32171 4641 32180 4675
rect 32128 4632 32180 4641
rect 32312 4607 32364 4616
rect 32312 4573 32321 4607
rect 32321 4573 32355 4607
rect 32355 4573 32364 4607
rect 32312 4564 32364 4573
rect 39580 4700 39632 4752
rect 43260 4743 43312 4752
rect 43260 4709 43269 4743
rect 43269 4709 43303 4743
rect 43303 4709 43312 4743
rect 43260 4700 43312 4709
rect 44180 4743 44232 4752
rect 44180 4709 44189 4743
rect 44189 4709 44223 4743
rect 44223 4709 44232 4743
rect 44180 4700 44232 4709
rect 45192 4700 45244 4752
rect 34428 4564 34480 4616
rect 34796 4564 34848 4616
rect 36176 4564 36228 4616
rect 37188 4607 37240 4616
rect 37188 4573 37197 4607
rect 37197 4573 37231 4607
rect 37231 4573 37240 4607
rect 37188 4564 37240 4573
rect 39488 4632 39540 4684
rect 45468 4632 45520 4684
rect 46848 4632 46900 4684
rect 56600 4632 56652 4684
rect 38568 4564 38620 4616
rect 39212 4564 39264 4616
rect 45928 4564 45980 4616
rect 32404 4496 32456 4548
rect 34612 4496 34664 4548
rect 37096 4496 37148 4548
rect 38936 4539 38988 4548
rect 38936 4505 38945 4539
rect 38945 4505 38979 4539
rect 38979 4505 38988 4539
rect 38936 4496 38988 4505
rect 29092 4428 29144 4437
rect 32312 4428 32364 4480
rect 35808 4428 35860 4480
rect 36084 4428 36136 4480
rect 38476 4428 38528 4480
rect 41420 4496 41472 4548
rect 42064 4496 42116 4548
rect 42892 4496 42944 4548
rect 42984 4496 43036 4548
rect 43168 4496 43220 4548
rect 44364 4496 44416 4548
rect 39120 4428 39172 4480
rect 45008 4428 45060 4480
rect 46572 4564 46624 4616
rect 47492 4564 47544 4616
rect 57980 4607 58032 4616
rect 57980 4573 57989 4607
rect 57989 4573 58023 4607
rect 58023 4573 58032 4607
rect 57980 4564 58032 4573
rect 58164 4607 58216 4616
rect 58164 4573 58173 4607
rect 58173 4573 58207 4607
rect 58207 4573 58216 4607
rect 58164 4564 58216 4573
rect 56600 4539 56652 4548
rect 56600 4505 56609 4539
rect 56609 4505 56643 4539
rect 56643 4505 56652 4539
rect 56600 4496 56652 4505
rect 45744 4428 45796 4480
rect 46204 4428 46256 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 7564 4224 7616 4276
rect 18512 4224 18564 4276
rect 7840 4156 7892 4208
rect 9496 4156 9548 4208
rect 8668 4088 8720 4140
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 10876 4156 10928 4208
rect 11336 4156 11388 4208
rect 10692 4131 10744 4140
rect 10692 4097 10701 4131
rect 10701 4097 10735 4131
rect 10735 4097 10744 4131
rect 10692 4088 10744 4097
rect 11152 4088 11204 4140
rect 12624 4156 12676 4208
rect 19524 4224 19576 4276
rect 19984 4224 20036 4276
rect 20536 4224 20588 4276
rect 22928 4224 22980 4276
rect 24584 4156 24636 4208
rect 25044 4224 25096 4276
rect 29552 4224 29604 4276
rect 30196 4224 30248 4276
rect 33048 4224 33100 4276
rect 58256 4224 58308 4276
rect 29092 4156 29144 4208
rect 30104 4156 30156 4208
rect 12348 4131 12400 4140
rect 12348 4097 12357 4131
rect 12357 4097 12391 4131
rect 12391 4097 12400 4131
rect 12348 4088 12400 4097
rect 13912 4088 13964 4140
rect 14740 4088 14792 4140
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 15660 4088 15712 4140
rect 16856 4131 16908 4140
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 7656 4020 7708 4072
rect 9588 4020 9640 4072
rect 9864 4020 9916 4072
rect 10508 4063 10560 4072
rect 10508 4029 10517 4063
rect 10517 4029 10551 4063
rect 10551 4029 10560 4063
rect 10508 4020 10560 4029
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 10968 4020 11020 4072
rect 11428 4020 11480 4072
rect 11612 4020 11664 4072
rect 12808 4020 12860 4072
rect 14096 4020 14148 4072
rect 16856 4097 16865 4131
rect 16865 4097 16899 4131
rect 16899 4097 16908 4131
rect 16856 4088 16908 4097
rect 17500 4088 17552 4140
rect 17868 4088 17920 4140
rect 19064 4131 19116 4140
rect 19064 4097 19073 4131
rect 19073 4097 19107 4131
rect 19107 4097 19116 4131
rect 19064 4088 19116 4097
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 20444 4088 20496 4140
rect 21088 4088 21140 4140
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 22284 4131 22336 4140
rect 22284 4097 22318 4131
rect 22318 4097 22336 4131
rect 23940 4131 23992 4140
rect 22284 4088 22336 4097
rect 23940 4097 23949 4131
rect 23949 4097 23983 4131
rect 23983 4097 23992 4131
rect 23940 4088 23992 4097
rect 9036 3884 9088 3936
rect 10140 3884 10192 3936
rect 13728 3952 13780 4004
rect 13820 3952 13872 4004
rect 14372 3952 14424 4004
rect 16396 3952 16448 4004
rect 16672 3952 16724 4004
rect 17316 4020 17368 4072
rect 18420 4020 18472 4072
rect 18696 4020 18748 4072
rect 20168 4063 20220 4072
rect 13084 3884 13136 3936
rect 13268 3884 13320 3936
rect 14096 3884 14148 3936
rect 17408 3884 17460 3936
rect 18696 3927 18748 3936
rect 18696 3893 18705 3927
rect 18705 3893 18739 3927
rect 18739 3893 18748 3927
rect 18696 3884 18748 3893
rect 20168 4029 20177 4063
rect 20177 4029 20211 4063
rect 20211 4029 20220 4063
rect 20168 4020 20220 4029
rect 20628 4020 20680 4072
rect 18972 3884 19024 3936
rect 19708 3927 19760 3936
rect 19708 3893 19717 3927
rect 19717 3893 19751 3927
rect 19751 3893 19760 3927
rect 19708 3884 19760 3893
rect 25504 4020 25556 4072
rect 26424 4088 26476 4140
rect 26884 4020 26936 4072
rect 26976 4020 27028 4072
rect 28540 4088 28592 4140
rect 28724 4088 28776 4140
rect 29736 4063 29788 4072
rect 29736 4029 29745 4063
rect 29745 4029 29779 4063
rect 29779 4029 29788 4063
rect 29736 4020 29788 4029
rect 30012 4088 30064 4140
rect 24952 3952 25004 4004
rect 31208 3952 31260 4004
rect 32036 4156 32088 4208
rect 33416 4156 33468 4208
rect 31760 4088 31812 4140
rect 32956 4088 33008 4140
rect 33600 4131 33652 4140
rect 33600 4097 33609 4131
rect 33609 4097 33643 4131
rect 33643 4097 33652 4131
rect 33600 4088 33652 4097
rect 36912 4156 36964 4208
rect 37188 4156 37240 4208
rect 35624 4088 35676 4140
rect 35716 4088 35768 4140
rect 23020 3884 23072 3936
rect 23204 3884 23256 3936
rect 25412 3884 25464 3936
rect 27160 3927 27212 3936
rect 27160 3893 27169 3927
rect 27169 3893 27203 3927
rect 27203 3893 27212 3927
rect 27160 3884 27212 3893
rect 28540 3884 28592 3936
rect 29276 3927 29328 3936
rect 29276 3893 29285 3927
rect 29285 3893 29319 3927
rect 29319 3893 29328 3927
rect 29276 3884 29328 3893
rect 30288 3884 30340 3936
rect 31668 3927 31720 3936
rect 31668 3893 31677 3927
rect 31677 3893 31711 3927
rect 31711 3893 31720 3927
rect 31668 3884 31720 3893
rect 33232 3884 33284 3936
rect 36268 4131 36320 4140
rect 36268 4097 36277 4131
rect 36277 4097 36311 4131
rect 36311 4097 36320 4131
rect 36268 4088 36320 4097
rect 37556 4088 37608 4140
rect 38568 4156 38620 4208
rect 38752 4156 38804 4208
rect 39948 4131 40000 4140
rect 36360 4020 36412 4072
rect 38200 4020 38252 4072
rect 38660 4020 38712 4072
rect 38844 4020 38896 4072
rect 39120 4020 39172 4072
rect 39948 4097 39957 4131
rect 39957 4097 39991 4131
rect 39991 4097 40000 4131
rect 39948 4088 40000 4097
rect 41512 4088 41564 4140
rect 42524 4088 42576 4140
rect 43260 4131 43312 4140
rect 43260 4097 43269 4131
rect 43269 4097 43303 4131
rect 43303 4097 43312 4131
rect 43260 4088 43312 4097
rect 40132 4020 40184 4072
rect 41788 4063 41840 4072
rect 41788 4029 41797 4063
rect 41797 4029 41831 4063
rect 41831 4029 41840 4063
rect 41788 4020 41840 4029
rect 43904 4088 43956 4140
rect 46204 4156 46256 4208
rect 46296 4156 46348 4208
rect 46848 4199 46900 4208
rect 45652 4131 45704 4140
rect 45652 4097 45661 4131
rect 45661 4097 45695 4131
rect 45695 4097 45704 4131
rect 45652 4088 45704 4097
rect 46848 4165 46857 4199
rect 46857 4165 46891 4199
rect 46891 4165 46900 4199
rect 46848 4156 46900 4165
rect 47032 4156 47084 4208
rect 43076 3952 43128 4004
rect 45192 4020 45244 4072
rect 46204 4020 46256 4072
rect 46388 3952 46440 4004
rect 55404 4131 55456 4140
rect 55404 4097 55413 4131
rect 55413 4097 55447 4131
rect 55447 4097 55456 4131
rect 55404 4088 55456 4097
rect 55588 4131 55640 4140
rect 55588 4097 55597 4131
rect 55597 4097 55631 4131
rect 55631 4097 55640 4131
rect 55588 4088 55640 4097
rect 47676 4020 47728 4072
rect 58072 4131 58124 4140
rect 58072 4097 58081 4131
rect 58081 4097 58115 4131
rect 58115 4097 58124 4131
rect 58072 4088 58124 4097
rect 53932 3952 53984 4004
rect 34336 3884 34388 3936
rect 36268 3884 36320 3936
rect 37188 3884 37240 3936
rect 37464 3884 37516 3936
rect 38660 3884 38712 3936
rect 40224 3884 40276 3936
rect 40684 3884 40736 3936
rect 42248 3884 42300 3936
rect 46664 3884 46716 3936
rect 47860 3884 47912 3936
rect 56692 3884 56744 3936
rect 57428 3927 57480 3936
rect 57428 3893 57437 3927
rect 57437 3893 57471 3927
rect 57471 3893 57480 3927
rect 57428 3884 57480 3893
rect 58256 3927 58308 3936
rect 58256 3893 58265 3927
rect 58265 3893 58299 3927
rect 58299 3893 58308 3927
rect 58256 3884 58308 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 9404 3680 9456 3732
rect 12256 3680 12308 3732
rect 20076 3680 20128 3732
rect 20168 3680 20220 3732
rect 22468 3680 22520 3732
rect 7472 3612 7524 3664
rect 7932 3612 7984 3664
rect 8668 3612 8720 3664
rect 10508 3612 10560 3664
rect 12348 3655 12400 3664
rect 12348 3621 12357 3655
rect 12357 3621 12391 3655
rect 12391 3621 12400 3655
rect 12348 3612 12400 3621
rect 12440 3612 12492 3664
rect 14464 3612 14516 3664
rect 15016 3655 15068 3664
rect 15016 3621 15025 3655
rect 15025 3621 15059 3655
rect 15059 3621 15068 3655
rect 15016 3612 15068 3621
rect 17408 3612 17460 3664
rect 18880 3612 18932 3664
rect 19064 3612 19116 3664
rect 9404 3544 9456 3596
rect 9864 3587 9916 3596
rect 9864 3553 9873 3587
rect 9873 3553 9907 3587
rect 9907 3553 9916 3587
rect 9864 3544 9916 3553
rect 9956 3587 10008 3596
rect 9956 3553 9965 3587
rect 9965 3553 9999 3587
rect 9999 3553 10008 3587
rect 10140 3587 10192 3596
rect 9956 3544 10008 3553
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 13268 3587 13320 3596
rect 13268 3553 13277 3587
rect 13277 3553 13311 3587
rect 13311 3553 13320 3587
rect 13268 3544 13320 3553
rect 13728 3587 13780 3596
rect 13728 3553 13737 3587
rect 13737 3553 13771 3587
rect 13771 3553 13780 3587
rect 13728 3544 13780 3553
rect 14924 3544 14976 3596
rect 17132 3544 17184 3596
rect 18972 3544 19024 3596
rect 20444 3612 20496 3664
rect 19432 3587 19484 3596
rect 19432 3553 19441 3587
rect 19441 3553 19475 3587
rect 19475 3553 19484 3587
rect 19432 3544 19484 3553
rect 21732 3587 21784 3596
rect 21732 3553 21741 3587
rect 21741 3553 21775 3587
rect 21775 3553 21784 3587
rect 21732 3544 21784 3553
rect 8300 3476 8352 3528
rect 9312 3476 9364 3528
rect 10692 3476 10744 3528
rect 11980 3476 12032 3528
rect 16212 3476 16264 3528
rect 16580 3519 16632 3528
rect 16580 3485 16589 3519
rect 16589 3485 16623 3519
rect 16623 3485 16632 3519
rect 16580 3476 16632 3485
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 1860 3408 1912 3417
rect 5908 3408 5960 3460
rect 8852 3340 8904 3392
rect 11060 3408 11112 3460
rect 17592 3476 17644 3528
rect 18420 3519 18472 3528
rect 18420 3485 18429 3519
rect 18429 3485 18463 3519
rect 18463 3485 18472 3519
rect 18420 3476 18472 3485
rect 19248 3476 19300 3528
rect 19524 3476 19576 3528
rect 19708 3519 19760 3528
rect 19708 3485 19742 3519
rect 19742 3485 19760 3519
rect 19708 3476 19760 3485
rect 20076 3476 20128 3528
rect 33508 3680 33560 3732
rect 34428 3680 34480 3732
rect 24584 3655 24636 3664
rect 24584 3621 24593 3655
rect 24593 3621 24627 3655
rect 24627 3621 24636 3655
rect 24584 3612 24636 3621
rect 26976 3612 27028 3664
rect 9772 3340 9824 3392
rect 11612 3383 11664 3392
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 11888 3340 11940 3392
rect 14464 3340 14516 3392
rect 17408 3340 17460 3392
rect 18972 3408 19024 3460
rect 19984 3408 20036 3460
rect 24860 3544 24912 3596
rect 25136 3587 25188 3596
rect 25136 3553 25145 3587
rect 25145 3553 25179 3587
rect 25179 3553 25188 3587
rect 25136 3544 25188 3553
rect 26884 3544 26936 3596
rect 29828 3612 29880 3664
rect 29368 3544 29420 3596
rect 30932 3544 30984 3596
rect 33508 3544 33560 3596
rect 23940 3476 23992 3528
rect 27160 3476 27212 3528
rect 28172 3476 28224 3528
rect 28540 3519 28592 3528
rect 28540 3485 28549 3519
rect 28549 3485 28583 3519
rect 28583 3485 28592 3519
rect 28540 3476 28592 3485
rect 29736 3476 29788 3528
rect 30288 3519 30340 3528
rect 30288 3485 30297 3519
rect 30297 3485 30331 3519
rect 30331 3485 30340 3519
rect 30288 3476 30340 3485
rect 19156 3340 19208 3392
rect 20812 3340 20864 3392
rect 24676 3408 24728 3460
rect 28356 3451 28408 3460
rect 27620 3340 27672 3392
rect 28356 3417 28365 3451
rect 28365 3417 28399 3451
rect 28399 3417 28408 3451
rect 28356 3408 28408 3417
rect 28908 3451 28960 3460
rect 28908 3417 28917 3451
rect 28917 3417 28951 3451
rect 28951 3417 28960 3451
rect 28908 3408 28960 3417
rect 30196 3408 30248 3460
rect 31944 3476 31996 3528
rect 32312 3519 32364 3528
rect 32312 3485 32346 3519
rect 32346 3485 32364 3519
rect 32312 3476 32364 3485
rect 32588 3476 32640 3528
rect 34520 3476 34572 3528
rect 34704 3476 34756 3528
rect 37556 3680 37608 3732
rect 44272 3680 44324 3732
rect 44456 3680 44508 3732
rect 46112 3680 46164 3732
rect 39396 3612 39448 3664
rect 39672 3612 39724 3664
rect 40408 3612 40460 3664
rect 35992 3587 36044 3596
rect 35992 3553 36001 3587
rect 36001 3553 36035 3587
rect 36035 3553 36044 3587
rect 35992 3544 36044 3553
rect 37648 3544 37700 3596
rect 38936 3544 38988 3596
rect 35900 3476 35952 3528
rect 36912 3476 36964 3528
rect 38108 3519 38160 3528
rect 31484 3383 31536 3392
rect 31484 3349 31493 3383
rect 31493 3349 31527 3383
rect 31527 3349 31536 3383
rect 31484 3340 31536 3349
rect 32036 3408 32088 3460
rect 33968 3408 34020 3460
rect 34796 3408 34848 3460
rect 38108 3485 38117 3519
rect 38117 3485 38151 3519
rect 38151 3485 38160 3519
rect 38108 3476 38160 3485
rect 39488 3476 39540 3528
rect 40132 3519 40184 3528
rect 40132 3485 40141 3519
rect 40141 3485 40175 3519
rect 40175 3485 40184 3519
rect 40132 3476 40184 3485
rect 32220 3340 32272 3392
rect 33048 3340 33100 3392
rect 33416 3383 33468 3392
rect 33416 3349 33425 3383
rect 33425 3349 33459 3383
rect 33459 3349 33468 3383
rect 33416 3340 33468 3349
rect 33692 3340 33744 3392
rect 34704 3340 34756 3392
rect 37188 3340 37240 3392
rect 38844 3408 38896 3460
rect 41052 3544 41104 3596
rect 41880 3587 41932 3596
rect 41880 3553 41889 3587
rect 41889 3553 41923 3587
rect 41923 3553 41932 3587
rect 41880 3544 41932 3553
rect 41788 3476 41840 3528
rect 42616 3587 42668 3596
rect 42616 3553 42625 3587
rect 42625 3553 42659 3587
rect 42659 3553 42668 3587
rect 42616 3544 42668 3553
rect 42892 3519 42944 3528
rect 42892 3485 42901 3519
rect 42901 3485 42935 3519
rect 42935 3485 42944 3519
rect 42892 3476 42944 3485
rect 43904 3544 43956 3596
rect 43444 3476 43496 3528
rect 43720 3519 43772 3528
rect 43720 3485 43727 3519
rect 43727 3485 43772 3519
rect 43720 3476 43772 3485
rect 44640 3544 44692 3596
rect 45100 3544 45152 3596
rect 45560 3544 45612 3596
rect 45836 3544 45888 3596
rect 44272 3476 44324 3528
rect 45192 3519 45244 3528
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 43352 3408 43404 3460
rect 43904 3451 43956 3460
rect 43904 3417 43913 3451
rect 43913 3417 43947 3451
rect 43947 3417 43956 3451
rect 45744 3519 45796 3528
rect 45744 3485 45753 3519
rect 45753 3485 45787 3519
rect 45787 3485 45796 3519
rect 46020 3519 46072 3528
rect 45744 3476 45796 3485
rect 46020 3485 46029 3519
rect 46029 3485 46063 3519
rect 46063 3485 46072 3519
rect 46020 3476 46072 3485
rect 46204 3476 46256 3528
rect 47584 3680 47636 3732
rect 48044 3723 48096 3732
rect 48044 3689 48053 3723
rect 48053 3689 48087 3723
rect 48087 3689 48096 3723
rect 48044 3680 48096 3689
rect 49884 3680 49936 3732
rect 51264 3723 51316 3732
rect 51264 3689 51273 3723
rect 51273 3689 51307 3723
rect 51307 3689 51316 3723
rect 51264 3680 51316 3689
rect 52736 3723 52788 3732
rect 52736 3689 52745 3723
rect 52745 3689 52779 3723
rect 52779 3689 52788 3723
rect 52736 3680 52788 3689
rect 52920 3680 52972 3732
rect 53564 3680 53616 3732
rect 58256 3680 58308 3732
rect 47124 3612 47176 3664
rect 50896 3612 50948 3664
rect 53196 3612 53248 3664
rect 46940 3544 46992 3596
rect 46848 3476 46900 3528
rect 43904 3408 43956 3417
rect 47124 3408 47176 3460
rect 39120 3340 39172 3392
rect 44548 3340 44600 3392
rect 47400 3408 47452 3460
rect 50804 3544 50856 3596
rect 50620 3476 50672 3528
rect 51724 3476 51776 3528
rect 49240 3408 49292 3460
rect 49516 3408 49568 3460
rect 50896 3408 50948 3460
rect 52276 3408 52328 3460
rect 56692 3544 56744 3596
rect 57428 3476 57480 3528
rect 53196 3408 53248 3460
rect 47308 3383 47360 3392
rect 47308 3349 47317 3383
rect 47317 3349 47351 3383
rect 47351 3349 47360 3383
rect 47308 3340 47360 3349
rect 47584 3340 47636 3392
rect 54668 3340 54720 3392
rect 57244 3340 57296 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 6000 3136 6052 3188
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 8392 3179 8444 3188
rect 8392 3145 8401 3179
rect 8401 3145 8435 3179
rect 8435 3145 8444 3179
rect 8392 3136 8444 3145
rect 9128 3179 9180 3188
rect 9128 3145 9137 3179
rect 9137 3145 9171 3179
rect 9171 3145 9180 3179
rect 9128 3136 9180 3145
rect 9680 3136 9732 3188
rect 11980 3136 12032 3188
rect 15016 3136 15068 3188
rect 8116 3068 8168 3120
rect 10692 3111 10744 3120
rect 8852 3000 8904 3052
rect 9036 3043 9088 3052
rect 9036 3009 9045 3043
rect 9045 3009 9079 3043
rect 9079 3009 9088 3043
rect 9036 3000 9088 3009
rect 9220 2932 9272 2984
rect 9680 3000 9732 3052
rect 10692 3077 10701 3111
rect 10701 3077 10735 3111
rect 10735 3077 10744 3111
rect 10692 3068 10744 3077
rect 11888 3111 11940 3120
rect 11888 3077 11897 3111
rect 11897 3077 11931 3111
rect 11931 3077 11940 3111
rect 11888 3068 11940 3077
rect 10140 3043 10192 3052
rect 10140 3009 10149 3043
rect 10149 3009 10183 3043
rect 10183 3009 10192 3043
rect 10140 3000 10192 3009
rect 9404 2932 9456 2984
rect 9864 2975 9916 2984
rect 9864 2941 9873 2975
rect 9873 2941 9907 2975
rect 9907 2941 9916 2975
rect 9864 2932 9916 2941
rect 12256 2932 12308 2984
rect 13820 3000 13872 3052
rect 14280 3000 14332 3052
rect 14832 3000 14884 3052
rect 17500 3068 17552 3120
rect 19340 3111 19392 3120
rect 19340 3077 19374 3111
rect 19374 3077 19392 3111
rect 19340 3068 19392 3077
rect 15568 3000 15620 3052
rect 16488 3000 16540 3052
rect 17224 3043 17276 3052
rect 17224 3009 17233 3043
rect 17233 3009 17267 3043
rect 17267 3009 17276 3043
rect 17224 3000 17276 3009
rect 8852 2796 8904 2848
rect 9864 2796 9916 2848
rect 10876 2864 10928 2916
rect 13544 2907 13596 2916
rect 13544 2873 13553 2907
rect 13553 2873 13587 2907
rect 13587 2873 13596 2907
rect 13544 2864 13596 2873
rect 12624 2796 12676 2848
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 19064 3043 19116 3052
rect 18144 3000 18196 3009
rect 19064 3009 19073 3043
rect 19073 3009 19107 3043
rect 19107 3009 19116 3043
rect 19064 3000 19116 3009
rect 20168 3000 20220 3052
rect 21180 3000 21232 3052
rect 22284 3136 22336 3188
rect 33416 3136 33468 3188
rect 33784 3136 33836 3188
rect 22192 3000 22244 3052
rect 23204 3068 23256 3120
rect 23940 3068 23992 3120
rect 16396 2864 16448 2916
rect 15016 2796 15068 2848
rect 21088 2932 21140 2984
rect 23572 3000 23624 3052
rect 24584 3000 24636 3052
rect 20260 2864 20312 2916
rect 20720 2796 20772 2848
rect 22744 2796 22796 2848
rect 26056 2932 26108 2984
rect 26424 2932 26476 2984
rect 24860 2907 24912 2916
rect 24860 2873 24869 2907
rect 24869 2873 24903 2907
rect 24903 2873 24912 2907
rect 24860 2864 24912 2873
rect 24952 2864 25004 2916
rect 27712 2864 27764 2916
rect 28080 3000 28132 3052
rect 29276 3068 29328 3120
rect 30748 3068 30800 3120
rect 32404 3068 32456 3120
rect 37924 3136 37976 3188
rect 39948 3136 40000 3188
rect 42800 3179 42852 3188
rect 42800 3145 42809 3179
rect 42809 3145 42843 3179
rect 42843 3145 42852 3179
rect 42800 3136 42852 3145
rect 43904 3136 43956 3188
rect 47952 3179 48004 3188
rect 47952 3145 47961 3179
rect 47961 3145 47995 3179
rect 47995 3145 48004 3179
rect 47952 3136 48004 3145
rect 48688 3179 48740 3188
rect 48688 3145 48697 3179
rect 48697 3145 48731 3179
rect 48731 3145 48740 3179
rect 48688 3136 48740 3145
rect 49792 3179 49844 3188
rect 49792 3145 49801 3179
rect 49801 3145 49835 3179
rect 49835 3145 49844 3179
rect 49792 3136 49844 3145
rect 50988 3136 51040 3188
rect 52184 3136 52236 3188
rect 52460 3136 52512 3188
rect 53932 3136 53984 3188
rect 58256 3179 58308 3188
rect 39396 3068 39448 3120
rect 39672 3068 39724 3120
rect 40868 3068 40920 3120
rect 41604 3111 41656 3120
rect 41604 3077 41613 3111
rect 41613 3077 41647 3111
rect 41647 3077 41656 3111
rect 41604 3068 41656 3077
rect 45008 3068 45060 3120
rect 31208 3000 31260 3052
rect 31484 3000 31536 3052
rect 33232 3043 33284 3052
rect 33232 3009 33241 3043
rect 33241 3009 33275 3043
rect 33275 3009 33284 3043
rect 33232 3000 33284 3009
rect 30748 2932 30800 2984
rect 31576 2932 31628 2984
rect 32956 2932 33008 2984
rect 33968 3000 34020 3052
rect 34520 3000 34572 3052
rect 35808 3000 35860 3052
rect 37464 3043 37516 3052
rect 37464 3009 37473 3043
rect 37473 3009 37507 3043
rect 37507 3009 37516 3043
rect 37464 3000 37516 3009
rect 24400 2796 24452 2848
rect 27988 2796 28040 2848
rect 29736 2864 29788 2916
rect 32128 2864 32180 2916
rect 35624 2932 35676 2984
rect 38660 3000 38712 3052
rect 39304 3043 39356 3052
rect 39304 3009 39313 3043
rect 39313 3009 39347 3043
rect 39347 3009 39356 3043
rect 39304 3000 39356 3009
rect 39580 3000 39632 3052
rect 40408 3000 40460 3052
rect 41328 3000 41380 3052
rect 44272 3000 44324 3052
rect 44916 3043 44968 3052
rect 35348 2864 35400 2916
rect 31760 2796 31812 2848
rect 31852 2796 31904 2848
rect 33416 2796 33468 2848
rect 33600 2796 33652 2848
rect 35992 2796 36044 2848
rect 36544 2796 36596 2848
rect 42340 2932 42392 2984
rect 44456 2932 44508 2984
rect 44916 3009 44925 3043
rect 44925 3009 44959 3043
rect 44959 3009 44968 3043
rect 44916 3000 44968 3009
rect 45100 3000 45152 3052
rect 45744 3000 45796 3052
rect 46112 3043 46164 3052
rect 46112 3009 46121 3043
rect 46121 3009 46155 3043
rect 46155 3009 46164 3043
rect 46112 3000 46164 3009
rect 51540 3068 51592 3120
rect 53380 3068 53432 3120
rect 56600 3111 56652 3120
rect 56600 3077 56609 3111
rect 56609 3077 56643 3111
rect 56643 3077 56652 3111
rect 56600 3068 56652 3077
rect 44824 2864 44876 2916
rect 45652 2932 45704 2984
rect 48412 3000 48464 3052
rect 48688 3000 48740 3052
rect 48136 2932 48188 2984
rect 49792 2932 49844 2984
rect 47308 2864 47360 2916
rect 50068 2864 50120 2916
rect 52000 3000 52052 3052
rect 54668 3043 54720 3052
rect 52552 2932 52604 2984
rect 54668 3009 54677 3043
rect 54677 3009 54711 3043
rect 54711 3009 54720 3043
rect 54668 3000 54720 3009
rect 56508 3000 56560 3052
rect 58256 3145 58265 3179
rect 58265 3145 58299 3179
rect 58299 3145 58308 3179
rect 58256 3136 58308 3145
rect 58164 3111 58216 3120
rect 58164 3077 58173 3111
rect 58173 3077 58207 3111
rect 58207 3077 58216 3111
rect 58164 3068 58216 3077
rect 57980 3000 58032 3052
rect 55312 2932 55364 2984
rect 40684 2796 40736 2848
rect 41420 2796 41472 2848
rect 43444 2796 43496 2848
rect 44916 2796 44968 2848
rect 45284 2796 45336 2848
rect 46388 2796 46440 2848
rect 51356 2796 51408 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 10784 2592 10836 2644
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 1860 2388 1912 2397
rect 6828 2388 6880 2440
rect 8484 2524 8536 2576
rect 8668 2524 8720 2576
rect 10416 2567 10468 2576
rect 10416 2533 10425 2567
rect 10425 2533 10459 2567
rect 10459 2533 10468 2567
rect 10416 2524 10468 2533
rect 10508 2524 10560 2576
rect 9588 2456 9640 2508
rect 10692 2456 10744 2508
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 7012 2295 7064 2304
rect 7012 2261 7021 2295
rect 7021 2261 7055 2295
rect 7055 2261 7064 2295
rect 7012 2252 7064 2261
rect 7748 2295 7800 2304
rect 7748 2261 7757 2295
rect 7757 2261 7791 2295
rect 7791 2261 7800 2295
rect 7748 2252 7800 2261
rect 9404 2320 9456 2372
rect 8944 2252 8996 2304
rect 9680 2363 9732 2372
rect 9680 2329 9689 2363
rect 9689 2329 9723 2363
rect 9723 2329 9732 2363
rect 9680 2320 9732 2329
rect 14740 2592 14792 2644
rect 18880 2592 18932 2644
rect 13176 2524 13228 2576
rect 14372 2524 14424 2576
rect 24952 2592 25004 2644
rect 16028 2456 16080 2508
rect 12440 2320 12492 2372
rect 14372 2320 14424 2372
rect 14004 2252 14056 2304
rect 15752 2388 15804 2440
rect 16304 2388 16356 2440
rect 22376 2456 22428 2508
rect 19156 2388 19208 2440
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 20996 2431 21048 2440
rect 20996 2397 21005 2431
rect 21005 2397 21039 2431
rect 21039 2397 21048 2431
rect 20996 2388 21048 2397
rect 15200 2363 15252 2372
rect 15200 2329 15209 2363
rect 15209 2329 15243 2363
rect 15243 2329 15252 2363
rect 15200 2320 15252 2329
rect 16120 2363 16172 2372
rect 16120 2329 16129 2363
rect 16129 2329 16163 2363
rect 16163 2329 16172 2363
rect 16120 2320 16172 2329
rect 18512 2320 18564 2372
rect 20260 2320 20312 2372
rect 24216 2524 24268 2576
rect 24952 2456 25004 2508
rect 23388 2388 23440 2440
rect 27068 2592 27120 2644
rect 41144 2635 41196 2644
rect 41144 2601 41153 2635
rect 41153 2601 41187 2635
rect 41187 2601 41196 2635
rect 41144 2592 41196 2601
rect 44640 2592 44692 2644
rect 45100 2592 45152 2644
rect 45284 2592 45336 2644
rect 45376 2592 45428 2644
rect 46480 2635 46532 2644
rect 46480 2601 46489 2635
rect 46489 2601 46523 2635
rect 46523 2601 46532 2635
rect 46480 2592 46532 2601
rect 49056 2592 49108 2644
rect 51448 2635 51500 2644
rect 51448 2601 51457 2635
rect 51457 2601 51491 2635
rect 51491 2601 51500 2635
rect 51448 2592 51500 2601
rect 53104 2635 53156 2644
rect 53104 2601 53113 2635
rect 53113 2601 53147 2635
rect 53147 2601 53156 2635
rect 53104 2592 53156 2601
rect 57980 2592 58032 2644
rect 27896 2524 27948 2576
rect 36820 2524 36872 2576
rect 28080 2456 28132 2508
rect 29184 2456 29236 2508
rect 26240 2388 26292 2440
rect 28172 2388 28224 2440
rect 30104 2388 30156 2440
rect 31208 2456 31260 2508
rect 33416 2499 33468 2508
rect 33416 2465 33425 2499
rect 33425 2465 33459 2499
rect 33459 2465 33468 2499
rect 33416 2456 33468 2465
rect 35992 2499 36044 2508
rect 35992 2465 36001 2499
rect 36001 2465 36035 2499
rect 36035 2465 36044 2499
rect 35992 2456 36044 2465
rect 46204 2524 46256 2576
rect 33048 2388 33100 2440
rect 34796 2388 34848 2440
rect 35716 2388 35768 2440
rect 51356 2524 51408 2576
rect 48964 2499 49016 2508
rect 18604 2252 18656 2304
rect 23480 2320 23532 2372
rect 25780 2320 25832 2372
rect 26608 2320 26660 2372
rect 26884 2320 26936 2372
rect 29920 2320 29972 2372
rect 30472 2363 30524 2372
rect 30472 2329 30481 2363
rect 30481 2329 30515 2363
rect 30515 2329 30524 2363
rect 30472 2320 30524 2329
rect 31024 2320 31076 2372
rect 24124 2252 24176 2304
rect 25228 2252 25280 2304
rect 29644 2252 29696 2304
rect 31300 2252 31352 2304
rect 32680 2320 32732 2372
rect 35440 2320 35492 2372
rect 37280 2320 37332 2372
rect 39396 2388 39448 2440
rect 39488 2388 39540 2440
rect 40132 2388 40184 2440
rect 41144 2388 41196 2440
rect 43536 2431 43588 2440
rect 43536 2397 43545 2431
rect 43545 2397 43579 2431
rect 43579 2397 43588 2431
rect 43536 2388 43588 2397
rect 48964 2465 48973 2499
rect 48973 2465 49007 2499
rect 49007 2465 49016 2499
rect 48964 2456 49016 2465
rect 54760 2499 54812 2508
rect 54760 2465 54769 2499
rect 54769 2465 54803 2499
rect 54803 2465 54812 2499
rect 54760 2456 54812 2465
rect 44272 2388 44324 2440
rect 45192 2431 45244 2440
rect 45192 2397 45201 2431
rect 45201 2397 45235 2431
rect 45235 2397 45244 2431
rect 45192 2388 45244 2397
rect 45284 2388 45336 2440
rect 45560 2431 45612 2440
rect 45560 2397 45574 2431
rect 45574 2397 45608 2431
rect 45608 2397 45612 2431
rect 45560 2388 45612 2397
rect 34336 2252 34388 2304
rect 40500 2320 40552 2372
rect 43352 2320 43404 2372
rect 44732 2320 44784 2372
rect 46664 2388 46716 2440
rect 48044 2388 48096 2440
rect 51172 2388 51224 2440
rect 53656 2388 53708 2440
rect 57244 2388 57296 2440
rect 58164 2431 58216 2440
rect 58164 2397 58173 2431
rect 58173 2397 58207 2431
rect 58207 2397 58216 2431
rect 58164 2388 58216 2397
rect 42616 2252 42668 2304
rect 47584 2320 47636 2372
rect 48964 2320 49016 2372
rect 51356 2363 51408 2372
rect 51356 2329 51365 2363
rect 51365 2329 51399 2363
rect 51399 2329 51408 2363
rect 51356 2320 51408 2329
rect 53932 2320 53984 2372
rect 47952 2295 48004 2304
rect 47952 2261 47961 2295
rect 47961 2261 47995 2295
rect 47995 2261 48004 2295
rect 47952 2252 48004 2261
rect 52828 2252 52880 2304
rect 57336 2363 57388 2372
rect 57336 2329 57345 2363
rect 57345 2329 57379 2363
rect 57379 2329 57388 2363
rect 57336 2320 57388 2329
rect 55680 2295 55732 2304
rect 55680 2261 55689 2295
rect 55689 2261 55723 2295
rect 55723 2261 55732 2295
rect 55680 2252 55732 2261
rect 56416 2295 56468 2304
rect 56416 2261 56425 2295
rect 56425 2261 56459 2295
rect 56459 2261 56468 2295
rect 56416 2252 56468 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 9404 2048 9456 2100
rect 12716 2048 12768 2100
rect 15200 2048 15252 2100
rect 19708 2048 19760 2100
rect 20996 2048 21048 2100
rect 24032 2048 24084 2100
rect 45192 2048 45244 2100
rect 55680 2048 55732 2100
rect 1584 1980 1636 2032
rect 7012 1912 7064 1964
rect 11520 1912 11572 1964
rect 12808 1912 12860 1964
rect 5172 1844 5224 1896
rect 17684 1844 17736 1896
rect 18512 1912 18564 1964
rect 21916 1912 21968 1964
rect 22376 1980 22428 2032
rect 31668 1980 31720 2032
rect 38108 1980 38160 2032
rect 56416 1980 56468 2032
rect 28356 1912 28408 1964
rect 31208 1844 31260 1896
rect 9680 1776 9732 1828
rect 14556 1776 14608 1828
rect 20628 1776 20680 1828
rect 40500 1912 40552 1964
rect 7748 1708 7800 1760
rect 12624 1708 12676 1760
rect 16120 1708 16172 1760
rect 20536 1708 20588 1760
rect 19248 1640 19300 1692
rect 26240 1640 26292 1692
rect 9312 1504 9364 1556
rect 10876 1504 10928 1556
rect 9864 1436 9916 1488
rect 12256 1436 12308 1488
rect 33232 1436 33284 1488
rect 33600 1436 33652 1488
rect 6828 1368 6880 1420
rect 7564 1368 7616 1420
rect 8484 1368 8536 1420
rect 11152 1368 11204 1420
rect 12440 1368 12492 1420
rect 13912 1368 13964 1420
rect 14372 1368 14424 1420
rect 15292 1368 15344 1420
rect 34060 1368 34112 1420
rect 35900 1368 35952 1420
rect 50344 1368 50396 1420
rect 51356 1368 51408 1420
rect 50712 1300 50764 1352
rect 56508 1300 56560 1352
<< metal2 >>
rect 846 63200 902 64000
rect 1582 63200 1638 64000
rect 2318 63322 2374 64000
rect 3054 63322 3110 64000
rect 3790 63322 3846 64000
rect 4526 63322 4582 64000
rect 5262 63322 5318 64000
rect 5998 63322 6054 64000
rect 2318 63294 2544 63322
rect 2318 63200 2374 63294
rect 860 59702 888 63200
rect 1596 60110 1624 63200
rect 1676 61124 1728 61130
rect 1676 61066 1728 61072
rect 1688 60897 1716 61066
rect 1674 60888 1730 60897
rect 1674 60823 1730 60832
rect 1676 60784 1728 60790
rect 1676 60726 1728 60732
rect 1688 60217 1716 60726
rect 1952 60512 2004 60518
rect 1952 60454 2004 60460
rect 1674 60208 1730 60217
rect 1674 60143 1730 60152
rect 1584 60104 1636 60110
rect 1584 60046 1636 60052
rect 848 59696 900 59702
rect 848 59638 900 59644
rect 1584 59628 1636 59634
rect 1584 59570 1636 59576
rect 1596 59537 1624 59570
rect 1582 59528 1638 59537
rect 1582 59463 1638 59472
rect 1964 59090 1992 60454
rect 2516 60110 2544 63294
rect 3054 63294 3280 63322
rect 3054 63200 3110 63294
rect 2778 61568 2834 61577
rect 2778 61503 2834 61512
rect 2792 61266 2820 61503
rect 2780 61260 2832 61266
rect 2780 61202 2832 61208
rect 3252 60790 3280 63294
rect 3790 63294 4016 63322
rect 3790 63200 3846 63294
rect 3988 60790 4016 63294
rect 4526 63294 4660 63322
rect 4526 63200 4582 63294
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 4632 61198 4660 63294
rect 5092 63294 5318 63322
rect 5092 61198 5120 63294
rect 5262 63200 5318 63294
rect 5828 63294 6054 63322
rect 5828 61198 5856 63294
rect 5998 63200 6054 63294
rect 6734 63200 6790 64000
rect 7470 63322 7526 64000
rect 7470 63294 7604 63322
rect 7470 63200 7526 63294
rect 6184 61328 6236 61334
rect 6184 61270 6236 61276
rect 4620 61192 4672 61198
rect 4620 61134 4672 61140
rect 5080 61192 5132 61198
rect 5080 61134 5132 61140
rect 5816 61192 5868 61198
rect 5816 61134 5868 61140
rect 4896 61124 4948 61130
rect 4896 61066 4948 61072
rect 3240 60784 3292 60790
rect 3240 60726 3292 60732
rect 3976 60784 4028 60790
rect 3976 60726 4028 60732
rect 4804 60580 4856 60586
rect 4804 60522 4856 60528
rect 3332 60512 3384 60518
rect 3332 60454 3384 60460
rect 2504 60104 2556 60110
rect 2504 60046 2556 60052
rect 2044 60036 2096 60042
rect 2044 59978 2096 59984
rect 1952 59084 2004 59090
rect 1952 59026 2004 59032
rect 1584 59016 1636 59022
rect 1584 58958 1636 58964
rect 1596 58857 1624 58958
rect 1768 58880 1820 58886
rect 1582 58848 1638 58857
rect 1768 58822 1820 58828
rect 1582 58783 1638 58792
rect 1676 58540 1728 58546
rect 1676 58482 1728 58488
rect 1688 58177 1716 58482
rect 1674 58168 1730 58177
rect 1674 58103 1730 58112
rect 1584 57928 1636 57934
rect 1584 57870 1636 57876
rect 1596 57497 1624 57870
rect 1582 57488 1638 57497
rect 1582 57423 1638 57432
rect 1780 57050 1808 58822
rect 1952 57792 2004 57798
rect 1952 57734 2004 57740
rect 1768 57044 1820 57050
rect 1768 56986 1820 56992
rect 1676 56840 1728 56846
rect 1674 56808 1676 56817
rect 1728 56808 1730 56817
rect 1674 56743 1730 56752
rect 1676 56364 1728 56370
rect 1676 56306 1728 56312
rect 1688 56137 1716 56306
rect 1768 56160 1820 56166
rect 1674 56128 1730 56137
rect 1768 56102 1820 56108
rect 1674 56063 1730 56072
rect 1780 55962 1808 56102
rect 1768 55956 1820 55962
rect 1768 55898 1820 55904
rect 1676 55684 1728 55690
rect 1676 55626 1728 55632
rect 1688 55457 1716 55626
rect 1674 55448 1730 55457
rect 1674 55383 1730 55392
rect 1584 55276 1636 55282
rect 1584 55218 1636 55224
rect 1596 54777 1624 55218
rect 1582 54768 1638 54777
rect 1582 54703 1638 54712
rect 1676 54188 1728 54194
rect 1676 54130 1728 54136
rect 1688 54097 1716 54130
rect 1674 54088 1730 54097
rect 1674 54023 1730 54032
rect 1584 53576 1636 53582
rect 1584 53518 1636 53524
rect 1596 53417 1624 53518
rect 1582 53408 1638 53417
rect 1582 53343 1638 53352
rect 1964 53174 1992 57734
rect 1952 53168 2004 53174
rect 1952 53110 2004 53116
rect 1584 53100 1636 53106
rect 1584 53042 1636 53048
rect 1596 52737 1624 53042
rect 1860 52896 1912 52902
rect 1860 52838 1912 52844
rect 1582 52728 1638 52737
rect 1582 52663 1638 52672
rect 1676 52420 1728 52426
rect 1676 52362 1728 52368
rect 1688 52057 1716 52362
rect 1674 52048 1730 52057
rect 1674 51983 1730 51992
rect 1674 51368 1730 51377
rect 1674 51303 1676 51312
rect 1728 51303 1730 51312
rect 1676 51274 1728 51280
rect 1676 50924 1728 50930
rect 1676 50866 1728 50872
rect 1688 50697 1716 50866
rect 1674 50688 1730 50697
rect 1674 50623 1730 50632
rect 1676 50244 1728 50250
rect 1676 50186 1728 50192
rect 1688 50017 1716 50186
rect 1674 50008 1730 50017
rect 1674 49943 1730 49952
rect 1676 49836 1728 49842
rect 1676 49778 1728 49784
rect 1688 49337 1716 49778
rect 1674 49328 1730 49337
rect 1674 49263 1730 49272
rect 1676 48748 1728 48754
rect 1676 48690 1728 48696
rect 1688 48657 1716 48690
rect 1674 48648 1730 48657
rect 1674 48583 1730 48592
rect 1676 48068 1728 48074
rect 1676 48010 1728 48016
rect 1688 47977 1716 48010
rect 1674 47968 1730 47977
rect 1674 47903 1730 47912
rect 1676 47660 1728 47666
rect 1676 47602 1728 47608
rect 1492 47456 1544 47462
rect 1492 47398 1544 47404
rect 1400 41132 1452 41138
rect 1400 41074 1452 41080
rect 1412 40497 1440 41074
rect 1398 40488 1454 40497
rect 1398 40423 1454 40432
rect 1400 39364 1452 39370
rect 1400 39306 1452 39312
rect 1412 38457 1440 39306
rect 1398 38448 1454 38457
rect 1398 38383 1454 38392
rect 1400 36780 1452 36786
rect 1400 36722 1452 36728
rect 1412 35737 1440 36722
rect 1398 35728 1454 35737
rect 1398 35663 1454 35672
rect 1504 35086 1532 47398
rect 1688 47297 1716 47602
rect 1674 47288 1730 47297
rect 1674 47223 1730 47232
rect 1676 46980 1728 46986
rect 1676 46922 1728 46928
rect 1688 46617 1716 46922
rect 1674 46608 1730 46617
rect 1674 46543 1730 46552
rect 1674 45928 1730 45937
rect 1674 45863 1676 45872
rect 1728 45863 1730 45872
rect 1676 45834 1728 45840
rect 1584 45484 1636 45490
rect 1584 45426 1636 45432
rect 1596 45257 1624 45426
rect 1582 45248 1638 45257
rect 1582 45183 1638 45192
rect 1676 44804 1728 44810
rect 1676 44746 1728 44752
rect 1688 44577 1716 44746
rect 1674 44568 1730 44577
rect 1674 44503 1730 44512
rect 1676 44396 1728 44402
rect 1676 44338 1728 44344
rect 1688 43897 1716 44338
rect 1674 43888 1730 43897
rect 1674 43823 1730 43832
rect 1584 43308 1636 43314
rect 1584 43250 1636 43256
rect 1596 43217 1624 43250
rect 1582 43208 1638 43217
rect 1582 43143 1638 43152
rect 1676 42628 1728 42634
rect 1676 42570 1728 42576
rect 1688 42537 1716 42570
rect 1674 42528 1730 42537
rect 1674 42463 1730 42472
rect 1676 42220 1728 42226
rect 1676 42162 1728 42168
rect 1688 41857 1716 42162
rect 1674 41848 1730 41857
rect 1674 41783 1730 41792
rect 1676 41540 1728 41546
rect 1676 41482 1728 41488
rect 1688 41177 1716 41482
rect 1674 41168 1730 41177
rect 1674 41103 1730 41112
rect 1676 40452 1728 40458
rect 1676 40394 1728 40400
rect 1584 40112 1636 40118
rect 1584 40054 1636 40060
rect 1596 39137 1624 40054
rect 1688 39817 1716 40394
rect 1674 39808 1730 39817
rect 1674 39743 1730 39752
rect 1582 39128 1638 39137
rect 1582 39063 1638 39072
rect 1676 38956 1728 38962
rect 1676 38898 1728 38904
rect 1688 37777 1716 38898
rect 1674 37768 1730 37777
rect 1674 37703 1730 37712
rect 1584 37256 1636 37262
rect 1584 37198 1636 37204
rect 1596 36417 1624 37198
rect 1768 36848 1820 36854
rect 1768 36790 1820 36796
rect 1582 36408 1638 36417
rect 1780 36378 1808 36790
rect 1582 36343 1638 36352
rect 1768 36372 1820 36378
rect 1768 36314 1820 36320
rect 1872 36310 1900 52838
rect 1952 37936 2004 37942
rect 1952 37878 2004 37884
rect 1860 36304 1912 36310
rect 1860 36246 1912 36252
rect 1676 36100 1728 36106
rect 1676 36042 1728 36048
rect 1492 35080 1544 35086
rect 1688 35057 1716 36042
rect 1860 35760 1912 35766
rect 1860 35702 1912 35708
rect 1492 35022 1544 35028
rect 1674 35048 1730 35057
rect 1674 34983 1730 34992
rect 1676 34604 1728 34610
rect 1676 34546 1728 34552
rect 1688 34377 1716 34546
rect 1674 34368 1730 34377
rect 1674 34303 1730 34312
rect 1872 34134 1900 35702
rect 1860 34128 1912 34134
rect 1860 34070 1912 34076
rect 1676 33924 1728 33930
rect 1676 33866 1728 33872
rect 1688 33697 1716 33866
rect 1674 33688 1730 33697
rect 1674 33623 1730 33632
rect 1964 33590 1992 37878
rect 2056 35698 2084 59978
rect 2412 59968 2464 59974
rect 2412 59910 2464 59916
rect 2424 40118 2452 59910
rect 2596 59492 2648 59498
rect 2596 59434 2648 59440
rect 2412 40112 2464 40118
rect 2412 40054 2464 40060
rect 2504 39364 2556 39370
rect 2504 39306 2556 39312
rect 2516 38350 2544 39306
rect 2608 38418 2636 59434
rect 2688 59424 2740 59430
rect 2688 59366 2740 59372
rect 2700 56914 2728 59366
rect 2688 56908 2740 56914
rect 2688 56850 2740 56856
rect 3344 48822 3372 60454
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4620 51944 4672 51950
rect 4620 51886 4672 51892
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 3332 48816 3384 48822
rect 3332 48758 3384 48764
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4068 43104 4120 43110
rect 4068 43046 4120 43052
rect 3792 42356 3844 42362
rect 3792 42298 3844 42304
rect 3804 41274 3832 42298
rect 4080 42090 4108 43046
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4632 42226 4660 51886
rect 4620 42220 4672 42226
rect 4620 42162 4672 42168
rect 4068 42084 4120 42090
rect 4068 42026 4120 42032
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 3976 41540 4028 41546
rect 3976 41482 4028 41488
rect 3884 41472 3936 41478
rect 3884 41414 3936 41420
rect 2964 41268 3016 41274
rect 2964 41210 3016 41216
rect 3792 41268 3844 41274
rect 3792 41210 3844 41216
rect 2780 40384 2832 40390
rect 2780 40326 2832 40332
rect 2792 40118 2820 40326
rect 2780 40112 2832 40118
rect 2780 40054 2832 40060
rect 2976 40050 3004 41210
rect 3896 41138 3924 41414
rect 3988 41206 4016 41482
rect 4632 41478 4660 42162
rect 4620 41472 4672 41478
rect 4620 41414 4672 41420
rect 3976 41200 4028 41206
rect 3976 41142 4028 41148
rect 3884 41132 3936 41138
rect 3884 41074 3936 41080
rect 3896 40186 3924 41074
rect 4816 41070 4844 60522
rect 4908 42158 4936 61066
rect 5172 61056 5224 61062
rect 5172 60998 5224 61004
rect 5908 61056 5960 61062
rect 5908 60998 5960 61004
rect 5184 52018 5212 60998
rect 5920 60858 5948 60998
rect 5908 60852 5960 60858
rect 5908 60794 5960 60800
rect 5448 52488 5500 52494
rect 5448 52430 5500 52436
rect 5460 52086 5488 52430
rect 5448 52080 5500 52086
rect 5448 52022 5500 52028
rect 5172 52012 5224 52018
rect 5172 51954 5224 51960
rect 5724 51808 5776 51814
rect 5724 51750 5776 51756
rect 5540 42628 5592 42634
rect 5540 42570 5592 42576
rect 4896 42152 4948 42158
rect 4896 42094 4948 42100
rect 4988 42016 5040 42022
rect 4988 41958 5040 41964
rect 5000 41750 5028 41958
rect 4988 41744 5040 41750
rect 4988 41686 5040 41692
rect 5552 41070 5580 42570
rect 4804 41064 4856 41070
rect 4804 41006 4856 41012
rect 5540 41064 5592 41070
rect 5540 41006 5592 41012
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 3884 40180 3936 40186
rect 3884 40122 3936 40128
rect 2688 40044 2740 40050
rect 2688 39986 2740 39992
rect 2964 40044 3016 40050
rect 2964 39986 3016 39992
rect 2700 38434 2728 39986
rect 2976 38486 3004 39986
rect 3056 39840 3108 39846
rect 3056 39782 3108 39788
rect 3068 39642 3096 39782
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 3056 39636 3108 39642
rect 3056 39578 3108 39584
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 2964 38480 3016 38486
rect 2596 38412 2648 38418
rect 2700 38406 2912 38434
rect 2964 38422 3016 38428
rect 3700 38480 3752 38486
rect 3700 38422 3752 38428
rect 2596 38354 2648 38360
rect 2504 38344 2556 38350
rect 2504 38286 2556 38292
rect 2688 38344 2740 38350
rect 2688 38286 2740 38292
rect 2700 38010 2728 38286
rect 2688 38004 2740 38010
rect 2688 37946 2740 37952
rect 2792 37890 2820 38406
rect 2884 38350 2912 38406
rect 2872 38344 2924 38350
rect 2872 38286 2924 38292
rect 2320 37868 2372 37874
rect 2320 37810 2372 37816
rect 2504 37868 2556 37874
rect 2504 37810 2556 37816
rect 2700 37862 2820 37890
rect 3712 37874 3740 38422
rect 3700 37868 3752 37874
rect 2136 37120 2188 37126
rect 2136 37062 2188 37068
rect 2044 35692 2096 35698
rect 2044 35634 2096 35640
rect 1952 33584 2004 33590
rect 1952 33526 2004 33532
rect 1676 33516 1728 33522
rect 1676 33458 1728 33464
rect 1688 33017 1716 33458
rect 1674 33008 1730 33017
rect 1674 32943 1730 32952
rect 1676 32428 1728 32434
rect 1676 32370 1728 32376
rect 1688 32337 1716 32370
rect 1674 32328 1730 32337
rect 1674 32263 1730 32272
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 1688 31657 1716 31758
rect 1674 31648 1730 31657
rect 1674 31583 1730 31592
rect 1676 31340 1728 31346
rect 1676 31282 1728 31288
rect 1688 30977 1716 31282
rect 1674 30968 1730 30977
rect 1674 30903 1730 30912
rect 1676 30660 1728 30666
rect 1676 30602 1728 30608
rect 1688 30297 1716 30602
rect 1674 30288 1730 30297
rect 1674 30223 1730 30232
rect 1858 29608 1914 29617
rect 1858 29543 1860 29552
rect 1912 29543 1914 29552
rect 1860 29514 1912 29520
rect 1768 29096 1820 29102
rect 1768 29038 1820 29044
rect 1780 28937 1808 29038
rect 1766 28928 1822 28937
rect 1766 28863 1822 28872
rect 1584 28552 1636 28558
rect 1584 28494 1636 28500
rect 1596 28218 1624 28494
rect 1860 28484 1912 28490
rect 1860 28426 1912 28432
rect 1872 28257 1900 28426
rect 1858 28248 1914 28257
rect 1584 28212 1636 28218
rect 1858 28183 1914 28192
rect 1584 28154 1636 28160
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 27674 1440 28018
rect 1584 28008 1636 28014
rect 1584 27950 1636 27956
rect 1400 27668 1452 27674
rect 1400 27610 1452 27616
rect 1596 27577 1624 27950
rect 1582 27568 1638 27577
rect 1582 27503 1638 27512
rect 1768 26920 1820 26926
rect 1766 26888 1768 26897
rect 1820 26888 1822 26897
rect 1766 26823 1822 26832
rect 1860 26308 1912 26314
rect 1860 26250 1912 26256
rect 1872 26217 1900 26250
rect 1858 26208 1914 26217
rect 1858 26143 1914 26152
rect 1768 25832 1820 25838
rect 1768 25774 1820 25780
rect 1780 25537 1808 25774
rect 1766 25528 1822 25537
rect 1766 25463 1822 25472
rect 1584 25288 1636 25294
rect 1584 25230 1636 25236
rect 1596 24954 1624 25230
rect 1860 25220 1912 25226
rect 1860 25162 1912 25168
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1872 24857 1900 25162
rect 1858 24848 1914 24857
rect 1858 24783 1914 24792
rect 1858 24168 1914 24177
rect 1858 24103 1860 24112
rect 1912 24103 1914 24112
rect 1860 24074 1912 24080
rect 1768 23656 1820 23662
rect 1768 23598 1820 23604
rect 1780 23497 1808 23598
rect 1766 23488 1822 23497
rect 1766 23423 1822 23432
rect 1860 23044 1912 23050
rect 1860 22986 1912 22992
rect 1872 22817 1900 22986
rect 1858 22808 1914 22817
rect 1858 22743 1914 22752
rect 1768 22568 1820 22574
rect 1768 22510 1820 22516
rect 1780 22137 1808 22510
rect 1766 22128 1822 22137
rect 1766 22063 1822 22072
rect 1860 21480 1912 21486
rect 1858 21448 1860 21457
rect 1912 21448 1914 21457
rect 1858 21383 1914 21392
rect 1860 20868 1912 20874
rect 1860 20810 1912 20816
rect 1872 20777 1900 20810
rect 1858 20768 1914 20777
rect 1858 20703 1914 20712
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 1780 20097 1808 20334
rect 1766 20088 1822 20097
rect 1766 20023 1822 20032
rect 1492 19848 1544 19854
rect 1492 19790 1544 19796
rect 1504 6914 1532 19790
rect 1860 19780 1912 19786
rect 1860 19722 1912 19728
rect 1872 19417 1900 19722
rect 1858 19408 1914 19417
rect 1858 19343 1914 19352
rect 1952 18760 2004 18766
rect 1858 18728 1914 18737
rect 1952 18702 2004 18708
rect 1858 18663 1860 18672
rect 1912 18663 1914 18672
rect 1860 18634 1912 18640
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1780 18057 1808 18158
rect 1766 18048 1822 18057
rect 1766 17983 1822 17992
rect 1860 17604 1912 17610
rect 1860 17546 1912 17552
rect 1872 17377 1900 17546
rect 1858 17368 1914 17377
rect 1858 17303 1914 17312
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 1780 16697 1808 17070
rect 1766 16688 1822 16697
rect 1766 16623 1822 16632
rect 1768 16040 1820 16046
rect 1766 16008 1768 16017
rect 1820 16008 1822 16017
rect 1766 15943 1822 15952
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1872 15337 1900 15370
rect 1858 15328 1914 15337
rect 1858 15263 1914 15272
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1780 14657 1808 14894
rect 1766 14648 1822 14657
rect 1766 14583 1822 14592
rect 1860 14340 1912 14346
rect 1860 14282 1912 14288
rect 1872 13977 1900 14282
rect 1858 13968 1914 13977
rect 1858 13903 1914 13912
rect 1584 13320 1636 13326
rect 1860 13320 1912 13326
rect 1584 13262 1636 13268
rect 1858 13288 1860 13297
rect 1912 13288 1914 13297
rect 1596 12986 1624 13262
rect 1858 13223 1914 13232
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1780 12617 1808 12718
rect 1766 12608 1822 12617
rect 1766 12543 1822 12552
rect 1860 12164 1912 12170
rect 1860 12106 1912 12112
rect 1872 11937 1900 12106
rect 1858 11928 1914 11937
rect 1858 11863 1914 11872
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1780 11257 1808 11630
rect 1766 11248 1822 11257
rect 1766 11183 1822 11192
rect 1768 10600 1820 10606
rect 1766 10568 1768 10577
rect 1820 10568 1822 10577
rect 1766 10503 1822 10512
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1872 9897 1900 9930
rect 1858 9888 1914 9897
rect 1858 9823 1914 9832
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1780 9217 1808 9454
rect 1766 9208 1822 9217
rect 1766 9143 1822 9152
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8537 1900 8842
rect 1858 8528 1914 8537
rect 1858 8463 1914 8472
rect 1858 7848 1914 7857
rect 1858 7783 1860 7792
rect 1912 7783 1914 7792
rect 1860 7754 1912 7760
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1780 7177 1808 7278
rect 1766 7168 1822 7177
rect 1766 7103 1822 7112
rect 1504 6886 1624 6914
rect 1596 5953 1624 6886
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1872 6497 1900 6666
rect 1858 6488 1914 6497
rect 1858 6423 1914 6432
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1582 5944 1638 5953
rect 1582 5879 1638 5888
rect 1780 5817 1808 6190
rect 1766 5808 1822 5817
rect 1766 5743 1822 5752
rect 1964 5681 1992 18702
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 2056 6769 2084 17614
rect 2148 17270 2176 37062
rect 2332 36242 2360 37810
rect 2412 37188 2464 37194
rect 2412 37130 2464 37136
rect 2424 37097 2452 37130
rect 2410 37088 2466 37097
rect 2410 37023 2466 37032
rect 2320 36236 2372 36242
rect 2320 36178 2372 36184
rect 2516 35894 2544 37810
rect 2596 36236 2648 36242
rect 2596 36178 2648 36184
rect 2424 35866 2544 35894
rect 2228 35828 2280 35834
rect 2228 35770 2280 35776
rect 2240 35086 2268 35770
rect 2424 35698 2452 35866
rect 2412 35692 2464 35698
rect 2412 35634 2464 35640
rect 2424 35086 2452 35634
rect 2228 35080 2280 35086
rect 2228 35022 2280 35028
rect 2412 35080 2464 35086
rect 2412 35022 2464 35028
rect 2320 35012 2372 35018
rect 2320 34954 2372 34960
rect 2332 32502 2360 34954
rect 2320 32496 2372 32502
rect 2320 32438 2372 32444
rect 2424 32314 2452 35022
rect 2240 32286 2452 32314
rect 2240 27470 2268 32286
rect 2504 28552 2556 28558
rect 2504 28494 2556 28500
rect 2516 28082 2544 28494
rect 2504 28076 2556 28082
rect 2504 28018 2556 28024
rect 2228 27464 2280 27470
rect 2228 27406 2280 27412
rect 2136 17264 2188 17270
rect 2136 17206 2188 17212
rect 2240 16658 2268 27406
rect 2516 27402 2544 28018
rect 2504 27396 2556 27402
rect 2504 27338 2556 27344
rect 2516 26994 2544 27338
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 2516 26382 2544 26930
rect 2608 26382 2636 36178
rect 2700 35630 2728 37862
rect 3700 37810 3752 37816
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 2688 35624 2740 35630
rect 2688 35566 2740 35572
rect 4712 35488 4764 35494
rect 4712 35430 4764 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4724 35290 4752 35430
rect 4712 35284 4764 35290
rect 4712 35226 4764 35232
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 5736 34134 5764 51750
rect 5724 34128 5776 34134
rect 5724 34070 5776 34076
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 6196 29714 6224 61270
rect 6748 61198 6776 63200
rect 7576 61198 7604 63294
rect 8206 63200 8262 64000
rect 8942 63322 8998 64000
rect 8942 63294 9168 63322
rect 8942 63200 8998 63294
rect 6736 61192 6788 61198
rect 6736 61134 6788 61140
rect 7564 61192 7616 61198
rect 7840 61192 7892 61198
rect 7564 61134 7616 61140
rect 7838 61160 7840 61169
rect 7892 61160 7894 61169
rect 7656 61124 7708 61130
rect 7838 61095 7894 61104
rect 7656 61066 7708 61072
rect 6920 61056 6972 61062
rect 6920 60998 6972 61004
rect 6932 30938 6960 60998
rect 6920 30932 6972 30938
rect 6920 30874 6972 30880
rect 6184 29708 6236 29714
rect 6184 29650 6236 29656
rect 2872 29164 2924 29170
rect 2872 29106 2924 29112
rect 2884 28694 2912 29106
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 2872 28688 2924 28694
rect 2872 28630 2924 28636
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 2504 26376 2556 26382
rect 2504 26318 2556 26324
rect 2596 26376 2648 26382
rect 2596 26318 2648 26324
rect 2516 25430 2544 26318
rect 2688 25900 2740 25906
rect 2688 25842 2740 25848
rect 2700 25498 2728 25842
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 2688 25492 2740 25498
rect 2688 25434 2740 25440
rect 2504 25424 2556 25430
rect 2504 25366 2556 25372
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 7668 21622 7696 61066
rect 8220 60874 8248 63200
rect 8220 60846 8340 60874
rect 8312 60790 8340 60846
rect 9140 60790 9168 63294
rect 9678 63200 9734 64000
rect 10414 63322 10470 64000
rect 10244 63294 10470 63322
rect 9692 61198 9720 63200
rect 10244 61198 10272 63294
rect 10414 63200 10470 63294
rect 11150 63200 11206 64000
rect 11886 63322 11942 64000
rect 12622 63322 12678 64000
rect 13358 63322 13414 64000
rect 11886 63294 12112 63322
rect 11886 63200 11942 63294
rect 11164 61198 11192 63200
rect 9680 61192 9732 61198
rect 9680 61134 9732 61140
rect 10232 61192 10284 61198
rect 10232 61134 10284 61140
rect 11152 61192 11204 61198
rect 11152 61134 11204 61140
rect 10324 61056 10376 61062
rect 10324 60998 10376 61004
rect 11980 61056 12032 61062
rect 11980 60998 12032 61004
rect 8300 60784 8352 60790
rect 8300 60726 8352 60732
rect 9128 60784 9180 60790
rect 9128 60726 9180 60732
rect 8576 60580 8628 60586
rect 8576 60522 8628 60528
rect 8588 56506 8616 60522
rect 8576 56500 8628 56506
rect 8576 56442 8628 56448
rect 9036 56364 9088 56370
rect 9036 56306 9088 56312
rect 8944 50788 8996 50794
rect 8944 50730 8996 50736
rect 8956 32910 8984 50730
rect 9048 45014 9076 56306
rect 9128 55412 9180 55418
rect 9128 55354 9180 55360
rect 9036 45008 9088 45014
rect 9036 44950 9088 44956
rect 9140 44878 9168 55354
rect 9128 44872 9180 44878
rect 9128 44814 9180 44820
rect 10336 39030 10364 60998
rect 11704 40928 11756 40934
rect 11704 40870 11756 40876
rect 11716 40730 11744 40870
rect 11704 40724 11756 40730
rect 11704 40666 11756 40672
rect 10324 39024 10376 39030
rect 10324 38966 10376 38972
rect 11704 38752 11756 38758
rect 11704 38694 11756 38700
rect 11716 37874 11744 38694
rect 11992 37942 12020 60998
rect 12084 60790 12112 63294
rect 12452 63294 12678 63322
rect 12452 61198 12480 63294
rect 12622 63200 12678 63294
rect 13280 63294 13414 63322
rect 13280 61198 13308 63294
rect 13358 63200 13414 63294
rect 14094 63322 14150 64000
rect 14094 63294 14412 63322
rect 14094 63200 14150 63294
rect 14384 61198 14412 63294
rect 14830 63200 14886 64000
rect 15566 63322 15622 64000
rect 16302 63322 16358 64000
rect 15396 63294 15622 63322
rect 12440 61192 12492 61198
rect 12440 61134 12492 61140
rect 13268 61192 13320 61198
rect 13268 61134 13320 61140
rect 14372 61192 14424 61198
rect 14372 61134 14424 61140
rect 13544 61124 13596 61130
rect 13544 61066 13596 61072
rect 12532 61056 12584 61062
rect 12532 60998 12584 61004
rect 12072 60784 12124 60790
rect 12072 60726 12124 60732
rect 12164 60512 12216 60518
rect 12164 60454 12216 60460
rect 12176 60314 12204 60454
rect 12164 60308 12216 60314
rect 12164 60250 12216 60256
rect 11980 37936 12032 37942
rect 11980 37878 12032 37884
rect 11704 37868 11756 37874
rect 11704 37810 11756 37816
rect 11336 37800 11388 37806
rect 11336 37742 11388 37748
rect 11348 37194 11376 37742
rect 11336 37188 11388 37194
rect 11336 37130 11388 37136
rect 8944 32904 8996 32910
rect 8944 32846 8996 32852
rect 7656 21616 7708 21622
rect 7656 21558 7708 21564
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 10796 18970 10824 20878
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11164 18358 11192 18770
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11256 18426 11284 18702
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 7564 18148 7616 18154
rect 7564 18090 7616 18096
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2700 7954 2728 16050
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 7576 12434 7604 18090
rect 11348 16658 11376 37130
rect 12348 36576 12400 36582
rect 12348 36518 12400 36524
rect 12360 34066 12388 36518
rect 12348 34060 12400 34066
rect 12348 34002 12400 34008
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 10508 16516 10560 16522
rect 10508 16458 10560 16464
rect 7484 12406 7604 12434
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 2042 6760 2098 6769
rect 2042 6695 2098 6704
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 1950 5672 2006 5681
rect 1950 5607 2006 5616
rect 1768 5160 1820 5166
rect 1766 5128 1768 5137
rect 1820 5128 1822 5137
rect 1766 5063 1822 5072
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 1860 4548 1912 4554
rect 1860 4490 1912 4496
rect 1872 4457 1900 4490
rect 1858 4448 1914 4457
rect 1858 4383 1914 4392
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1780 3777 1808 4014
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 1766 3768 1822 3777
rect 4214 3771 4522 3780
rect 1766 3703 1822 3712
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 1872 3097 1900 3402
rect 1858 3088 1914 3097
rect 1858 3023 1914 3032
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 1584 2440 1636 2446
rect 1860 2440 1912 2446
rect 1584 2382 1636 2388
rect 1858 2408 1860 2417
rect 1912 2408 1914 2417
rect 1596 2038 1624 2382
rect 1858 2343 1914 2352
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 1584 2032 1636 2038
rect 1584 1974 1636 1980
rect 5184 1902 5212 2246
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 5920 800 5948 3402
rect 6012 3194 6040 10474
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6932 3194 6960 4694
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6840 1426 6868 2382
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7024 1970 7052 2246
rect 7012 1964 7064 1970
rect 7012 1906 7064 1912
rect 6828 1420 6880 1426
rect 6828 1362 6880 1368
rect 7300 800 7328 4490
rect 7484 3670 7512 12406
rect 9128 11280 9180 11286
rect 9128 11222 9180 11228
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 7656 7472 7708 7478
rect 7656 7414 7708 7420
rect 7564 4480 7616 4486
rect 7564 4422 7616 4428
rect 7576 4282 7604 4422
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7668 4078 7696 7414
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 7840 4208 7892 4214
rect 7840 4150 7892 4156
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 1766 7788 2246
rect 7748 1760 7800 1766
rect 7748 1702 7800 1708
rect 7564 1420 7616 1426
rect 7564 1362 7616 1368
rect 7576 800 7604 1362
rect 7852 800 7880 4150
rect 7944 3670 7972 5102
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 3913 8340 4558
rect 8298 3904 8354 3913
rect 8298 3839 8354 3848
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8116 3120 8168 3126
rect 8116 3062 8168 3068
rect 8128 800 8156 3062
rect 8312 2774 8340 3470
rect 8404 3194 8432 10066
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8392 3188 8444 3194
rect 8392 3130 8444 3136
rect 8312 2746 8432 2774
rect 8404 800 8432 2746
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8496 1426 8524 2518
rect 8484 1420 8536 1426
rect 8484 1362 8536 1368
rect 8588 1170 8616 4490
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8772 4146 8800 4422
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8680 3670 8708 4082
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8864 3398 8892 6122
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8956 3210 8984 10134
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 8680 3182 8984 3210
rect 8680 2582 8708 3182
rect 9048 3058 9076 3878
rect 9140 3194 9168 11222
rect 10520 9722 10548 16458
rect 11256 15570 11284 16526
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11072 10810 11100 11698
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9416 3738 9444 6734
rect 9508 6322 9536 6734
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 8864 2854 8892 2994
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8588 1142 8708 1170
rect 8680 800 8708 1142
rect 8956 800 8984 2246
rect 9232 800 9260 2926
rect 9324 1562 9352 3470
rect 9416 2990 9444 3538
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 9416 2106 9444 2314
rect 9404 2100 9456 2106
rect 9404 2042 9456 2048
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 9508 800 9536 4150
rect 9600 4078 9628 4558
rect 9876 4078 9904 5170
rect 9968 4826 9996 6666
rect 10152 6118 10180 6666
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9954 3768 10010 3777
rect 9954 3703 10010 3712
rect 9968 3602 9996 3703
rect 9864 3596 9916 3602
rect 9864 3538 9916 3544
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9678 3224 9734 3233
rect 9678 3159 9680 3168
rect 9732 3159 9734 3168
rect 9680 3130 9732 3136
rect 9678 3088 9734 3097
rect 9678 3023 9680 3032
rect 9732 3023 9734 3032
rect 9680 2994 9732 3000
rect 9586 2816 9642 2825
rect 9586 2751 9642 2760
rect 9600 2514 9628 2751
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9692 1834 9720 2314
rect 9680 1828 9732 1834
rect 9680 1770 9732 1776
rect 9784 800 9812 3334
rect 9876 2990 9904 3538
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9876 1494 9904 2790
rect 9864 1488 9916 1494
rect 9864 1430 9916 1436
rect 10060 800 10088 5170
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3602 10180 3878
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10140 3052 10192 3058
rect 10244 3040 10272 4422
rect 10192 3012 10272 3040
rect 10140 2994 10192 3000
rect 10336 2774 10364 4490
rect 10152 2746 10364 2774
rect 10152 1442 10180 2746
rect 10428 2582 10456 5034
rect 10520 4078 10548 9658
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11072 6866 11100 7346
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11072 6254 11100 6666
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10704 4758 10732 5034
rect 10692 4752 10744 4758
rect 10692 4694 10744 4700
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10508 3664 10560 3670
rect 10508 3606 10560 3612
rect 10520 2582 10548 3606
rect 10704 3534 10732 4082
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10598 3224 10654 3233
rect 10598 3159 10654 3168
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10152 1414 10364 1442
rect 10336 800 10364 1414
rect 10612 800 10640 3159
rect 10704 3126 10732 3470
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10704 2514 10732 3062
rect 10796 2650 10824 4014
rect 10888 2922 10916 4150
rect 10980 4078 11008 5170
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 11072 3466 11100 6190
rect 11164 5302 11192 7958
rect 11256 6866 11284 15506
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11256 4826 11284 6802
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11164 4146 11192 4558
rect 11256 4486 11284 4762
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11348 4214 11376 16594
rect 11624 16590 11652 17206
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 12360 16454 12388 17138
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12544 16250 12572 60998
rect 13556 31754 13584 61066
rect 14464 61056 14516 61062
rect 14464 60998 14516 61004
rect 13912 38276 13964 38282
rect 13912 38218 13964 38224
rect 13924 37942 13952 38218
rect 14004 38208 14056 38214
rect 14004 38150 14056 38156
rect 14016 37942 14044 38150
rect 13912 37936 13964 37942
rect 13912 37878 13964 37884
rect 14004 37936 14056 37942
rect 14004 37878 14056 37884
rect 14476 32978 14504 60998
rect 14844 60790 14872 63200
rect 15396 61198 15424 63294
rect 15566 63200 15622 63294
rect 16132 63294 16358 63322
rect 16132 61198 16160 63294
rect 16302 63200 16358 63294
rect 17038 63322 17094 64000
rect 17774 63322 17830 64000
rect 18510 63322 18566 64000
rect 17038 63294 17264 63322
rect 17038 63200 17094 63294
rect 17132 61328 17184 61334
rect 17132 61270 17184 61276
rect 15384 61192 15436 61198
rect 15384 61134 15436 61140
rect 16120 61192 16172 61198
rect 16120 61134 16172 61140
rect 15660 61124 15712 61130
rect 15660 61066 15712 61072
rect 16396 61124 16448 61130
rect 16396 61066 16448 61072
rect 14832 60784 14884 60790
rect 14832 60726 14884 60732
rect 15108 60648 15160 60654
rect 15108 60590 15160 60596
rect 15120 58614 15148 60590
rect 15108 58608 15160 58614
rect 15108 58550 15160 58556
rect 15384 58336 15436 58342
rect 15384 58278 15436 58284
rect 15108 43648 15160 43654
rect 15108 43590 15160 43596
rect 14464 32972 14516 32978
rect 14464 32914 14516 32920
rect 13464 31726 13584 31754
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 13096 18426 13124 24142
rect 13464 22094 13492 31726
rect 14372 31680 14424 31686
rect 14372 31622 14424 31628
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 13924 23118 13952 23598
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13556 22234 13584 22578
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 13464 22066 13584 22094
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13372 21690 13400 21966
rect 13360 21684 13412 21690
rect 13360 21626 13412 21632
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12360 12442 12388 12786
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13004 11898 13032 12174
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11808 8634 11836 8910
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 12176 8430 12204 9454
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12544 8430 12572 9386
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 11992 8294 12020 8366
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11808 7546 11836 7822
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11992 7410 12020 8230
rect 12176 7818 12204 8366
rect 12268 8090 12296 8366
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11532 6458 11560 6734
rect 12268 6458 12296 7278
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11336 4208 11388 4214
rect 11336 4150 11388 4156
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 10876 2916 10928 2922
rect 10876 2858 10928 2864
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 10876 1556 10928 1562
rect 10876 1498 10928 1504
rect 10888 800 10916 1498
rect 11152 1420 11204 1426
rect 11152 1362 11204 1368
rect 11164 800 11192 1362
rect 11440 800 11468 4014
rect 11532 1970 11560 6122
rect 11624 4826 11652 6326
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11624 4078 11652 4626
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 11610 3496 11666 3505
rect 11610 3431 11666 3440
rect 11624 3398 11652 3431
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11520 1964 11572 1970
rect 11520 1906 11572 1912
rect 11716 800 11744 5578
rect 12360 5370 12388 6190
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11992 4622 12020 4762
rect 12360 4622 12388 5306
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 11992 3534 12020 4558
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11900 3126 11928 3334
rect 12084 3210 12112 4558
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12360 4146 12388 4422
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 11992 3194 12112 3210
rect 11980 3188 12112 3194
rect 12032 3182 12112 3188
rect 11980 3130 12032 3136
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 12268 2990 12296 3674
rect 12452 3670 12480 4490
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12360 3097 12388 3606
rect 12346 3088 12402 3097
rect 12346 3023 12402 3032
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 11978 2816 12034 2825
rect 11978 2751 12034 2760
rect 11992 800 12020 2751
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12256 1488 12308 1494
rect 12256 1430 12308 1436
rect 12268 800 12296 1430
rect 12452 1426 12480 2314
rect 12440 1420 12492 1426
rect 12440 1362 12492 1368
rect 12544 800 12572 5578
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12636 2854 12664 4150
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12728 2394 12756 9386
rect 12820 5098 12848 11154
rect 13096 10674 13124 17478
rect 13556 17241 13584 22066
rect 13728 21616 13780 21622
rect 13728 21558 13780 21564
rect 13740 20806 13768 21558
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13542 17232 13598 17241
rect 13542 17167 13598 17176
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 10062 12940 10406
rect 13004 10062 13032 10542
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 13004 5846 13032 9386
rect 13096 8566 13124 10610
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 13096 5914 13124 7210
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 12992 5840 13044 5846
rect 12992 5782 13044 5788
rect 12808 5092 12860 5098
rect 12808 5034 12860 5040
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12636 2366 12756 2394
rect 12636 1766 12664 2366
rect 12716 2100 12768 2106
rect 12716 2042 12768 2048
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 12728 1170 12756 2042
rect 12820 1970 12848 4014
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 12808 1964 12860 1970
rect 12808 1906 12860 1912
rect 12728 1142 12848 1170
rect 12820 800 12848 1142
rect 13096 800 13124 3878
rect 13188 2582 13216 14826
rect 13832 14822 13860 14894
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13832 12442 13860 14758
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13832 12306 13860 12378
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13280 11830 13308 12174
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13360 10600 13412 10606
rect 13360 10542 13412 10548
rect 13372 9518 13400 10542
rect 13464 10266 13492 11630
rect 13556 11354 13584 12174
rect 13832 11762 13860 12242
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13924 9081 13952 14350
rect 14016 12434 14044 15438
rect 14016 12406 14136 12434
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 9994 14044 10610
rect 14004 9988 14056 9994
rect 14004 9930 14056 9936
rect 14016 9654 14044 9930
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 13910 9072 13966 9081
rect 13910 9007 13966 9016
rect 14108 8945 14136 12406
rect 14094 8936 14150 8945
rect 14094 8871 14150 8880
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13280 7546 13308 8366
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13280 6798 13308 7346
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13280 6390 13308 6734
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13280 5166 13308 6326
rect 13556 5846 13584 6802
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13360 5636 13412 5642
rect 13360 5578 13412 5584
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 13280 3942 13308 5102
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13280 3602 13308 3878
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13372 800 13400 5578
rect 13832 5302 13860 6802
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13542 2952 13598 2961
rect 13542 2887 13544 2896
rect 13596 2887 13598 2896
rect 13544 2858 13596 2864
rect 13648 800 13676 5170
rect 13924 4146 13952 8298
rect 14004 6860 14056 6866
rect 14004 6802 14056 6808
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13726 4040 13782 4049
rect 13726 3975 13728 3984
rect 13780 3975 13782 3984
rect 13820 4004 13872 4010
rect 13728 3946 13780 3952
rect 13820 3946 13872 3952
rect 13726 3632 13782 3641
rect 13726 3567 13728 3576
rect 13780 3567 13782 3576
rect 13728 3538 13780 3544
rect 13832 3058 13860 3946
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 14016 2310 14044 6802
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14108 3942 14136 4014
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14004 2304 14056 2310
rect 14004 2246 14056 2252
rect 13912 1420 13964 1426
rect 13912 1362 13964 1368
rect 13924 800 13952 1362
rect 14200 800 14228 5578
rect 14292 3058 14320 22170
rect 14384 22030 14412 31622
rect 15120 22094 15148 43590
rect 15396 35018 15424 58278
rect 15672 56438 15700 61066
rect 16028 60580 16080 60586
rect 16028 60522 16080 60528
rect 15752 56772 15804 56778
rect 15752 56714 15804 56720
rect 15660 56432 15712 56438
rect 15660 56374 15712 56380
rect 15764 56370 15792 56714
rect 15568 56364 15620 56370
rect 15568 56306 15620 56312
rect 15752 56364 15804 56370
rect 15752 56306 15804 56312
rect 15580 52018 15608 56306
rect 15568 52012 15620 52018
rect 15568 51954 15620 51960
rect 15476 44192 15528 44198
rect 15476 44134 15528 44140
rect 15488 43858 15516 44134
rect 15476 43852 15528 43858
rect 15476 43794 15528 43800
rect 16040 43790 16068 60522
rect 16028 43784 16080 43790
rect 16028 43726 16080 43732
rect 16408 35154 16436 61066
rect 16580 61056 16632 61062
rect 16580 60998 16632 61004
rect 16592 58410 16620 60998
rect 16672 58608 16724 58614
rect 17144 58596 17172 61270
rect 17236 61198 17264 63294
rect 17774 63294 17908 63322
rect 17774 63200 17830 63294
rect 17224 61192 17276 61198
rect 17880 61180 17908 63294
rect 18510 63294 18736 63322
rect 18510 63200 18566 63294
rect 18708 61198 18736 63294
rect 19246 63200 19302 64000
rect 19982 63322 20038 64000
rect 19812 63294 20038 63322
rect 17960 61192 18012 61198
rect 17880 61152 17960 61180
rect 17224 61134 17276 61140
rect 17960 61134 18012 61140
rect 18696 61192 18748 61198
rect 18696 61134 18748 61140
rect 18144 61124 18196 61130
rect 18144 61066 18196 61072
rect 17224 58608 17276 58614
rect 16672 58550 16724 58556
rect 16762 58576 16818 58585
rect 16580 58404 16632 58410
rect 16580 58346 16632 58352
rect 16684 58138 16712 58550
rect 17144 58568 17224 58596
rect 17224 58550 17276 58556
rect 17406 58576 17462 58585
rect 16762 58511 16764 58520
rect 16816 58511 16818 58520
rect 17406 58511 17408 58520
rect 16764 58482 16816 58488
rect 17460 58511 17462 58520
rect 17408 58482 17460 58488
rect 16856 58472 16908 58478
rect 17224 58472 17276 58478
rect 16908 58420 17224 58426
rect 16856 58414 17276 58420
rect 16868 58398 17264 58414
rect 17500 58336 17552 58342
rect 17500 58278 17552 58284
rect 16672 58132 16724 58138
rect 16672 58074 16724 58080
rect 17132 58132 17184 58138
rect 17132 58074 17184 58080
rect 17144 56778 17172 58074
rect 17132 56772 17184 56778
rect 17132 56714 17184 56720
rect 16580 48000 16632 48006
rect 16580 47942 16632 47948
rect 16592 39574 16620 47942
rect 17224 47048 17276 47054
rect 17224 46990 17276 46996
rect 16580 39568 16632 39574
rect 16580 39510 16632 39516
rect 17236 37874 17264 46990
rect 17224 37868 17276 37874
rect 17224 37810 17276 37816
rect 16764 36644 16816 36650
rect 16764 36586 16816 36592
rect 16396 35148 16448 35154
rect 16396 35090 16448 35096
rect 16212 35080 16264 35086
rect 16212 35022 16264 35028
rect 16304 35080 16356 35086
rect 16304 35022 16356 35028
rect 15384 35012 15436 35018
rect 15384 34954 15436 34960
rect 15844 34944 15896 34950
rect 15844 34886 15896 34892
rect 15856 34746 15884 34886
rect 15844 34740 15896 34746
rect 15844 34682 15896 34688
rect 16224 34610 16252 35022
rect 16212 34604 16264 34610
rect 16212 34546 16264 34552
rect 16316 30598 16344 35022
rect 16488 31952 16540 31958
rect 16488 31894 16540 31900
rect 16304 30592 16356 30598
rect 16304 30534 16356 30540
rect 15200 29640 15252 29646
rect 15200 29582 15252 29588
rect 15212 25362 15240 29582
rect 16304 28688 16356 28694
rect 16304 28630 16356 28636
rect 15200 25356 15252 25362
rect 15200 25298 15252 25304
rect 15212 24818 15240 25298
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 15028 22066 15148 22094
rect 14372 22024 14424 22030
rect 14372 21966 14424 21972
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14752 18154 14780 19178
rect 14936 18834 14964 19246
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14936 18290 14964 18770
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14752 17134 14780 18090
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14752 16658 14780 17070
rect 14844 16794 14872 17818
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 14740 16652 14792 16658
rect 14740 16594 14792 16600
rect 14936 16590 14964 18226
rect 14924 16584 14976 16590
rect 14844 16532 14924 16538
rect 14844 16526 14976 16532
rect 14844 16510 14964 16526
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14660 13870 14688 14894
rect 14844 14822 14872 16510
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14936 15162 14964 16390
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14936 14074 14964 14894
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 14660 13394 14688 13806
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14660 12850 14688 13330
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 15028 11801 15056 22066
rect 15212 21554 15240 23734
rect 15580 23730 15608 24754
rect 15568 23724 15620 23730
rect 15568 23666 15620 23672
rect 15580 21690 15608 23666
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15948 21894 15976 23054
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15948 21622 15976 21830
rect 15936 21616 15988 21622
rect 15936 21558 15988 21564
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15212 21026 15240 21490
rect 15212 20998 15608 21026
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15120 19514 15148 20402
rect 15212 20058 15240 20878
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 15580 18222 15608 20998
rect 15672 20534 15700 21490
rect 15948 21010 15976 21558
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 15936 21004 15988 21010
rect 15936 20946 15988 20952
rect 15660 20528 15712 20534
rect 15660 20470 15712 20476
rect 16040 20398 16068 21422
rect 16028 20392 16080 20398
rect 16028 20334 16080 20340
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15948 19854 15976 20198
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15844 18692 15896 18698
rect 15844 18634 15896 18640
rect 15856 18290 15884 18634
rect 16132 18358 16160 24754
rect 16212 21888 16264 21894
rect 16212 21830 16264 21836
rect 16224 21622 16252 21830
rect 16212 21616 16264 21622
rect 16212 21558 16264 21564
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16224 18766 16252 18906
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16120 18352 16172 18358
rect 16120 18294 16172 18300
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15120 12782 15148 15302
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15014 11792 15070 11801
rect 15014 11727 15070 11736
rect 15212 11676 15240 16934
rect 14936 11648 15240 11676
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14384 2582 14412 3946
rect 14476 3670 14504 5510
rect 14464 3664 14516 3670
rect 14464 3606 14516 3612
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14372 2576 14424 2582
rect 14372 2518 14424 2524
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 14384 1426 14412 2314
rect 14372 1420 14424 1426
rect 14372 1362 14424 1368
rect 14476 800 14504 3334
rect 14568 1834 14596 6122
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14752 4593 14780 4966
rect 14738 4584 14794 4593
rect 14738 4519 14794 4528
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14752 4146 14780 4422
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14844 3058 14872 11086
rect 14936 10606 14964 11648
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 14936 10198 14964 10542
rect 14924 10192 14976 10198
rect 14924 10134 14976 10140
rect 15212 9518 15240 10542
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15304 6866 15332 18158
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15488 14618 15516 15438
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15396 11762 15424 14418
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15580 6254 15608 18158
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15672 17338 15700 17614
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16028 16448 16080 16454
rect 16028 16390 16080 16396
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15764 11762 15792 15846
rect 16040 14414 16068 16390
rect 16224 16114 16252 16526
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15856 14074 15884 14350
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15948 11898 15976 13874
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 16040 11898 16068 12582
rect 16120 12232 16172 12238
rect 16120 12174 16172 12180
rect 16132 12102 16160 12174
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 16040 11150 16068 11834
rect 16224 11286 16252 14758
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 14924 4548 14976 4554
rect 14924 4490 14976 4496
rect 14936 4146 14964 4490
rect 15672 4146 15700 6190
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 14936 3602 14964 4082
rect 15016 3664 15068 3670
rect 15016 3606 15068 3612
rect 14924 3596 14976 3602
rect 14924 3538 14976 3544
rect 15028 3194 15056 3606
rect 15016 3188 15068 3194
rect 15016 3130 15068 3136
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14556 1828 14608 1834
rect 14556 1770 14608 1776
rect 14752 800 14780 2586
rect 15028 800 15056 2790
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 15212 2106 15240 2314
rect 15200 2100 15252 2106
rect 15200 2042 15252 2048
rect 15292 1420 15344 1426
rect 15292 1362 15344 1368
rect 15304 800 15332 1362
rect 15580 800 15608 2994
rect 15764 2446 15792 9386
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 16132 5914 16160 6122
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16132 4758 16160 5102
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15856 800 15884 4490
rect 16224 3534 16252 11222
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 16040 1170 16068 2450
rect 16316 2446 16344 28630
rect 16500 25362 16528 31894
rect 16776 31890 16804 36586
rect 17224 33992 17276 33998
rect 17224 33934 17276 33940
rect 17236 33114 17264 33934
rect 17316 33924 17368 33930
rect 17316 33866 17368 33872
rect 17328 33318 17356 33866
rect 17316 33312 17368 33318
rect 17316 33254 17368 33260
rect 17224 33108 17276 33114
rect 17224 33050 17276 33056
rect 17316 33108 17368 33114
rect 17316 33050 17368 33056
rect 17328 32994 17356 33050
rect 17236 32978 17356 32994
rect 17224 32972 17356 32978
rect 17276 32966 17356 32972
rect 17224 32914 17276 32920
rect 17224 32768 17276 32774
rect 17224 32710 17276 32716
rect 16764 31884 16816 31890
rect 16764 31826 16816 31832
rect 16488 25356 16540 25362
rect 16488 25298 16540 25304
rect 16500 24818 16528 25298
rect 17236 25294 17264 32710
rect 17408 32428 17460 32434
rect 17408 32370 17460 32376
rect 17420 31822 17448 32370
rect 17512 32026 17540 58278
rect 18156 57866 18184 61066
rect 18512 61056 18564 61062
rect 18512 60998 18564 61004
rect 18144 57860 18196 57866
rect 18144 57802 18196 57808
rect 17868 49768 17920 49774
rect 17868 49710 17920 49716
rect 17880 49230 17908 49710
rect 17868 49224 17920 49230
rect 17868 49166 17920 49172
rect 18052 40724 18104 40730
rect 18052 40666 18104 40672
rect 17960 37664 18012 37670
rect 17960 37606 18012 37612
rect 17972 35834 18000 37606
rect 17960 35828 18012 35834
rect 17960 35770 18012 35776
rect 17960 34604 18012 34610
rect 17960 34546 18012 34552
rect 17776 34060 17828 34066
rect 17776 34002 17828 34008
rect 17500 32020 17552 32026
rect 17500 31962 17552 31968
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 17500 31748 17552 31754
rect 17500 31690 17552 31696
rect 17512 30802 17540 31690
rect 17500 30796 17552 30802
rect 17500 30738 17552 30744
rect 17408 30660 17460 30666
rect 17408 30602 17460 30608
rect 17224 25288 17276 25294
rect 17224 25230 17276 25236
rect 16488 24812 16540 24818
rect 16488 24754 16540 24760
rect 16856 24132 16908 24138
rect 16856 24074 16908 24080
rect 16868 22234 16896 24074
rect 17316 22772 17368 22778
rect 17316 22714 17368 22720
rect 16856 22228 16908 22234
rect 16856 22170 16908 22176
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16592 20942 16620 21830
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16684 20602 16712 21966
rect 16948 21412 17000 21418
rect 16948 21354 17000 21360
rect 16672 20596 16724 20602
rect 16672 20538 16724 20544
rect 16960 20398 16988 21354
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16396 19304 16448 19310
rect 16396 19246 16448 19252
rect 16408 4010 16436 19246
rect 17052 18630 17080 20742
rect 17224 18896 17276 18902
rect 17224 18838 17276 18844
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16868 18426 16896 18566
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16960 17338 16988 18158
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16794 16712 16934
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16592 16182 16620 16458
rect 16580 16176 16632 16182
rect 16580 16118 16632 16124
rect 16684 15366 16712 16526
rect 16764 16516 16816 16522
rect 16764 16458 16816 16464
rect 16776 16250 16804 16458
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 13326 16620 14758
rect 16776 13433 16804 14962
rect 16762 13424 16818 13433
rect 16762 13359 16818 13368
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16684 12238 16712 12378
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16500 11898 16528 12038
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16500 3058 16528 8842
rect 16868 8022 16896 16050
rect 16960 8090 16988 17274
rect 17052 17202 17080 18566
rect 17144 18290 17172 18702
rect 17236 18630 17264 18838
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17328 18290 17356 22714
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17144 17610 17172 18226
rect 17420 17678 17448 30602
rect 17512 30326 17540 30738
rect 17788 30666 17816 34002
rect 17868 33992 17920 33998
rect 17868 33934 17920 33940
rect 17880 32910 17908 33934
rect 17972 33930 18000 34546
rect 17960 33924 18012 33930
rect 17960 33866 18012 33872
rect 17972 33454 18000 33866
rect 17960 33448 18012 33454
rect 17960 33390 18012 33396
rect 17960 33312 18012 33318
rect 17960 33254 18012 33260
rect 17972 32910 18000 33254
rect 17868 32904 17920 32910
rect 17868 32846 17920 32852
rect 17960 32904 18012 32910
rect 17960 32846 18012 32852
rect 17880 32502 17908 32846
rect 17972 32570 18000 32846
rect 18064 32774 18092 40666
rect 18420 36916 18472 36922
rect 18420 36858 18472 36864
rect 18328 32904 18380 32910
rect 18328 32846 18380 32852
rect 18052 32768 18104 32774
rect 18052 32710 18104 32716
rect 17960 32564 18012 32570
rect 17960 32506 18012 32512
rect 17868 32496 17920 32502
rect 17868 32438 17920 32444
rect 17880 31754 17908 32438
rect 17972 31890 18000 32506
rect 18236 32360 18288 32366
rect 18236 32302 18288 32308
rect 17960 31884 18012 31890
rect 17960 31826 18012 31832
rect 17880 31726 18000 31754
rect 17972 31414 18000 31726
rect 18144 31748 18196 31754
rect 18144 31690 18196 31696
rect 17960 31408 18012 31414
rect 17960 31350 18012 31356
rect 17972 30870 18000 31350
rect 18156 31346 18184 31690
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 17960 30864 18012 30870
rect 17960 30806 18012 30812
rect 17776 30660 17828 30666
rect 17776 30602 17828 30608
rect 18156 30598 18184 31282
rect 18144 30592 18196 30598
rect 18144 30534 18196 30540
rect 17500 30320 17552 30326
rect 17500 30262 17552 30268
rect 17868 30320 17920 30326
rect 17868 30262 17920 30268
rect 17684 29708 17736 29714
rect 17684 29650 17736 29656
rect 17592 26852 17644 26858
rect 17592 26794 17644 26800
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17512 22778 17540 24142
rect 17604 23798 17632 26794
rect 17696 24206 17724 29650
rect 17880 29646 17908 30262
rect 17868 29640 17920 29646
rect 17868 29582 17920 29588
rect 18144 29096 18196 29102
rect 18144 29038 18196 29044
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 17972 27606 18000 28018
rect 18052 27668 18104 27674
rect 18052 27610 18104 27616
rect 17960 27600 18012 27606
rect 17960 27542 18012 27548
rect 17972 27470 18000 27542
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17868 27328 17920 27334
rect 17868 27270 17920 27276
rect 17880 26994 17908 27270
rect 18064 27062 18092 27610
rect 18052 27056 18104 27062
rect 18052 26998 18104 27004
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 17684 24200 17736 24206
rect 17684 24142 17736 24148
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 17592 23792 17644 23798
rect 17592 23734 17644 23740
rect 17788 23730 17816 24074
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 17592 23180 17644 23186
rect 17592 23122 17644 23128
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17500 22636 17552 22642
rect 17500 22578 17552 22584
rect 17512 18766 17540 22578
rect 17604 19378 17632 23122
rect 17776 23044 17828 23050
rect 17776 22986 17828 22992
rect 17684 22636 17736 22642
rect 17684 22578 17736 22584
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17696 18834 17724 22578
rect 17788 21146 17816 22986
rect 17880 22642 17908 26930
rect 18156 23730 18184 29038
rect 18248 28558 18276 32302
rect 18340 31754 18368 32846
rect 18432 32366 18460 36858
rect 18524 35698 18552 60998
rect 19260 60772 19288 63200
rect 19812 61198 19840 63294
rect 19982 63200 20038 63294
rect 20718 63200 20774 64000
rect 21454 63322 21510 64000
rect 21284 63294 21510 63322
rect 20732 61198 20760 63200
rect 21284 61198 21312 63294
rect 21454 63200 21510 63294
rect 22190 63322 22246 64000
rect 22926 63322 22982 64000
rect 23662 63322 23718 64000
rect 24398 63322 24454 64000
rect 22190 63294 22416 63322
rect 22190 63200 22246 63294
rect 21732 61328 21784 61334
rect 21732 61270 21784 61276
rect 19800 61192 19852 61198
rect 19800 61134 19852 61140
rect 20720 61192 20772 61198
rect 20720 61134 20772 61140
rect 21272 61192 21324 61198
rect 21272 61134 21324 61140
rect 20352 61124 20404 61130
rect 20352 61066 20404 61072
rect 19574 60956 19882 60965
rect 19574 60954 19580 60956
rect 19636 60954 19660 60956
rect 19716 60954 19740 60956
rect 19796 60954 19820 60956
rect 19876 60954 19882 60956
rect 19636 60902 19638 60954
rect 19818 60902 19820 60954
rect 19574 60900 19580 60902
rect 19636 60900 19660 60902
rect 19716 60900 19740 60902
rect 19796 60900 19820 60902
rect 19876 60900 19882 60902
rect 19574 60891 19882 60900
rect 19340 60784 19392 60790
rect 19260 60744 19340 60772
rect 19340 60726 19392 60732
rect 19574 59868 19882 59877
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59803 19882 59812
rect 19574 58780 19882 58789
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58715 19882 58724
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 20168 57452 20220 57458
rect 20168 57394 20220 57400
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 18604 53440 18656 53446
rect 18604 53382 18656 53388
rect 18616 41070 18644 53382
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19340 53168 19392 53174
rect 19340 53110 19392 53116
rect 18604 41064 18656 41070
rect 18604 41006 18656 41012
rect 18880 38412 18932 38418
rect 18880 38354 18932 38360
rect 18892 37874 18920 38354
rect 18880 37868 18932 37874
rect 18880 37810 18932 37816
rect 18972 37868 19024 37874
rect 18972 37810 19024 37816
rect 18788 37732 18840 37738
rect 18788 37674 18840 37680
rect 18604 36168 18656 36174
rect 18604 36110 18656 36116
rect 18512 35692 18564 35698
rect 18512 35634 18564 35640
rect 18616 35630 18644 36110
rect 18800 35698 18828 37674
rect 18892 37670 18920 37810
rect 18880 37664 18932 37670
rect 18880 37606 18932 37612
rect 18984 37398 19012 37810
rect 18972 37392 19024 37398
rect 18972 37334 19024 37340
rect 18788 35692 18840 35698
rect 18788 35634 18840 35640
rect 18604 35624 18656 35630
rect 18656 35572 18736 35578
rect 18604 35566 18736 35572
rect 18616 35550 18736 35566
rect 18708 35018 18736 35550
rect 18696 35012 18748 35018
rect 18696 34954 18748 34960
rect 18708 34542 18736 34954
rect 18696 34536 18748 34542
rect 18696 34478 18748 34484
rect 18420 32360 18472 32366
rect 18420 32302 18472 32308
rect 18328 31748 18380 31754
rect 18328 31690 18380 31696
rect 18328 30728 18380 30734
rect 18328 30670 18380 30676
rect 18340 30258 18368 30670
rect 18328 30252 18380 30258
rect 18328 30194 18380 30200
rect 18420 29164 18472 29170
rect 18420 29106 18472 29112
rect 18328 29096 18380 29102
rect 18328 29038 18380 29044
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18236 26920 18288 26926
rect 18236 26862 18288 26868
rect 18144 23724 18196 23730
rect 18144 23666 18196 23672
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 18248 22574 18276 26862
rect 18340 26382 18368 29038
rect 18432 28966 18460 29106
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 18432 27538 18460 28902
rect 18420 27532 18472 27538
rect 18420 27474 18472 27480
rect 18604 27396 18656 27402
rect 18604 27338 18656 27344
rect 18616 27062 18644 27338
rect 18604 27056 18656 27062
rect 18604 26998 18656 27004
rect 18616 26450 18644 26998
rect 18604 26444 18656 26450
rect 18604 26386 18656 26392
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18236 22568 18288 22574
rect 18236 22510 18288 22516
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17972 21554 18000 22374
rect 18248 22094 18276 22510
rect 18156 22066 18276 22094
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 18156 21162 18184 22066
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 17972 21134 18184 21162
rect 17868 20460 17920 20466
rect 17868 20402 17920 20408
rect 17880 20330 17908 20402
rect 17868 20324 17920 20330
rect 17868 20266 17920 20272
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17788 19446 17816 19926
rect 17880 19786 17908 20266
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17776 19440 17828 19446
rect 17776 19382 17828 19388
rect 17972 18970 18000 21134
rect 18340 21026 18368 26318
rect 18708 22094 18736 34478
rect 19352 33998 19380 53110
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 20076 48748 20128 48754
rect 20076 48690 20128 48696
rect 19984 48612 20036 48618
rect 19984 48554 20036 48560
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19432 44872 19484 44878
rect 19432 44814 19484 44820
rect 19340 33992 19392 33998
rect 19340 33934 19392 33940
rect 18972 33856 19024 33862
rect 18972 33798 19024 33804
rect 19340 33856 19392 33862
rect 19340 33798 19392 33804
rect 18880 33516 18932 33522
rect 18880 33458 18932 33464
rect 18788 32904 18840 32910
rect 18788 32846 18840 32852
rect 18800 32570 18828 32846
rect 18788 32564 18840 32570
rect 18788 32506 18840 32512
rect 18800 32434 18828 32506
rect 18788 32428 18840 32434
rect 18788 32370 18840 32376
rect 18892 30870 18920 33458
rect 18984 32978 19012 33798
rect 19064 33652 19116 33658
rect 19064 33594 19116 33600
rect 18972 32972 19024 32978
rect 18972 32914 19024 32920
rect 19076 32230 19104 33594
rect 19352 32910 19380 33798
rect 19444 33522 19472 44814
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19708 37868 19760 37874
rect 19708 37810 19760 37816
rect 19720 37777 19748 37810
rect 19706 37768 19762 37777
rect 19706 37703 19762 37712
rect 19708 37664 19760 37670
rect 19708 37606 19760 37612
rect 19720 37262 19748 37606
rect 19708 37256 19760 37262
rect 19708 37198 19760 37204
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 19432 33312 19484 33318
rect 19432 33254 19484 33260
rect 19340 32904 19392 32910
rect 19340 32846 19392 32852
rect 19444 32774 19472 33254
rect 19522 33144 19578 33153
rect 19522 33079 19578 33088
rect 19536 32842 19564 33079
rect 19616 33040 19668 33046
rect 19614 33008 19616 33017
rect 19668 33008 19670 33017
rect 19614 32943 19670 32952
rect 19890 33008 19946 33017
rect 19890 32943 19946 32952
rect 19904 32842 19932 32943
rect 19524 32836 19576 32842
rect 19524 32778 19576 32784
rect 19892 32836 19944 32842
rect 19892 32778 19944 32784
rect 19340 32768 19392 32774
rect 19338 32736 19340 32745
rect 19432 32768 19484 32774
rect 19392 32736 19394 32745
rect 19432 32710 19484 32716
rect 19338 32671 19394 32680
rect 19340 32564 19392 32570
rect 19340 32506 19392 32512
rect 19248 32360 19300 32366
rect 19248 32302 19300 32308
rect 19064 32224 19116 32230
rect 19064 32166 19116 32172
rect 19076 31346 19104 32166
rect 19260 31754 19288 32302
rect 19352 31890 19380 32506
rect 19444 32502 19472 32710
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19996 32570 20024 48554
rect 20088 43790 20116 48690
rect 20076 43784 20128 43790
rect 20076 43726 20128 43732
rect 20088 42770 20116 43726
rect 20076 42764 20128 42770
rect 20076 42706 20128 42712
rect 20076 35760 20128 35766
rect 20076 35702 20128 35708
rect 20088 34474 20116 35702
rect 20076 34468 20128 34474
rect 20076 34410 20128 34416
rect 20076 33856 20128 33862
rect 20076 33798 20128 33804
rect 20088 33590 20116 33798
rect 20076 33584 20128 33590
rect 20076 33526 20128 33532
rect 20074 33144 20130 33153
rect 20074 33079 20130 33088
rect 20088 32910 20116 33079
rect 20076 32904 20128 32910
rect 20076 32846 20128 32852
rect 19984 32564 20036 32570
rect 19984 32506 20036 32512
rect 19432 32496 19484 32502
rect 19432 32438 19484 32444
rect 19984 32428 20036 32434
rect 19984 32370 20036 32376
rect 19892 32360 19944 32366
rect 19892 32302 19944 32308
rect 19432 32292 19484 32298
rect 19432 32234 19484 32240
rect 19340 31884 19392 31890
rect 19340 31826 19392 31832
rect 19248 31748 19300 31754
rect 19248 31690 19300 31696
rect 19064 31340 19116 31346
rect 19064 31282 19116 31288
rect 18880 30864 18932 30870
rect 18880 30806 18932 30812
rect 18788 30592 18840 30598
rect 18788 30534 18840 30540
rect 18800 29578 18828 30534
rect 18788 29572 18840 29578
rect 18788 29514 18840 29520
rect 18800 29170 18828 29514
rect 18892 29510 18920 30806
rect 18880 29504 18932 29510
rect 18880 29446 18932 29452
rect 18788 29164 18840 29170
rect 18788 29106 18840 29112
rect 18800 27470 18828 29106
rect 19076 28966 19104 31282
rect 19352 30598 19380 31826
rect 19444 31346 19472 32234
rect 19798 32056 19854 32065
rect 19904 32026 19932 32302
rect 19798 31991 19800 32000
rect 19852 31991 19854 32000
rect 19892 32020 19944 32026
rect 19800 31962 19852 31968
rect 19892 31962 19944 31968
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19444 30734 19472 31282
rect 19996 30734 20024 32370
rect 20088 30802 20116 32846
rect 20180 31754 20208 57394
rect 20364 48822 20392 61066
rect 20812 61056 20864 61062
rect 20812 60998 20864 61004
rect 20444 60580 20496 60586
rect 20444 60522 20496 60528
rect 20456 57526 20484 60522
rect 20444 57520 20496 57526
rect 20444 57462 20496 57468
rect 20628 57452 20680 57458
rect 20628 57394 20680 57400
rect 20640 57254 20668 57394
rect 20628 57248 20680 57254
rect 20628 57190 20680 57196
rect 20640 56778 20668 57190
rect 20628 56772 20680 56778
rect 20628 56714 20680 56720
rect 20444 52012 20496 52018
rect 20444 51954 20496 51960
rect 20456 51338 20484 51954
rect 20444 51332 20496 51338
rect 20444 51274 20496 51280
rect 20456 49910 20484 51274
rect 20536 50176 20588 50182
rect 20536 50118 20588 50124
rect 20444 49904 20496 49910
rect 20444 49846 20496 49852
rect 20456 49162 20484 49846
rect 20548 49842 20576 50118
rect 20536 49836 20588 49842
rect 20536 49778 20588 49784
rect 20640 49774 20668 56714
rect 20824 49910 20852 60998
rect 21272 57928 21324 57934
rect 21272 57870 21324 57876
rect 21364 57928 21416 57934
rect 21364 57870 21416 57876
rect 21640 57928 21692 57934
rect 21640 57870 21692 57876
rect 20904 57792 20956 57798
rect 20904 57734 20956 57740
rect 20812 49904 20864 49910
rect 20812 49846 20864 49852
rect 20628 49768 20680 49774
rect 20628 49710 20680 49716
rect 20444 49156 20496 49162
rect 20444 49098 20496 49104
rect 20352 48816 20404 48822
rect 20352 48758 20404 48764
rect 20456 48686 20484 49098
rect 20640 48754 20668 49710
rect 20628 48748 20680 48754
rect 20628 48690 20680 48696
rect 20444 48680 20496 48686
rect 20444 48622 20496 48628
rect 20720 48680 20772 48686
rect 20720 48622 20772 48628
rect 20260 48544 20312 48550
rect 20260 48486 20312 48492
rect 20272 34202 20300 48486
rect 20352 47592 20404 47598
rect 20352 47534 20404 47540
rect 20364 37670 20392 47534
rect 20456 43722 20484 48622
rect 20444 43716 20496 43722
rect 20444 43658 20496 43664
rect 20628 43716 20680 43722
rect 20628 43658 20680 43664
rect 20536 39092 20588 39098
rect 20536 39034 20588 39040
rect 20444 38956 20496 38962
rect 20444 38898 20496 38904
rect 20456 37738 20484 38898
rect 20444 37732 20496 37738
rect 20444 37674 20496 37680
rect 20352 37664 20404 37670
rect 20352 37606 20404 37612
rect 20548 37346 20576 39034
rect 20640 38418 20668 43658
rect 20732 38962 20760 48622
rect 20720 38956 20772 38962
rect 20720 38898 20772 38904
rect 20732 38826 20760 38898
rect 20720 38820 20772 38826
rect 20720 38762 20772 38768
rect 20628 38412 20680 38418
rect 20628 38354 20680 38360
rect 20640 37466 20668 38354
rect 20916 37806 20944 57734
rect 21284 57458 21312 57870
rect 21376 57526 21404 57870
rect 21652 57594 21680 57870
rect 21640 57588 21692 57594
rect 21640 57530 21692 57536
rect 21364 57520 21416 57526
rect 21364 57462 21416 57468
rect 21272 57452 21324 57458
rect 21272 57394 21324 57400
rect 21548 57316 21600 57322
rect 21548 57258 21600 57264
rect 21364 56772 21416 56778
rect 21364 56714 21416 56720
rect 20996 56296 21048 56302
rect 20996 56238 21048 56244
rect 21008 38962 21036 56238
rect 21272 44872 21324 44878
rect 21272 44814 21324 44820
rect 20996 38956 21048 38962
rect 20996 38898 21048 38904
rect 21008 38282 21036 38898
rect 21088 38752 21140 38758
rect 21088 38694 21140 38700
rect 21100 38486 21128 38694
rect 21088 38480 21140 38486
rect 21088 38422 21140 38428
rect 20996 38276 21048 38282
rect 20996 38218 21048 38224
rect 20812 37800 20864 37806
rect 20812 37742 20864 37748
rect 20904 37800 20956 37806
rect 20904 37742 20956 37748
rect 20628 37460 20680 37466
rect 20628 37402 20680 37408
rect 20456 37318 20576 37346
rect 20824 37330 20852 37742
rect 21008 37618 21036 38218
rect 20916 37590 21036 37618
rect 20812 37324 20864 37330
rect 20456 36038 20484 37318
rect 20812 37266 20864 37272
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 20548 36922 20576 37198
rect 20720 37120 20772 37126
rect 20720 37062 20772 37068
rect 20536 36916 20588 36922
rect 20536 36858 20588 36864
rect 20732 36786 20760 37062
rect 20720 36780 20772 36786
rect 20720 36722 20772 36728
rect 20444 36032 20496 36038
rect 20444 35974 20496 35980
rect 20260 34196 20312 34202
rect 20260 34138 20312 34144
rect 20260 33992 20312 33998
rect 20260 33934 20312 33940
rect 20272 33522 20300 33934
rect 20352 33856 20404 33862
rect 20352 33798 20404 33804
rect 20260 33516 20312 33522
rect 20260 33458 20312 33464
rect 20272 32910 20300 33458
rect 20364 33318 20392 33798
rect 20352 33312 20404 33318
rect 20352 33254 20404 33260
rect 20350 33008 20406 33017
rect 20350 32943 20406 32952
rect 20260 32904 20312 32910
rect 20260 32846 20312 32852
rect 20260 32428 20312 32434
rect 20364 32416 20392 32943
rect 20312 32388 20392 32416
rect 20260 32370 20312 32376
rect 20456 32026 20484 35974
rect 20628 35828 20680 35834
rect 20628 35770 20680 35776
rect 20536 33652 20588 33658
rect 20536 33594 20588 33600
rect 20548 32298 20576 33594
rect 20640 32586 20668 35770
rect 20812 35692 20864 35698
rect 20812 35634 20864 35640
rect 20824 32978 20852 35634
rect 20916 34490 20944 37590
rect 21088 36848 21140 36854
rect 21088 36790 21140 36796
rect 20996 36780 21048 36786
rect 20996 36722 21048 36728
rect 21008 36106 21036 36722
rect 21100 36650 21128 36790
rect 21180 36780 21232 36786
rect 21180 36722 21232 36728
rect 21088 36644 21140 36650
rect 21088 36586 21140 36592
rect 20996 36100 21048 36106
rect 20996 36042 21048 36048
rect 21008 35766 21036 36042
rect 21192 35986 21220 36722
rect 21284 36174 21312 44814
rect 21376 38350 21404 56714
rect 21560 49230 21588 57258
rect 21744 56846 21772 61270
rect 22388 61198 22416 63294
rect 22926 63294 23152 63322
rect 22926 63200 22982 63294
rect 23124 61198 23152 63294
rect 23662 63294 23888 63322
rect 23662 63200 23718 63294
rect 23860 61198 23888 63294
rect 24398 63294 24624 63322
rect 24398 63200 24454 63294
rect 22376 61192 22428 61198
rect 22376 61134 22428 61140
rect 23112 61192 23164 61198
rect 23112 61134 23164 61140
rect 23848 61192 23900 61198
rect 23848 61134 23900 61140
rect 22284 61056 22336 61062
rect 22284 60998 22336 61004
rect 22928 61056 22980 61062
rect 22928 60998 22980 61004
rect 23940 61056 23992 61062
rect 23940 60998 23992 61004
rect 21824 60308 21876 60314
rect 21824 60250 21876 60256
rect 21836 57866 21864 60250
rect 21916 58540 21968 58546
rect 21916 58482 21968 58488
rect 21928 57916 21956 58482
rect 22008 57928 22060 57934
rect 21928 57888 22008 57916
rect 22008 57870 22060 57876
rect 21824 57860 21876 57866
rect 21824 57802 21876 57808
rect 21824 57520 21876 57526
rect 21824 57462 21876 57468
rect 21640 56840 21692 56846
rect 21640 56782 21692 56788
rect 21732 56840 21784 56846
rect 21732 56782 21784 56788
rect 21652 49434 21680 56782
rect 21836 56778 21864 57462
rect 21916 57248 21968 57254
rect 21916 57190 21968 57196
rect 21928 56846 21956 57190
rect 21916 56840 21968 56846
rect 21916 56782 21968 56788
rect 21824 56772 21876 56778
rect 21824 56714 21876 56720
rect 22020 56302 22048 57870
rect 22192 57452 22244 57458
rect 22192 57394 22244 57400
rect 22100 56976 22152 56982
rect 22100 56918 22152 56924
rect 22008 56296 22060 56302
rect 22008 56238 22060 56244
rect 22008 49632 22060 49638
rect 22008 49574 22060 49580
rect 21640 49428 21692 49434
rect 21640 49370 21692 49376
rect 21548 49224 21600 49230
rect 21548 49166 21600 49172
rect 21456 49156 21508 49162
rect 21456 49098 21508 49104
rect 21468 47666 21496 49098
rect 21560 48686 21588 49166
rect 22020 48754 22048 49574
rect 22008 48748 22060 48754
rect 22008 48690 22060 48696
rect 21548 48680 21600 48686
rect 21548 48622 21600 48628
rect 21732 48272 21784 48278
rect 21732 48214 21784 48220
rect 21456 47660 21508 47666
rect 21456 47602 21508 47608
rect 21640 46028 21692 46034
rect 21640 45970 21692 45976
rect 21548 45620 21600 45626
rect 21548 45562 21600 45568
rect 21364 38344 21416 38350
rect 21364 38286 21416 38292
rect 21456 38344 21508 38350
rect 21456 38286 21508 38292
rect 21468 37874 21496 38286
rect 21456 37868 21508 37874
rect 21456 37810 21508 37816
rect 21364 37460 21416 37466
rect 21364 37402 21416 37408
rect 21376 37194 21404 37402
rect 21364 37188 21416 37194
rect 21364 37130 21416 37136
rect 21468 36836 21496 37810
rect 21560 37262 21588 45562
rect 21652 38486 21680 45970
rect 21640 38480 21692 38486
rect 21640 38422 21692 38428
rect 21640 38344 21692 38350
rect 21640 38286 21692 38292
rect 21548 37256 21600 37262
rect 21548 37198 21600 37204
rect 21376 36808 21496 36836
rect 21272 36168 21324 36174
rect 21272 36110 21324 36116
rect 21272 36032 21324 36038
rect 21192 35980 21272 35986
rect 21192 35974 21324 35980
rect 21192 35958 21312 35974
rect 20996 35760 21048 35766
rect 20996 35702 21048 35708
rect 21284 35698 21312 35958
rect 21272 35692 21324 35698
rect 21272 35634 21324 35640
rect 20996 35624 21048 35630
rect 20996 35566 21048 35572
rect 21008 34678 21036 35566
rect 21180 34944 21232 34950
rect 21180 34886 21232 34892
rect 20996 34672 21048 34678
rect 20996 34614 21048 34620
rect 21192 34610 21220 34886
rect 21284 34678 21312 35634
rect 21272 34672 21324 34678
rect 21272 34614 21324 34620
rect 21180 34604 21232 34610
rect 21180 34546 21232 34552
rect 20916 34462 21036 34490
rect 20812 32972 20864 32978
rect 20812 32914 20864 32920
rect 20812 32836 20864 32842
rect 20812 32778 20864 32784
rect 20640 32558 20760 32586
rect 20628 32496 20680 32502
rect 20628 32438 20680 32444
rect 20536 32292 20588 32298
rect 20536 32234 20588 32240
rect 20444 32020 20496 32026
rect 20444 31962 20496 31968
rect 20548 31754 20576 32234
rect 20180 31726 20300 31754
rect 20076 30796 20128 30802
rect 20076 30738 20128 30744
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 19984 30728 20036 30734
rect 19984 30670 20036 30676
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 19444 30410 19472 30670
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19352 30382 19472 30410
rect 19616 30388 19668 30394
rect 19352 29646 19380 30382
rect 19616 30330 19668 30336
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 19156 29640 19208 29646
rect 19156 29582 19208 29588
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19168 29102 19196 29582
rect 19444 29306 19472 30126
rect 19628 30122 19656 30330
rect 19996 30190 20024 30670
rect 20088 30394 20116 30738
rect 20076 30388 20128 30394
rect 20076 30330 20128 30336
rect 20076 30252 20128 30258
rect 20076 30194 20128 30200
rect 19984 30184 20036 30190
rect 19984 30126 20036 30132
rect 19616 30116 19668 30122
rect 19616 30058 19668 30064
rect 19982 30016 20038 30025
rect 19982 29951 20038 29960
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 29300 19484 29306
rect 19432 29242 19484 29248
rect 19524 29164 19576 29170
rect 19524 29106 19576 29112
rect 19156 29096 19208 29102
rect 19536 29050 19564 29106
rect 19156 29038 19208 29044
rect 19260 29022 19564 29050
rect 19616 29096 19668 29102
rect 19616 29038 19668 29044
rect 19064 28960 19116 28966
rect 19064 28902 19116 28908
rect 18880 27600 18932 27606
rect 18880 27542 18932 27548
rect 18788 27464 18840 27470
rect 18788 27406 18840 27412
rect 18892 26330 18920 27542
rect 19260 26926 19288 29022
rect 19628 28914 19656 29038
rect 19352 28886 19656 28914
rect 19352 27538 19380 28886
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 19352 26994 19380 27474
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19340 26988 19392 26994
rect 19340 26930 19392 26936
rect 19248 26920 19300 26926
rect 19248 26862 19300 26868
rect 18064 20998 18368 21026
rect 18524 22066 18736 22094
rect 18800 26302 18920 26330
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17512 18358 17540 18702
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 18064 18290 18092 20998
rect 18144 20868 18196 20874
rect 18144 20810 18196 20816
rect 18420 20868 18472 20874
rect 18420 20810 18472 20816
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 17684 17808 17736 17814
rect 17684 17750 17736 17756
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17316 17604 17368 17610
rect 17316 17546 17368 17552
rect 17040 17196 17092 17202
rect 17328 17184 17356 17546
rect 17408 17196 17460 17202
rect 17328 17156 17408 17184
rect 17040 17138 17092 17144
rect 17408 17138 17460 17144
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17144 14793 17172 17002
rect 17314 16552 17370 16561
rect 17314 16487 17370 16496
rect 17328 16114 17356 16487
rect 17420 16250 17448 17138
rect 17500 17060 17552 17066
rect 17500 17002 17552 17008
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17512 16182 17540 17002
rect 17604 16590 17632 17750
rect 17696 17542 17724 17750
rect 18156 17678 18184 20810
rect 18236 20528 18288 20534
rect 18432 20482 18460 20810
rect 18288 20476 18460 20482
rect 18236 20470 18460 20476
rect 18248 20466 18460 20470
rect 18248 20460 18472 20466
rect 18248 20454 18420 20460
rect 18236 20324 18288 20330
rect 18236 20266 18288 20272
rect 18248 19378 18276 20266
rect 18340 19514 18368 20454
rect 18420 20402 18472 20408
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18432 19378 18460 19722
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 17960 17604 18012 17610
rect 17960 17546 18012 17552
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17500 16176 17552 16182
rect 17500 16118 17552 16124
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17604 16046 17632 16526
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17236 14958 17264 15982
rect 17696 15502 17724 17206
rect 17868 17196 17920 17202
rect 17788 17156 17868 17184
rect 17788 16590 17816 17156
rect 17868 17138 17920 17144
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17130 14784 17186 14793
rect 17130 14719 17186 14728
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17144 12442 17172 13806
rect 17236 13530 17264 14894
rect 17406 14784 17462 14793
rect 17406 14719 17462 14728
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17052 11898 17080 12242
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 17144 11218 17172 12242
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 17144 10538 17172 10678
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 16856 8016 16908 8022
rect 16856 7958 16908 7964
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 16592 3534 16620 5578
rect 16868 4146 16896 6938
rect 16946 6352 17002 6361
rect 16946 6287 16948 6296
rect 17000 6287 17002 6296
rect 16948 6258 17000 6264
rect 17144 5574 17172 8026
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 16948 4548 17000 4554
rect 16948 4490 17000 4496
rect 16856 4140 16908 4146
rect 16856 4082 16908 4088
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 16132 1766 16160 2314
rect 16120 1760 16172 1766
rect 16120 1702 16172 1708
rect 16040 1142 16160 1170
rect 16132 800 16160 1142
rect 16408 800 16436 2858
rect 16684 800 16712 3946
rect 16960 800 16988 4490
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17144 2774 17172 3538
rect 17236 3058 17264 13194
rect 17420 11830 17448 14719
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17512 11898 17540 12786
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17328 3233 17356 4014
rect 17420 3942 17448 8026
rect 17512 4146 17540 11018
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 17420 3398 17448 3606
rect 17604 3534 17632 13670
rect 17788 11898 17816 16526
rect 17972 16114 18000 17546
rect 18156 16561 18184 17614
rect 18340 17542 18368 18906
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18142 16552 18198 16561
rect 18142 16487 18198 16496
rect 18234 16144 18290 16153
rect 17960 16108 18012 16114
rect 18234 16079 18236 16088
rect 17960 16050 18012 16056
rect 18288 16079 18290 16088
rect 18236 16050 18288 16056
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17880 13258 17908 13738
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 18156 12986 18184 14826
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17972 11694 18000 12106
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17684 11620 17736 11626
rect 17684 11562 17736 11568
rect 17696 11354 17724 11562
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17788 10266 17816 10542
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17972 8838 18000 11630
rect 18340 11626 18368 17478
rect 18432 17338 18460 18022
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18524 16590 18552 22066
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18616 21146 18644 21286
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18616 19446 18644 20334
rect 18604 19440 18656 19446
rect 18604 19382 18656 19388
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18616 18834 18644 19110
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18616 18086 18644 18770
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18524 15434 18552 15846
rect 18512 15428 18564 15434
rect 18512 15370 18564 15376
rect 18524 15094 18552 15370
rect 18512 15088 18564 15094
rect 18512 15030 18564 15036
rect 18420 14884 18472 14890
rect 18420 14826 18472 14832
rect 18432 14618 18460 14826
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18512 13864 18564 13870
rect 18512 13806 18564 13812
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 18328 11620 18380 11626
rect 18328 11562 18380 11568
rect 18156 11218 18184 11562
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18064 10538 18092 10950
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 18156 8498 18184 9454
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 17960 8424 18012 8430
rect 18248 8378 18276 9114
rect 18340 8566 18368 11562
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 17960 8366 18012 8372
rect 17972 7546 18000 8366
rect 18156 8350 18276 8378
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 6458 17816 6598
rect 17866 6488 17922 6497
rect 17776 6452 17828 6458
rect 17866 6423 17868 6432
rect 17776 6394 17828 6400
rect 17920 6423 17922 6432
rect 17868 6394 17920 6400
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17314 3224 17370 3233
rect 17314 3159 17370 3168
rect 17500 3120 17552 3126
rect 17500 3062 17552 3068
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17144 2746 17264 2774
rect 17236 800 17264 2746
rect 17512 800 17540 3062
rect 17696 1902 17724 5170
rect 17684 1896 17736 1902
rect 17684 1838 17736 1844
rect 17788 800 17816 5646
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17880 3097 17908 4082
rect 17866 3088 17922 3097
rect 17866 3023 17922 3032
rect 17972 2530 18000 4966
rect 18064 4690 18092 4966
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18156 3058 18184 8350
rect 18340 7750 18368 8502
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18248 6866 18276 7686
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18248 6390 18276 6802
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18340 5370 18368 6190
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 17972 2502 18092 2530
rect 18064 800 18092 2502
rect 18340 800 18368 5034
rect 18432 4078 18460 12174
rect 18524 10742 18552 13806
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18616 11150 18644 11630
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18524 7342 18552 10542
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18524 6390 18552 7278
rect 18512 6384 18564 6390
rect 18512 6326 18564 6332
rect 18616 6254 18644 8366
rect 18708 7562 18736 18362
rect 18800 16590 18828 26302
rect 19248 25492 19300 25498
rect 19248 25434 19300 25440
rect 19260 25158 19288 25434
rect 19248 25152 19300 25158
rect 19248 25094 19300 25100
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18892 22642 18920 23122
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18984 19310 19012 19790
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 19076 17678 19104 23734
rect 19168 21554 19196 24550
rect 19260 24206 19288 25094
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 19260 23798 19288 24142
rect 19248 23792 19300 23798
rect 19248 23734 19300 23740
rect 19352 23254 19380 24754
rect 19444 24698 19472 26318
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19996 25498 20024 29951
rect 20088 26382 20116 30194
rect 20168 26988 20220 26994
rect 20168 26930 20220 26936
rect 20180 26450 20208 26930
rect 20168 26444 20220 26450
rect 20168 26386 20220 26392
rect 20076 26376 20128 26382
rect 20076 26318 20128 26324
rect 20076 25696 20128 25702
rect 20076 25638 20128 25644
rect 19984 25492 20036 25498
rect 19984 25434 20036 25440
rect 19984 25220 20036 25226
rect 19984 25162 20036 25168
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19708 24744 19760 24750
rect 19444 24670 19564 24698
rect 19708 24686 19760 24692
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19444 24274 19472 24550
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19536 24154 19564 24670
rect 19444 24126 19564 24154
rect 19340 23248 19392 23254
rect 19340 23190 19392 23196
rect 19444 23066 19472 24126
rect 19720 24070 19748 24686
rect 19708 24064 19760 24070
rect 19708 24006 19760 24012
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23866 20024 25162
rect 20088 24206 20116 25638
rect 20168 25288 20220 25294
rect 20168 25230 20220 25236
rect 20180 24818 20208 25230
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20180 24410 20208 24754
rect 20168 24404 20220 24410
rect 20168 24346 20220 24352
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19984 23860 20036 23866
rect 19984 23802 20036 23808
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 19812 23322 19840 23462
rect 19800 23316 19852 23322
rect 19800 23258 19852 23264
rect 19812 23118 19840 23258
rect 19352 23038 19472 23066
rect 19800 23112 19852 23118
rect 19800 23054 19852 23060
rect 19352 22710 19380 23038
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19444 22778 19472 22918
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19340 22704 19392 22710
rect 19340 22646 19392 22652
rect 20272 22094 20300 31726
rect 20536 31748 20588 31754
rect 20536 31690 20588 31696
rect 20548 31362 20576 31690
rect 20456 31346 20576 31362
rect 20444 31340 20576 31346
rect 20496 31334 20576 31340
rect 20444 31282 20496 31288
rect 20456 29850 20484 31282
rect 20536 31272 20588 31278
rect 20536 31214 20588 31220
rect 20548 30734 20576 31214
rect 20640 30734 20668 32438
rect 20732 31822 20760 32558
rect 20824 31822 20852 32778
rect 20902 32056 20958 32065
rect 20902 31991 20904 32000
rect 20956 31991 20958 32000
rect 20904 31962 20956 31968
rect 20720 31816 20772 31822
rect 20720 31758 20772 31764
rect 20812 31816 20864 31822
rect 20812 31758 20864 31764
rect 20536 30728 20588 30734
rect 20536 30670 20588 30676
rect 20628 30728 20680 30734
rect 20628 30670 20680 30676
rect 20536 30592 20588 30598
rect 20536 30534 20588 30540
rect 20444 29844 20496 29850
rect 20444 29786 20496 29792
rect 20456 29646 20484 29786
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20456 29238 20484 29582
rect 20444 29232 20496 29238
rect 20444 29174 20496 29180
rect 20548 27606 20576 30534
rect 20640 30326 20668 30670
rect 21008 30598 21036 34462
rect 21180 34196 21232 34202
rect 21180 34138 21232 34144
rect 21192 33590 21220 34138
rect 21180 33584 21232 33590
rect 21180 33526 21232 33532
rect 21180 32904 21232 32910
rect 21178 32872 21180 32881
rect 21232 32872 21234 32881
rect 21376 32842 21404 36808
rect 21456 36100 21508 36106
rect 21456 36042 21508 36048
rect 21468 35630 21496 36042
rect 21456 35624 21508 35630
rect 21456 35566 21508 35572
rect 21560 35154 21588 37198
rect 21652 36922 21680 38286
rect 21640 36916 21692 36922
rect 21640 36858 21692 36864
rect 21640 36576 21692 36582
rect 21640 36518 21692 36524
rect 21652 36174 21680 36518
rect 21640 36168 21692 36174
rect 21640 36110 21692 36116
rect 21548 35148 21600 35154
rect 21468 35108 21548 35136
rect 21178 32807 21234 32816
rect 21364 32836 21416 32842
rect 21364 32778 21416 32784
rect 20996 30592 21048 30598
rect 20996 30534 21048 30540
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20996 30116 21048 30122
rect 20996 30058 21048 30064
rect 21008 29646 21036 30058
rect 20996 29640 21048 29646
rect 20996 29582 21048 29588
rect 20720 29572 20772 29578
rect 20720 29514 20772 29520
rect 20536 27600 20588 27606
rect 20536 27542 20588 27548
rect 20732 27402 20760 29514
rect 21008 29034 21036 29582
rect 20996 29028 21048 29034
rect 20996 28970 21048 28976
rect 20720 27396 20772 27402
rect 20720 27338 20772 27344
rect 20732 26994 20760 27338
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 21468 26858 21496 35108
rect 21548 35090 21600 35096
rect 21640 34196 21692 34202
rect 21640 34138 21692 34144
rect 21652 34066 21680 34138
rect 21640 34060 21692 34066
rect 21640 34002 21692 34008
rect 21744 32910 21772 48214
rect 21916 39568 21968 39574
rect 21916 39510 21968 39516
rect 21824 38208 21876 38214
rect 21824 38150 21876 38156
rect 21548 32904 21600 32910
rect 21548 32846 21600 32852
rect 21732 32904 21784 32910
rect 21732 32846 21784 32852
rect 21560 31210 21588 32846
rect 21836 31754 21864 38150
rect 21928 37262 21956 39510
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 22008 35692 22060 35698
rect 22008 35634 22060 35640
rect 21916 34536 21968 34542
rect 21916 34478 21968 34484
rect 21928 32910 21956 34478
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 21652 31726 21864 31754
rect 21548 31204 21600 31210
rect 21548 31146 21600 31152
rect 21560 30802 21588 31146
rect 21548 30796 21600 30802
rect 21548 30738 21600 30744
rect 21456 26852 21508 26858
rect 21456 26794 21508 26800
rect 20536 25900 20588 25906
rect 20536 25842 20588 25848
rect 21088 25900 21140 25906
rect 21088 25842 21140 25848
rect 20444 25832 20496 25838
rect 20444 25774 20496 25780
rect 20456 25362 20484 25774
rect 20444 25356 20496 25362
rect 20444 25298 20496 25304
rect 20352 24948 20404 24954
rect 20352 24890 20404 24896
rect 20364 23168 20392 24890
rect 20456 23662 20484 25298
rect 20548 24954 20576 25842
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20536 24948 20588 24954
rect 20536 24890 20588 24896
rect 20640 23866 20668 25094
rect 21100 24070 21128 25842
rect 21272 25220 21324 25226
rect 21272 25162 21324 25168
rect 21284 24614 21312 25162
rect 21364 25152 21416 25158
rect 21364 25094 21416 25100
rect 21376 24818 21404 25094
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21180 24200 21232 24206
rect 21180 24142 21232 24148
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20444 23656 20496 23662
rect 20444 23598 20496 23604
rect 20536 23588 20588 23594
rect 20536 23530 20588 23536
rect 20548 23254 20576 23530
rect 20536 23248 20588 23254
rect 20536 23190 20588 23196
rect 20364 23140 20484 23168
rect 20456 23050 20484 23140
rect 20352 23044 20404 23050
rect 20352 22986 20404 22992
rect 20444 23044 20496 23050
rect 20444 22986 20496 22992
rect 20364 22710 20392 22986
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 20548 22574 20576 22918
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20180 22066 20300 22094
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19444 21622 19472 21966
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 21616 19484 21622
rect 19432 21558 19484 21564
rect 19156 21548 19208 21554
rect 19156 21490 19208 21496
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 19168 20466 19196 21354
rect 19352 21078 19380 21354
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 19444 20942 19472 21558
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19168 19514 19196 20198
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18880 17264 18932 17270
rect 18880 17206 18932 17212
rect 18892 17066 18920 17206
rect 18880 17060 18932 17066
rect 18880 17002 18932 17008
rect 18984 16674 19012 17478
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19064 17264 19116 17270
rect 19064 17206 19116 17212
rect 18892 16658 19012 16674
rect 18892 16652 19024 16658
rect 18892 16646 18972 16652
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18800 16114 18828 16390
rect 18892 16114 18920 16646
rect 18972 16594 19024 16600
rect 19076 16590 19104 17206
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 18984 16250 19012 16458
rect 19076 16250 19104 16526
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 18892 13462 18920 15914
rect 19168 15858 19196 17274
rect 19260 17134 19288 18362
rect 19352 17678 19380 19654
rect 19444 18834 19472 20878
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 18828 19484 18834
rect 19432 18770 19484 18776
rect 19800 18828 19852 18834
rect 19852 18788 20024 18816
rect 19800 18770 19852 18776
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19444 17134 19472 18634
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18426 20024 18788
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20076 18352 20128 18358
rect 20076 18294 20128 18300
rect 19892 17808 19944 17814
rect 19944 17768 20024 17796
rect 19892 17750 19944 17756
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19260 15978 19288 16526
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19248 15972 19300 15978
rect 19248 15914 19300 15920
rect 19168 15830 19288 15858
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19168 13938 19196 14758
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18800 11762 18828 13262
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18984 12986 19012 13126
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 19076 11558 19104 11834
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 18880 10736 18932 10742
rect 18880 10678 18932 10684
rect 18708 7534 18828 7562
rect 18696 7268 18748 7274
rect 18696 7210 18748 7216
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18616 5778 18644 6190
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18524 5166 18552 5510
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18616 4826 18644 5510
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18524 4282 18552 4422
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18708 4078 18736 7210
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18432 3534 18460 4014
rect 18696 3936 18748 3942
rect 18694 3904 18696 3913
rect 18748 3904 18750 3913
rect 18694 3839 18750 3848
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18800 2774 18828 7534
rect 18892 7274 18920 10678
rect 19168 10169 19196 11154
rect 19154 10160 19210 10169
rect 19154 10095 19210 10104
rect 18972 8424 19024 8430
rect 19168 8412 19196 10095
rect 19024 8384 19196 8412
rect 18972 8366 19024 8372
rect 19064 8288 19116 8294
rect 19062 8256 19064 8265
rect 19116 8256 19118 8265
rect 19062 8191 19118 8200
rect 19156 8016 19208 8022
rect 19156 7958 19208 7964
rect 18880 7268 18932 7274
rect 18880 7210 18932 7216
rect 19168 6322 19196 7958
rect 19260 6934 19288 15830
rect 19352 15570 19380 15982
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19352 15162 19380 15506
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19444 15065 19472 17070
rect 19904 16658 19932 17138
rect 19996 16833 20024 17768
rect 20088 17202 20116 18294
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 19982 16824 20038 16833
rect 19982 16759 20038 16768
rect 19892 16652 19944 16658
rect 19892 16594 19944 16600
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19996 15502 20024 16050
rect 19524 15496 19576 15502
rect 19522 15464 19524 15473
rect 19984 15496 20036 15502
rect 19576 15464 19578 15473
rect 19984 15438 20036 15444
rect 19522 15399 19578 15408
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20088 15178 20116 17138
rect 20180 15348 20208 22066
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 20272 17882 20300 19926
rect 20456 19922 20484 21626
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 20352 18692 20404 18698
rect 20352 18634 20404 18640
rect 20364 18426 20392 18634
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 20640 18222 20668 23802
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20732 20398 20760 21898
rect 20824 20534 20852 23054
rect 20904 23044 20956 23050
rect 20904 22986 20956 22992
rect 20916 21350 20944 22986
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 21008 20058 21036 20810
rect 20996 20052 21048 20058
rect 20996 19994 21048 20000
rect 20904 18896 20956 18902
rect 20904 18838 20956 18844
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20352 17604 20404 17610
rect 20352 17546 20404 17552
rect 20364 17202 20392 17546
rect 20456 17542 20484 18158
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20640 16590 20668 18022
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20444 16516 20496 16522
rect 20444 16458 20496 16464
rect 20180 15320 20300 15348
rect 20088 15150 20208 15178
rect 19984 15088 20036 15094
rect 19430 15056 19486 15065
rect 19340 15020 19392 15026
rect 19984 15030 20036 15036
rect 19430 14991 19486 15000
rect 19340 14962 19392 14968
rect 19352 13394 19380 14962
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19444 14414 19472 14894
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19444 13938 19472 14350
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19996 13988 20024 15030
rect 19904 13960 20024 13988
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19352 11830 19380 13330
rect 19628 13172 19656 13874
rect 19904 13190 19932 13960
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19444 13144 19656 13172
rect 19892 13184 19944 13190
rect 19444 12442 19472 13144
rect 19892 13126 19944 13132
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19892 12368 19944 12374
rect 19890 12336 19892 12345
rect 19944 12336 19946 12345
rect 19890 12271 19946 12280
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19340 11824 19392 11830
rect 19340 11766 19392 11772
rect 19444 11286 19472 11834
rect 19800 11688 19852 11694
rect 19798 11656 19800 11665
rect 19852 11656 19854 11665
rect 19996 11626 20024 13194
rect 19798 11591 19854 11600
rect 19984 11620 20036 11626
rect 19984 11562 20036 11568
rect 19432 11280 19484 11286
rect 19338 11248 19394 11257
rect 19432 11222 19484 11228
rect 19338 11183 19394 11192
rect 19248 6928 19300 6934
rect 19248 6870 19300 6876
rect 19246 6488 19302 6497
rect 19246 6423 19302 6432
rect 19260 6390 19288 6423
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19064 6180 19116 6186
rect 19064 6122 19116 6128
rect 18972 5840 19024 5846
rect 18972 5782 19024 5788
rect 18984 5642 19012 5782
rect 18972 5636 19024 5642
rect 18972 5578 19024 5584
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 18892 3670 18920 5510
rect 19076 5166 19104 6122
rect 19352 5386 19380 11183
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 9674 19472 11086
rect 19996 11014 20024 11562
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 20074 10296 20130 10305
rect 20074 10231 20130 10240
rect 20088 10198 20116 10231
rect 20076 10192 20128 10198
rect 20076 10134 20128 10140
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19444 9646 19564 9674
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 9110 19472 9318
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19432 8968 19484 8974
rect 19536 8956 19564 9646
rect 19484 8928 19564 8956
rect 19432 8910 19484 8916
rect 19444 8566 19472 8910
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19996 8634 20024 8774
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19444 7954 19472 8502
rect 19708 8288 19760 8294
rect 19708 8230 19760 8236
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19444 7546 19472 7890
rect 19616 7812 19668 7818
rect 19720 7800 19748 8230
rect 19668 7772 19748 7800
rect 19984 7812 20036 7818
rect 19616 7754 19668 7760
rect 19984 7754 20036 7760
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19798 7304 19854 7313
rect 19996 7274 20024 7754
rect 19798 7239 19800 7248
rect 19852 7239 19854 7248
rect 19984 7268 20036 7274
rect 19800 7210 19852 7216
rect 19984 7210 20036 7216
rect 20180 6866 20208 15150
rect 20272 7290 20300 15320
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20364 14074 20392 14350
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20456 13954 20484 16458
rect 20534 16416 20590 16425
rect 20534 16351 20590 16360
rect 20364 13926 20484 13954
rect 20364 11257 20392 13926
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20456 12170 20484 12582
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20350 11248 20406 11257
rect 20350 11183 20406 11192
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20364 8276 20392 11018
rect 20456 8430 20484 11290
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20364 8248 20484 8276
rect 20352 7812 20404 7818
rect 20352 7754 20404 7760
rect 20364 7410 20392 7754
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20272 7262 20392 7290
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19432 5772 19484 5778
rect 19536 5760 19564 6394
rect 19996 6390 20024 6598
rect 20088 6458 20116 6666
rect 20258 6624 20314 6633
rect 20258 6559 20314 6568
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 19484 5732 19564 5760
rect 19432 5714 19484 5720
rect 19260 5358 19380 5386
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19076 4690 19104 5102
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 19076 4146 19104 4626
rect 19154 4584 19210 4593
rect 19154 4519 19210 4528
rect 19168 4146 19196 4519
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 18972 3936 19024 3942
rect 18970 3904 18972 3913
rect 19024 3904 19026 3913
rect 18970 3839 19026 3848
rect 19076 3754 19104 4082
rect 19260 3913 19288 5358
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19246 3904 19302 3913
rect 19246 3839 19302 3848
rect 18984 3726 19104 3754
rect 19246 3768 19302 3777
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 18984 3602 19012 3726
rect 19246 3703 19302 3712
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 18972 3596 19024 3602
rect 18972 3538 19024 3544
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 18984 3369 19012 3402
rect 18970 3360 19026 3369
rect 18970 3295 19026 3304
rect 19076 3058 19104 3606
rect 19260 3534 19288 3703
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19156 3392 19208 3398
rect 19154 3360 19156 3369
rect 19208 3360 19210 3369
rect 19154 3295 19210 3304
rect 19246 3224 19302 3233
rect 19246 3159 19302 3168
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19260 2938 19288 3159
rect 19352 3126 19380 4422
rect 19444 3777 19472 5714
rect 20272 5574 20300 6559
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19798 5264 19854 5273
rect 19798 5199 19854 5208
rect 19812 4622 19840 5199
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19996 4282 20024 4422
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19430 3768 19486 3777
rect 19430 3703 19486 3712
rect 19444 3602 19472 3703
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19536 3534 19564 4218
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19720 3534 19748 3878
rect 20180 3738 20208 4014
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20088 3534 20116 3674
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 19260 2910 19472 2938
rect 18800 2746 19288 2774
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 18512 2372 18564 2378
rect 18512 2314 18564 2320
rect 18524 1970 18552 2314
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18512 1964 18564 1970
rect 18512 1906 18564 1912
rect 18616 800 18644 2246
rect 18892 800 18920 2586
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 19168 800 19196 2382
rect 19260 1698 19288 2746
rect 19248 1692 19300 1698
rect 19248 1634 19300 1640
rect 19444 800 19472 2910
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19708 2100 19760 2106
rect 19708 2042 19760 2048
rect 19720 800 19748 2042
rect 19996 800 20024 3402
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 20074 2680 20130 2689
rect 20074 2615 20130 2624
rect 20088 2446 20116 2615
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 20180 1578 20208 2994
rect 20260 2916 20312 2922
rect 20260 2858 20312 2864
rect 20272 2378 20300 2858
rect 20364 2774 20392 7262
rect 20456 6934 20484 8248
rect 20548 7818 20576 16351
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20732 15502 20760 15846
rect 20916 15722 20944 18838
rect 21100 18630 21128 24006
rect 21192 23186 21220 24142
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21192 21690 21220 23122
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 21284 21570 21312 24550
rect 21456 24268 21508 24274
rect 21456 24210 21508 24216
rect 21468 23526 21496 24210
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 21456 23520 21508 23526
rect 21456 23462 21508 23468
rect 21364 22636 21416 22642
rect 21468 22624 21496 23462
rect 21560 23050 21588 24142
rect 21548 23044 21600 23050
rect 21548 22986 21600 22992
rect 21416 22596 21496 22624
rect 21364 22578 21416 22584
rect 21192 21542 21312 21570
rect 21192 19242 21220 21542
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21284 19786 21312 21286
rect 21272 19780 21324 19786
rect 21272 19722 21324 19728
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21272 19236 21324 19242
rect 21272 19178 21324 19184
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21008 16454 21036 18226
rect 21086 17368 21142 17377
rect 21086 17303 21142 17312
rect 21100 17270 21128 17303
rect 21088 17264 21140 17270
rect 21088 17206 21140 17212
rect 21180 17264 21232 17270
rect 21180 17206 21232 17212
rect 21192 16998 21220 17206
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21192 16114 21220 16458
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 20916 15694 21036 15722
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 20640 11354 20668 13194
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20640 11150 20668 11181
rect 20628 11144 20680 11150
rect 20732 11098 20760 12786
rect 20824 12170 20852 15302
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20812 12164 20864 12170
rect 20812 12106 20864 12112
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20824 11354 20852 11698
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20916 11150 20944 12854
rect 21008 12434 21036 15694
rect 21192 15570 21220 16050
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21100 13326 21128 14758
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 21284 12434 21312 19178
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21376 16726 21404 19110
rect 21364 16720 21416 16726
rect 21364 16662 21416 16668
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21468 16017 21496 16050
rect 21454 16008 21510 16017
rect 21454 15943 21510 15952
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21468 15094 21496 15302
rect 21456 15088 21508 15094
rect 21456 15030 21508 15036
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21376 14521 21404 14758
rect 21362 14512 21418 14521
rect 21362 14447 21418 14456
rect 21468 13734 21496 14758
rect 21652 14532 21680 31726
rect 21928 30190 21956 31758
rect 21916 30184 21968 30190
rect 21916 30126 21968 30132
rect 22020 27674 22048 35634
rect 22112 35086 22140 56918
rect 22204 56846 22232 57394
rect 22192 56840 22244 56846
rect 22192 56782 22244 56788
rect 22204 51542 22232 56782
rect 22192 51536 22244 51542
rect 22192 51478 22244 51484
rect 22192 51400 22244 51406
rect 22192 51342 22244 51348
rect 22204 37874 22232 51342
rect 22296 48278 22324 60998
rect 22468 57928 22520 57934
rect 22468 57870 22520 57876
rect 22480 57458 22508 57870
rect 22468 57452 22520 57458
rect 22468 57394 22520 57400
rect 22480 51406 22508 57394
rect 22468 51400 22520 51406
rect 22468 51342 22520 51348
rect 22376 48544 22428 48550
rect 22376 48486 22428 48492
rect 22284 48272 22336 48278
rect 22284 48214 22336 48220
rect 22284 39636 22336 39642
rect 22284 39578 22336 39584
rect 22192 37868 22244 37874
rect 22192 37810 22244 37816
rect 22192 37188 22244 37194
rect 22192 37130 22244 37136
rect 22204 36854 22232 37130
rect 22192 36848 22244 36854
rect 22192 36790 22244 36796
rect 22296 35986 22324 39578
rect 22388 36174 22416 48486
rect 22836 42764 22888 42770
rect 22836 42706 22888 42712
rect 22744 42696 22796 42702
rect 22744 42638 22796 42644
rect 22652 42220 22704 42226
rect 22652 42162 22704 42168
rect 22664 41818 22692 42162
rect 22652 41812 22704 41818
rect 22652 41754 22704 41760
rect 22560 41064 22612 41070
rect 22560 41006 22612 41012
rect 22376 36168 22428 36174
rect 22376 36110 22428 36116
rect 22296 35958 22416 35986
rect 22192 35828 22244 35834
rect 22192 35770 22244 35776
rect 22204 35290 22232 35770
rect 22388 35290 22416 35958
rect 22192 35284 22244 35290
rect 22192 35226 22244 35232
rect 22376 35284 22428 35290
rect 22376 35226 22428 35232
rect 22468 35148 22520 35154
rect 22468 35090 22520 35096
rect 22100 35080 22152 35086
rect 22100 35022 22152 35028
rect 22480 34202 22508 35090
rect 22468 34196 22520 34202
rect 22468 34138 22520 34144
rect 22572 34082 22600 41006
rect 22652 40928 22704 40934
rect 22652 40870 22704 40876
rect 22664 40526 22692 40870
rect 22652 40520 22704 40526
rect 22652 40462 22704 40468
rect 22652 39840 22704 39846
rect 22652 39782 22704 39788
rect 22664 38962 22692 39782
rect 22756 39098 22784 42638
rect 22848 41614 22876 42706
rect 22940 41614 22968 60998
rect 23480 60852 23532 60858
rect 23480 60794 23532 60800
rect 23112 58676 23164 58682
rect 23112 58618 23164 58624
rect 23020 57928 23072 57934
rect 23020 57870 23072 57876
rect 23032 57254 23060 57870
rect 23124 57254 23152 58618
rect 23492 57934 23520 60794
rect 23204 57928 23256 57934
rect 23204 57870 23256 57876
rect 23480 57928 23532 57934
rect 23480 57870 23532 57876
rect 23216 57390 23244 57870
rect 23388 57792 23440 57798
rect 23388 57734 23440 57740
rect 23400 57526 23428 57734
rect 23388 57520 23440 57526
rect 23388 57462 23440 57468
rect 23204 57384 23256 57390
rect 23204 57326 23256 57332
rect 23020 57248 23072 57254
rect 23020 57190 23072 57196
rect 23112 57248 23164 57254
rect 23112 57190 23164 57196
rect 23124 55214 23152 57190
rect 23124 55186 23244 55214
rect 23020 51400 23072 51406
rect 23020 51342 23072 51348
rect 22836 41608 22888 41614
rect 22836 41550 22888 41556
rect 22928 41608 22980 41614
rect 22928 41550 22980 41556
rect 23032 40526 23060 51342
rect 23112 51264 23164 51270
rect 23112 51206 23164 51212
rect 23124 42226 23152 51206
rect 23216 45966 23244 55186
rect 23204 45960 23256 45966
rect 23204 45902 23256 45908
rect 23216 45626 23244 45902
rect 23296 45824 23348 45830
rect 23296 45766 23348 45772
rect 23204 45620 23256 45626
rect 23204 45562 23256 45568
rect 23112 42220 23164 42226
rect 23112 42162 23164 42168
rect 23020 40520 23072 40526
rect 23020 40462 23072 40468
rect 22836 40452 22888 40458
rect 22836 40394 22888 40400
rect 22744 39092 22796 39098
rect 22744 39034 22796 39040
rect 22848 38962 22876 40394
rect 23032 39506 23060 40462
rect 23020 39500 23072 39506
rect 23020 39442 23072 39448
rect 23032 38962 23060 39442
rect 23112 39432 23164 39438
rect 23112 39374 23164 39380
rect 22652 38956 22704 38962
rect 22652 38898 22704 38904
rect 22836 38956 22888 38962
rect 22836 38898 22888 38904
rect 23020 38956 23072 38962
rect 23020 38898 23072 38904
rect 22652 37868 22704 37874
rect 22652 37810 22704 37816
rect 22664 37754 22692 37810
rect 22664 37726 22784 37754
rect 22652 36576 22704 36582
rect 22652 36518 22704 36524
rect 22664 36174 22692 36518
rect 22652 36168 22704 36174
rect 22652 36110 22704 36116
rect 22756 35986 22784 37726
rect 22848 37126 22876 38898
rect 23020 37256 23072 37262
rect 23020 37198 23072 37204
rect 22836 37120 22888 37126
rect 22836 37062 22888 37068
rect 23032 36786 23060 37198
rect 23020 36780 23072 36786
rect 22204 34054 22600 34082
rect 22664 35958 22784 35986
rect 22940 36740 23020 36768
rect 22204 32434 22232 34054
rect 22192 32428 22244 32434
rect 22192 32370 22244 32376
rect 22560 32428 22612 32434
rect 22560 32370 22612 32376
rect 22192 31816 22244 31822
rect 22192 31758 22244 31764
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 22112 30598 22140 31214
rect 22204 30734 22232 31758
rect 22572 31754 22600 32370
rect 22664 31958 22692 35958
rect 22940 35329 22968 36740
rect 23020 36722 23072 36728
rect 22926 35320 22982 35329
rect 22926 35255 22982 35264
rect 22744 34944 22796 34950
rect 22744 34886 22796 34892
rect 22652 31952 22704 31958
rect 22652 31894 22704 31900
rect 22560 31748 22612 31754
rect 22560 31690 22612 31696
rect 22192 30728 22244 30734
rect 22192 30670 22244 30676
rect 22100 30592 22152 30598
rect 22100 30534 22152 30540
rect 22112 30138 22140 30534
rect 22204 30258 22232 30670
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22112 30110 22232 30138
rect 22008 27668 22060 27674
rect 22008 27610 22060 27616
rect 22204 26790 22232 30110
rect 22756 29209 22784 34886
rect 22940 33998 22968 35255
rect 23124 34626 23152 39374
rect 23204 37868 23256 37874
rect 23204 37810 23256 37816
rect 23216 37466 23244 37810
rect 23204 37460 23256 37466
rect 23204 37402 23256 37408
rect 23032 34598 23152 34626
rect 22928 33992 22980 33998
rect 22928 33934 22980 33940
rect 22836 33924 22888 33930
rect 22836 33866 22888 33872
rect 22848 29714 22876 33866
rect 23032 32298 23060 34598
rect 23112 34536 23164 34542
rect 23112 34478 23164 34484
rect 23020 32292 23072 32298
rect 23020 32234 23072 32240
rect 23032 31890 23060 32234
rect 23020 31884 23072 31890
rect 23020 31826 23072 31832
rect 23020 30728 23072 30734
rect 23020 30670 23072 30676
rect 23032 30190 23060 30670
rect 23020 30184 23072 30190
rect 23020 30126 23072 30132
rect 22836 29708 22888 29714
rect 22836 29650 22888 29656
rect 22742 29200 22798 29209
rect 22742 29135 22798 29144
rect 23032 28422 23060 30126
rect 23020 28416 23072 28422
rect 23020 28358 23072 28364
rect 22192 26784 22244 26790
rect 22192 26726 22244 26732
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21836 23730 21864 24006
rect 21824 23724 21876 23730
rect 21824 23666 21876 23672
rect 21732 23520 21784 23526
rect 21732 23462 21784 23468
rect 21744 20942 21772 23462
rect 21836 22642 21864 23666
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 22112 23474 22140 23598
rect 22020 23446 22140 23474
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 22020 21894 22048 23446
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 21732 20936 21784 20942
rect 21732 20878 21784 20884
rect 21824 19780 21876 19786
rect 21824 19722 21876 19728
rect 21732 16584 21784 16590
rect 21732 16526 21784 16532
rect 21744 15638 21772 16526
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21836 15473 21864 19722
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 22112 18358 22140 19246
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21928 17202 21956 17478
rect 21916 17196 21968 17202
rect 21916 17138 21968 17144
rect 21822 15464 21878 15473
rect 21822 15399 21878 15408
rect 21824 14544 21876 14550
rect 21652 14504 21824 14532
rect 21824 14486 21876 14492
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21362 13016 21418 13025
rect 21362 12951 21418 12960
rect 21008 12406 21128 12434
rect 20996 12368 21048 12374
rect 20994 12336 20996 12345
rect 21048 12336 21050 12345
rect 20994 12271 21050 12280
rect 20996 12164 21048 12170
rect 20996 12106 21048 12112
rect 20680 11092 20760 11098
rect 20628 11086 20760 11092
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20640 11070 20760 11086
rect 21008 11082 21036 12106
rect 20996 11076 21048 11082
rect 20640 10742 20668 11070
rect 20996 11018 21048 11024
rect 20628 10736 20680 10742
rect 20628 10678 20680 10684
rect 20640 10062 20668 10678
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20640 7342 20668 9454
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20824 9178 20852 9386
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20718 8256 20774 8265
rect 20718 8191 20774 8200
rect 20732 8090 20760 8191
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20916 7410 20944 7686
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 20548 7002 20576 7142
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20444 6928 20496 6934
rect 20444 6870 20496 6876
rect 20456 4146 20484 6870
rect 20640 4690 20668 7278
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20824 5234 20852 5510
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21008 4826 21036 5170
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20640 4486 20668 4626
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20444 3664 20496 3670
rect 20444 3606 20496 3612
rect 20456 2961 20484 3606
rect 20442 2952 20498 2961
rect 20442 2887 20498 2896
rect 20548 2836 20576 4218
rect 20640 4078 20668 4422
rect 21100 4146 21128 12406
rect 21192 12406 21312 12434
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20720 2848 20772 2854
rect 20548 2808 20720 2836
rect 20720 2790 20772 2796
rect 20364 2746 20668 2774
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 20640 1834 20668 2746
rect 20628 1828 20680 1834
rect 20628 1770 20680 1776
rect 20536 1760 20588 1766
rect 20536 1702 20588 1708
rect 20180 1550 20300 1578
rect 20272 800 20300 1550
rect 20548 800 20576 1702
rect 20824 800 20852 3334
rect 21192 3058 21220 12406
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21284 10674 21312 11290
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21284 10062 21312 10406
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21376 8514 21404 12951
rect 21468 11286 21496 13126
rect 21640 12776 21692 12782
rect 21640 12718 21692 12724
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21456 11280 21508 11286
rect 21456 11222 21508 11228
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21468 10810 21496 11086
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21456 10600 21508 10606
rect 21456 10542 21508 10548
rect 21284 8486 21404 8514
rect 21284 4622 21312 8486
rect 21468 8090 21496 10542
rect 21560 10538 21588 12650
rect 21652 10810 21680 12718
rect 21744 11898 21772 14350
rect 21836 13802 21864 14486
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21824 13388 21876 13394
rect 21824 13330 21876 13336
rect 21836 12442 21864 13330
rect 21824 12436 21876 12442
rect 21928 12434 21956 17138
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 22020 13938 22048 14894
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 22112 12918 22140 13466
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 21928 12406 22048 12434
rect 21824 12378 21876 12384
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 21640 10804 21692 10810
rect 21640 10746 21692 10752
rect 21640 10668 21692 10674
rect 21640 10610 21692 10616
rect 21548 10532 21600 10538
rect 21548 10474 21600 10480
rect 21546 10432 21602 10441
rect 21546 10367 21602 10376
rect 21560 10266 21588 10367
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21652 10062 21680 10610
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21744 9994 21772 11494
rect 21732 9988 21784 9994
rect 21732 9930 21784 9936
rect 21836 8430 21864 11562
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 21928 10198 21956 10746
rect 22020 10606 22048 12406
rect 22112 11762 22140 12854
rect 22204 12170 22232 26726
rect 22836 25152 22888 25158
rect 22836 25094 22888 25100
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22296 23866 22324 24006
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22296 22982 22324 23802
rect 22480 23322 22508 24754
rect 22560 24676 22612 24682
rect 22560 24618 22612 24624
rect 22572 24342 22600 24618
rect 22744 24608 22796 24614
rect 22744 24550 22796 24556
rect 22560 24336 22612 24342
rect 22560 24278 22612 24284
rect 22652 24336 22704 24342
rect 22652 24278 22704 24284
rect 22664 23662 22692 24278
rect 22756 23730 22784 24550
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 22652 23656 22704 23662
rect 22848 23610 22876 25094
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 23032 24070 23060 24142
rect 23020 24064 23072 24070
rect 23020 24006 23072 24012
rect 22652 23598 22704 23604
rect 22756 23582 22876 23610
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 22284 22976 22336 22982
rect 22284 22918 22336 22924
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 22388 22030 22416 22510
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22296 20058 22324 21966
rect 22388 21554 22416 21966
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22388 20466 22416 21490
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22388 19922 22416 20402
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22388 19310 22416 19858
rect 22664 19786 22692 20878
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 22480 18426 22508 19246
rect 22560 18896 22612 18902
rect 22560 18838 22612 18844
rect 22572 18630 22600 18838
rect 22560 18624 22612 18630
rect 22560 18566 22612 18572
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22480 17746 22508 18226
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22480 16046 22508 17682
rect 22664 17377 22692 19722
rect 22650 17368 22706 17377
rect 22650 17303 22706 17312
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22664 17105 22692 17138
rect 22650 17096 22706 17105
rect 22650 17031 22706 17040
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 22468 16040 22520 16046
rect 22468 15982 22520 15988
rect 22480 15570 22508 15982
rect 22572 15638 22600 16730
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22560 15632 22612 15638
rect 22560 15574 22612 15580
rect 22468 15564 22520 15570
rect 22468 15506 22520 15512
rect 22480 14958 22508 15506
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22296 13530 22324 13874
rect 22284 13524 22336 13530
rect 22284 13466 22336 13472
rect 22284 12980 22336 12986
rect 22284 12922 22336 12928
rect 22296 12866 22324 12922
rect 22480 12866 22508 14010
rect 22296 12838 22508 12866
rect 22664 12850 22692 16186
rect 22652 12844 22704 12850
rect 22192 12164 22244 12170
rect 22192 12106 22244 12112
rect 22388 12102 22416 12838
rect 22652 12786 22704 12792
rect 22560 12776 22612 12782
rect 22756 12764 22784 23582
rect 22928 22976 22980 22982
rect 22928 22918 22980 22924
rect 22940 22710 22968 22918
rect 22928 22704 22980 22710
rect 22928 22646 22980 22652
rect 23124 22094 23152 34478
rect 23308 31822 23336 45766
rect 23480 40384 23532 40390
rect 23480 40326 23532 40332
rect 23492 36786 23520 40326
rect 23848 38752 23900 38758
rect 23848 38694 23900 38700
rect 23388 36780 23440 36786
rect 23388 36722 23440 36728
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23400 34610 23428 36722
rect 23572 35488 23624 35494
rect 23572 35430 23624 35436
rect 23388 34604 23440 34610
rect 23388 34546 23440 34552
rect 23584 33522 23612 35430
rect 23860 34610 23888 38694
rect 23664 34604 23716 34610
rect 23664 34546 23716 34552
rect 23848 34604 23900 34610
rect 23848 34546 23900 34552
rect 23676 34474 23704 34546
rect 23664 34468 23716 34474
rect 23664 34410 23716 34416
rect 23572 33516 23624 33522
rect 23572 33458 23624 33464
rect 23584 32910 23612 33458
rect 23676 33454 23704 34410
rect 23952 33862 23980 60998
rect 24596 60790 24624 63294
rect 25134 63200 25190 64000
rect 25870 63322 25926 64000
rect 25870 63294 26096 63322
rect 25870 63200 25926 63294
rect 25148 61198 25176 63200
rect 26068 61198 26096 63294
rect 26606 63200 26662 64000
rect 27342 63322 27398 64000
rect 28078 63322 28134 64000
rect 28814 63322 28870 64000
rect 29550 63322 29606 64000
rect 27342 63294 27568 63322
rect 27342 63200 27398 63294
rect 25136 61192 25188 61198
rect 25136 61134 25188 61140
rect 26056 61192 26108 61198
rect 26056 61134 26108 61140
rect 25136 61056 25188 61062
rect 25136 60998 25188 61004
rect 24584 60784 24636 60790
rect 24584 60726 24636 60732
rect 24768 57860 24820 57866
rect 24768 57802 24820 57808
rect 24860 57860 24912 57866
rect 24860 57802 24912 57808
rect 24780 48618 24808 57802
rect 24872 56982 24900 57802
rect 24860 56976 24912 56982
rect 24860 56918 24912 56924
rect 24768 48612 24820 48618
rect 24768 48554 24820 48560
rect 25148 45554 25176 60998
rect 26620 60722 26648 63200
rect 27540 61198 27568 63294
rect 28078 63294 28396 63322
rect 28078 63200 28134 63294
rect 28368 61198 28396 63294
rect 28814 63294 28948 63322
rect 28814 63200 28870 63294
rect 27528 61192 27580 61198
rect 27528 61134 27580 61140
rect 28356 61192 28408 61198
rect 28920 61180 28948 63294
rect 29550 63294 29684 63322
rect 29550 63200 29606 63294
rect 29000 61192 29052 61198
rect 28920 61152 29000 61180
rect 28356 61134 28408 61140
rect 29000 61134 29052 61140
rect 27620 61056 27672 61062
rect 27620 60998 27672 61004
rect 28540 61056 28592 61062
rect 28540 60998 28592 61004
rect 26884 60852 26936 60858
rect 26884 60794 26936 60800
rect 26608 60716 26660 60722
rect 26608 60658 26660 60664
rect 25320 60580 25372 60586
rect 25320 60522 25372 60528
rect 25056 45526 25176 45554
rect 24124 45280 24176 45286
rect 24124 45222 24176 45228
rect 24136 37262 24164 45222
rect 24860 41608 24912 41614
rect 24860 41550 24912 41556
rect 24872 39370 24900 41550
rect 24860 39364 24912 39370
rect 24860 39306 24912 39312
rect 24952 38820 25004 38826
rect 24952 38762 25004 38768
rect 24124 37256 24176 37262
rect 24124 37198 24176 37204
rect 24964 36174 24992 38762
rect 24952 36168 25004 36174
rect 24766 36136 24822 36145
rect 24952 36110 25004 36116
rect 24766 36071 24768 36080
rect 24820 36071 24822 36080
rect 24768 36042 24820 36048
rect 24860 35692 24912 35698
rect 24860 35634 24912 35640
rect 24032 35624 24084 35630
rect 24032 35566 24084 35572
rect 24044 35086 24072 35566
rect 24308 35488 24360 35494
rect 24308 35430 24360 35436
rect 24032 35080 24084 35086
rect 24032 35022 24084 35028
rect 24122 35048 24178 35057
rect 24122 34983 24124 34992
rect 24176 34983 24178 34992
rect 24216 35012 24268 35018
rect 24124 34954 24176 34960
rect 24216 34954 24268 34960
rect 24228 34474 24256 34954
rect 24216 34468 24268 34474
rect 24216 34410 24268 34416
rect 23940 33856 23992 33862
rect 23940 33798 23992 33804
rect 23664 33448 23716 33454
rect 23664 33390 23716 33396
rect 23940 33448 23992 33454
rect 23940 33390 23992 33396
rect 23572 32904 23624 32910
rect 23492 32864 23572 32892
rect 23296 31816 23348 31822
rect 23296 31758 23348 31764
rect 23296 31136 23348 31142
rect 23296 31078 23348 31084
rect 23308 30734 23336 31078
rect 23296 30728 23348 30734
rect 23296 30670 23348 30676
rect 23492 30326 23520 32864
rect 23572 32846 23624 32852
rect 23572 31748 23624 31754
rect 23572 31690 23624 31696
rect 23584 30870 23612 31690
rect 23572 30864 23624 30870
rect 23572 30806 23624 30812
rect 23480 30320 23532 30326
rect 23480 30262 23532 30268
rect 23388 26036 23440 26042
rect 23388 25978 23440 25984
rect 23204 24744 23256 24750
rect 23204 24686 23256 24692
rect 23216 24070 23244 24686
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23296 24064 23348 24070
rect 23296 24006 23348 24012
rect 23216 23730 23244 24006
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 23308 22642 23336 24006
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 22848 22066 23152 22094
rect 22848 17649 22876 22066
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 22940 21622 22968 21830
rect 22928 21616 22980 21622
rect 22928 21558 22980 21564
rect 22928 20800 22980 20806
rect 22928 20742 22980 20748
rect 22940 20534 22968 20742
rect 22928 20528 22980 20534
rect 22928 20470 22980 20476
rect 23400 19174 23428 25978
rect 23572 24812 23624 24818
rect 23572 24754 23624 24760
rect 23584 22438 23612 24754
rect 23952 24750 23980 33390
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 24216 29164 24268 29170
rect 24216 29106 24268 29112
rect 24136 29073 24164 29106
rect 24122 29064 24178 29073
rect 24122 28999 24178 29008
rect 24032 27600 24084 27606
rect 24032 27542 24084 27548
rect 23940 24744 23992 24750
rect 23940 24686 23992 24692
rect 23848 23044 23900 23050
rect 23848 22986 23900 22992
rect 23860 22778 23888 22986
rect 23848 22772 23900 22778
rect 23848 22714 23900 22720
rect 23572 22432 23624 22438
rect 23572 22374 23624 22380
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 23664 18760 23716 18766
rect 23664 18702 23716 18708
rect 22928 18624 22980 18630
rect 22928 18566 22980 18572
rect 22940 18358 22968 18566
rect 22928 18352 22980 18358
rect 22928 18294 22980 18300
rect 23388 18148 23440 18154
rect 23388 18090 23440 18096
rect 23400 17678 23428 18090
rect 23676 18086 23704 18702
rect 23664 18080 23716 18086
rect 23664 18022 23716 18028
rect 23388 17672 23440 17678
rect 22834 17640 22890 17649
rect 23388 17614 23440 17620
rect 22834 17575 22890 17584
rect 22928 17604 22980 17610
rect 22560 12718 22612 12724
rect 22747 12736 22784 12764
rect 22468 12708 22520 12714
rect 22468 12650 22520 12656
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22296 11830 22324 12038
rect 22284 11824 22336 11830
rect 22284 11766 22336 11772
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22008 10600 22060 10606
rect 22008 10542 22060 10548
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 22006 10296 22062 10305
rect 22006 10231 22008 10240
rect 22060 10231 22062 10240
rect 22008 10202 22060 10208
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 22098 10160 22154 10169
rect 22098 10095 22154 10104
rect 22112 10062 22140 10095
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21364 7268 21416 7274
rect 21364 7210 21416 7216
rect 21376 6934 21404 7210
rect 22204 7041 22232 10542
rect 22190 7032 22246 7041
rect 22190 6967 22246 6976
rect 21364 6928 21416 6934
rect 21364 6870 21416 6876
rect 22098 6896 22154 6905
rect 22098 6831 22154 6840
rect 22112 6798 22140 6831
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 21638 6488 21694 6497
rect 21638 6423 21694 6432
rect 21652 6322 21680 6423
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 22006 6080 22062 6089
rect 22006 6015 22062 6024
rect 22020 5778 22048 6015
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 21364 5636 21416 5642
rect 21824 5636 21876 5642
rect 21364 5578 21416 5584
rect 21744 5596 21824 5624
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 21088 2984 21140 2990
rect 21088 2926 21140 2932
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 21008 2106 21036 2382
rect 20996 2100 21048 2106
rect 20996 2042 21048 2048
rect 21100 800 21128 2926
rect 21376 800 21404 5578
rect 21640 5160 21692 5166
rect 21640 5102 21692 5108
rect 21652 800 21680 5102
rect 21744 4554 21772 5596
rect 21824 5578 21876 5584
rect 22008 5160 22060 5166
rect 22008 5102 22060 5108
rect 21732 4548 21784 4554
rect 21732 4490 21784 4496
rect 21744 3602 21772 4490
rect 22020 4146 22048 5102
rect 22204 4690 22232 6967
rect 22296 5710 22324 10610
rect 22480 10130 22508 12650
rect 22572 11354 22600 12718
rect 22747 12696 22775 12736
rect 22747 12668 22784 12696
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22572 10588 22600 11086
rect 22652 10600 22704 10606
rect 22572 10560 22652 10588
rect 22652 10542 22704 10548
rect 22664 10266 22692 10542
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22468 10124 22520 10130
rect 22468 10066 22520 10072
rect 22376 6928 22428 6934
rect 22376 6870 22428 6876
rect 22388 6769 22416 6870
rect 22374 6760 22430 6769
rect 22374 6695 22430 6704
rect 22560 6724 22612 6730
rect 22612 6684 22692 6712
rect 22560 6666 22612 6672
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22388 5642 22416 6598
rect 22560 6180 22612 6186
rect 22560 6122 22612 6128
rect 22466 5808 22522 5817
rect 22466 5743 22468 5752
rect 22520 5743 22522 5752
rect 22468 5714 22520 5720
rect 22376 5636 22428 5642
rect 22376 5578 22428 5584
rect 22466 4856 22522 4865
rect 22466 4791 22522 4800
rect 22284 4752 22336 4758
rect 22284 4694 22336 4700
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 22296 4146 22324 4694
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22020 3777 22048 4082
rect 22006 3768 22062 3777
rect 22480 3738 22508 4791
rect 22006 3703 22062 3712
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 21732 3596 21784 3602
rect 21732 3538 21784 3544
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 22296 3097 22324 3130
rect 22282 3088 22338 3097
rect 22192 3052 22244 3058
rect 22282 3023 22338 3032
rect 22192 2994 22244 3000
rect 21916 1964 21968 1970
rect 21916 1906 21968 1912
rect 21928 800 21956 1906
rect 22204 800 22232 2994
rect 22572 2774 22600 6122
rect 22664 5710 22692 6684
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22756 5574 22784 12668
rect 22848 10674 22876 17575
rect 22928 17546 22980 17552
rect 22940 16794 22968 17546
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 23952 17270 23980 17478
rect 23940 17264 23992 17270
rect 23940 17206 23992 17212
rect 22928 16788 22980 16794
rect 22928 16730 22980 16736
rect 23202 16008 23258 16017
rect 23202 15943 23258 15952
rect 23216 15366 23244 15943
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23308 15366 23336 15642
rect 23204 15360 23256 15366
rect 23204 15302 23256 15308
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 23020 14612 23072 14618
rect 23020 14554 23072 14560
rect 23032 14498 23060 14554
rect 22940 14470 23060 14498
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22836 6860 22888 6866
rect 22836 6802 22888 6808
rect 22848 6633 22876 6802
rect 22834 6624 22890 6633
rect 22834 6559 22890 6568
rect 22940 6322 22968 14470
rect 23216 12782 23244 15302
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 23112 12640 23164 12646
rect 23112 12582 23164 12588
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23032 11694 23060 12038
rect 23124 11762 23152 12582
rect 23204 12164 23256 12170
rect 23204 12106 23256 12112
rect 23112 11756 23164 11762
rect 23112 11698 23164 11704
rect 23020 11688 23072 11694
rect 23020 11630 23072 11636
rect 23112 9444 23164 9450
rect 23112 9386 23164 9392
rect 23020 8424 23072 8430
rect 23020 8366 23072 8372
rect 23032 6798 23060 8366
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 22928 6316 22980 6322
rect 22928 6258 22980 6264
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22848 5914 22876 6190
rect 22836 5908 22888 5914
rect 22836 5850 22888 5856
rect 23020 5636 23072 5642
rect 23020 5578 23072 5584
rect 22744 5568 22796 5574
rect 22744 5510 22796 5516
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 22834 4720 22890 4729
rect 22940 4690 22968 4966
rect 23032 4826 23060 5578
rect 23124 5302 23152 9386
rect 23216 7342 23244 12106
rect 23308 11150 23336 15302
rect 23492 13938 23520 15846
rect 23572 15496 23624 15502
rect 23570 15464 23572 15473
rect 23624 15464 23626 15473
rect 23570 15399 23626 15408
rect 23848 15428 23900 15434
rect 23848 15370 23900 15376
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23676 11762 23704 13806
rect 23860 13530 23888 15370
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 23952 12918 23980 14350
rect 23940 12912 23992 12918
rect 23940 12854 23992 12860
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 23768 11898 23796 12786
rect 23952 12434 23980 12854
rect 23860 12406 23980 12434
rect 23756 11892 23808 11898
rect 23756 11834 23808 11840
rect 23860 11762 23888 12406
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23860 11354 23888 11698
rect 23848 11348 23900 11354
rect 23848 11290 23900 11296
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 23112 5296 23164 5302
rect 23112 5238 23164 5244
rect 23296 5160 23348 5166
rect 23296 5102 23348 5108
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 22834 4655 22890 4664
rect 22928 4684 22980 4690
rect 22848 4622 22876 4655
rect 22928 4626 22980 4632
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22940 4282 22968 4626
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 22744 2848 22796 2854
rect 22744 2790 22796 2796
rect 22480 2746 22600 2774
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 22388 2038 22416 2450
rect 22376 2032 22428 2038
rect 22376 1974 22428 1980
rect 22480 800 22508 2746
rect 22756 800 22784 2790
rect 23032 800 23060 3878
rect 23216 3126 23244 3878
rect 23204 3120 23256 3126
rect 23204 3062 23256 3068
rect 23308 800 23336 5102
rect 23400 2446 23428 11086
rect 23952 10674 23980 12038
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23664 10056 23716 10062
rect 23756 10056 23808 10062
rect 23664 9998 23716 10004
rect 23754 10024 23756 10033
rect 23808 10024 23810 10033
rect 23570 9752 23626 9761
rect 23676 9722 23704 9998
rect 23754 9959 23810 9968
rect 23570 9687 23572 9696
rect 23624 9687 23626 9696
rect 23664 9716 23716 9722
rect 23572 9658 23624 9664
rect 23664 9658 23716 9664
rect 23664 9036 23716 9042
rect 23664 8978 23716 8984
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23584 7002 23612 8910
rect 23676 7818 23704 8978
rect 23664 7812 23716 7818
rect 23664 7754 23716 7760
rect 23572 6996 23624 7002
rect 23572 6938 23624 6944
rect 23570 6896 23626 6905
rect 23570 6831 23626 6840
rect 23584 5846 23612 6831
rect 23676 6322 23704 7754
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23676 5846 23704 6258
rect 23572 5840 23624 5846
rect 23572 5782 23624 5788
rect 23664 5840 23716 5846
rect 23664 5782 23716 5788
rect 23676 5642 23704 5782
rect 23664 5636 23716 5642
rect 23664 5578 23716 5584
rect 23768 5216 23796 7482
rect 23860 6186 23888 10406
rect 24044 10248 24072 27542
rect 24228 24682 24256 29106
rect 24320 29034 24348 35430
rect 24872 35290 24900 35634
rect 24964 35306 24992 36110
rect 25056 35578 25084 45526
rect 25136 36304 25188 36310
rect 25136 36246 25188 36252
rect 25148 35698 25176 36246
rect 25332 35698 25360 60522
rect 25412 57792 25464 57798
rect 25412 57734 25464 57740
rect 25504 57792 25556 57798
rect 25504 57734 25556 57740
rect 25424 55214 25452 57734
rect 25516 57594 25544 57734
rect 25504 57588 25556 57594
rect 25504 57530 25556 57536
rect 25780 57384 25832 57390
rect 25608 57332 25780 57338
rect 25608 57326 25832 57332
rect 25608 57310 25820 57326
rect 25608 57254 25636 57310
rect 25596 57248 25648 57254
rect 25596 57190 25648 57196
rect 25424 55186 25544 55214
rect 25136 35692 25188 35698
rect 25136 35634 25188 35640
rect 25320 35692 25372 35698
rect 25320 35634 25372 35640
rect 25412 35624 25464 35630
rect 25056 35550 25176 35578
rect 25412 35566 25464 35572
rect 24860 35284 24912 35290
rect 24964 35278 25084 35306
rect 24860 35226 24912 35232
rect 24952 35216 25004 35222
rect 24952 35158 25004 35164
rect 24768 35148 24820 35154
rect 24768 35090 24820 35096
rect 24780 34950 24808 35090
rect 24860 35080 24912 35086
rect 24860 35022 24912 35028
rect 24768 34944 24820 34950
rect 24768 34886 24820 34892
rect 24872 34678 24900 35022
rect 24768 34672 24820 34678
rect 24768 34614 24820 34620
rect 24860 34672 24912 34678
rect 24860 34614 24912 34620
rect 24492 34536 24544 34542
rect 24492 34478 24544 34484
rect 24400 31884 24452 31890
rect 24400 31826 24452 31832
rect 24412 29306 24440 31826
rect 24400 29300 24452 29306
rect 24400 29242 24452 29248
rect 24308 29028 24360 29034
rect 24308 28970 24360 28976
rect 24216 24676 24268 24682
rect 24216 24618 24268 24624
rect 24308 24676 24360 24682
rect 24308 24618 24360 24624
rect 24216 23792 24268 23798
rect 24216 23734 24268 23740
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 24136 19378 24164 20198
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 24124 15904 24176 15910
rect 24124 15846 24176 15852
rect 24136 15094 24164 15846
rect 24124 15088 24176 15094
rect 24124 15030 24176 15036
rect 24124 12844 24176 12850
rect 24124 12786 24176 12792
rect 23952 10220 24072 10248
rect 23952 6934 23980 10220
rect 23940 6928 23992 6934
rect 23940 6870 23992 6876
rect 24032 6928 24084 6934
rect 24032 6870 24084 6876
rect 24044 6497 24072 6870
rect 24030 6488 24086 6497
rect 23940 6452 23992 6458
rect 24030 6423 24086 6432
rect 23940 6394 23992 6400
rect 23848 6180 23900 6186
rect 23848 6122 23900 6128
rect 23952 5574 23980 6394
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 24044 5710 24072 6054
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 23940 5568 23992 5574
rect 23940 5510 23992 5516
rect 23940 5228 23992 5234
rect 23768 5188 23940 5216
rect 23940 5170 23992 5176
rect 23952 4146 23980 5170
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 23952 3534 23980 4082
rect 23940 3528 23992 3534
rect 23940 3470 23992 3476
rect 23952 3126 23980 3470
rect 23940 3120 23992 3126
rect 23940 3062 23992 3068
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 23584 2774 23612 2994
rect 24136 2774 24164 12786
rect 24228 11150 24256 23734
rect 24320 23526 24348 24618
rect 24308 23520 24360 23526
rect 24308 23462 24360 23468
rect 24320 22642 24348 23462
rect 24308 22636 24360 22642
rect 24308 22578 24360 22584
rect 24400 22092 24452 22098
rect 24400 22034 24452 22040
rect 24308 21548 24360 21554
rect 24308 21490 24360 21496
rect 24320 21078 24348 21490
rect 24412 21486 24440 22034
rect 24400 21480 24452 21486
rect 24400 21422 24452 21428
rect 24308 21072 24360 21078
rect 24308 21014 24360 21020
rect 24308 19372 24360 19378
rect 24308 19314 24360 19320
rect 24320 17338 24348 19314
rect 24308 17332 24360 17338
rect 24308 17274 24360 17280
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 24412 16658 24440 17274
rect 24504 16658 24532 34478
rect 24780 34066 24808 34614
rect 24964 34610 24992 35158
rect 24952 34604 25004 34610
rect 24952 34546 25004 34552
rect 25056 34134 25084 35278
rect 25044 34128 25096 34134
rect 25044 34070 25096 34076
rect 24768 34060 24820 34066
rect 24768 34002 24820 34008
rect 24676 33992 24728 33998
rect 24676 33934 24728 33940
rect 24860 33992 24912 33998
rect 25056 33980 25084 34070
rect 24912 33952 25084 33980
rect 24860 33934 24912 33940
rect 24584 31476 24636 31482
rect 24584 31418 24636 31424
rect 24596 31278 24624 31418
rect 24584 31272 24636 31278
rect 24584 31214 24636 31220
rect 24584 31136 24636 31142
rect 24584 31078 24636 31084
rect 24596 30734 24624 31078
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24688 26994 24716 33934
rect 24768 32224 24820 32230
rect 24768 32166 24820 32172
rect 24780 30734 24808 32166
rect 25148 31414 25176 35550
rect 25226 35320 25282 35329
rect 25282 35264 25360 35272
rect 25226 35255 25228 35264
rect 25280 35244 25360 35264
rect 25228 35226 25280 35232
rect 25228 33856 25280 33862
rect 25228 33798 25280 33804
rect 25240 32502 25268 33798
rect 25332 33590 25360 35244
rect 25424 34474 25452 35566
rect 25516 35154 25544 55186
rect 26896 39030 26924 60794
rect 27344 60512 27396 60518
rect 27344 60454 27396 60460
rect 27356 55214 27384 60454
rect 27356 55186 27476 55214
rect 26884 39024 26936 39030
rect 26884 38966 26936 38972
rect 26148 38888 26200 38894
rect 26148 38830 26200 38836
rect 26160 37942 26188 38830
rect 26148 37936 26200 37942
rect 26148 37878 26200 37884
rect 26516 37800 26568 37806
rect 26516 37742 26568 37748
rect 25596 37256 25648 37262
rect 25596 37198 25648 37204
rect 25504 35148 25556 35154
rect 25504 35090 25556 35096
rect 25502 35048 25558 35057
rect 25502 34983 25504 34992
rect 25556 34983 25558 34992
rect 25504 34954 25556 34960
rect 25412 34468 25464 34474
rect 25412 34410 25464 34416
rect 25424 33998 25452 34410
rect 25412 33992 25464 33998
rect 25412 33934 25464 33940
rect 25320 33584 25372 33590
rect 25320 33526 25372 33532
rect 25228 32496 25280 32502
rect 25228 32438 25280 32444
rect 25136 31408 25188 31414
rect 25136 31350 25188 31356
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 24768 30728 24820 30734
rect 24768 30670 24820 30676
rect 24860 30592 24912 30598
rect 24860 30534 24912 30540
rect 24676 26988 24728 26994
rect 24676 26930 24728 26936
rect 24872 26042 24900 30534
rect 24964 28490 24992 31282
rect 25332 29170 25360 33526
rect 25412 33516 25464 33522
rect 25412 33458 25464 33464
rect 25320 29164 25372 29170
rect 25320 29106 25372 29112
rect 25424 28558 25452 33458
rect 25608 32910 25636 37198
rect 26424 36032 26476 36038
rect 26424 35974 26476 35980
rect 25688 34536 25740 34542
rect 25688 34478 25740 34484
rect 25700 33318 25728 34478
rect 25780 34128 25832 34134
rect 25780 34070 25832 34076
rect 25792 33522 25820 34070
rect 26056 33992 26108 33998
rect 26056 33934 26108 33940
rect 25780 33516 25832 33522
rect 25780 33458 25832 33464
rect 25688 33312 25740 33318
rect 25688 33254 25740 33260
rect 25504 32904 25556 32910
rect 25504 32846 25556 32852
rect 25596 32904 25648 32910
rect 25596 32846 25648 32852
rect 25792 32892 25820 33458
rect 25964 32904 26016 32910
rect 25792 32864 25964 32892
rect 25516 32774 25544 32846
rect 25504 32768 25556 32774
rect 25504 32710 25556 32716
rect 25792 31754 25820 32864
rect 25964 32846 26016 32852
rect 25964 32292 26016 32298
rect 25964 32234 26016 32240
rect 25872 31952 25924 31958
rect 25872 31894 25924 31900
rect 25780 31748 25832 31754
rect 25780 31690 25832 31696
rect 25792 31278 25820 31690
rect 25884 31414 25912 31894
rect 25976 31890 26004 32234
rect 25964 31884 26016 31890
rect 25964 31826 26016 31832
rect 26068 31754 26096 33934
rect 26148 32904 26200 32910
rect 26148 32846 26200 32852
rect 25964 31748 26096 31754
rect 26016 31726 26096 31748
rect 25964 31690 26016 31696
rect 25872 31408 25924 31414
rect 25872 31350 25924 31356
rect 25976 31278 26004 31690
rect 26056 31680 26108 31686
rect 26056 31622 26108 31628
rect 26068 31346 26096 31622
rect 26056 31340 26108 31346
rect 26056 31282 26108 31288
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 25964 31272 26016 31278
rect 25964 31214 26016 31220
rect 26160 28762 26188 32846
rect 26332 31272 26384 31278
rect 26332 31214 26384 31220
rect 26148 28756 26200 28762
rect 26148 28698 26200 28704
rect 25412 28552 25464 28558
rect 25412 28494 25464 28500
rect 24952 28484 25004 28490
rect 24952 28426 25004 28432
rect 25320 27328 25372 27334
rect 25320 27270 25372 27276
rect 24860 26036 24912 26042
rect 24860 25978 24912 25984
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24584 23112 24636 23118
rect 24584 23054 24636 23060
rect 24596 22778 24624 23054
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24688 19854 24716 24550
rect 24964 24410 24992 25230
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 25228 24064 25280 24070
rect 25228 24006 25280 24012
rect 25044 23656 25096 23662
rect 25044 23598 25096 23604
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24780 23186 24808 23258
rect 25056 23254 25084 23598
rect 25044 23248 25096 23254
rect 25044 23190 25096 23196
rect 24768 23180 24820 23186
rect 24768 23122 24820 23128
rect 24780 19854 24808 23122
rect 25148 22030 25176 24006
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24872 20602 24900 20878
rect 24860 20596 24912 20602
rect 24860 20538 24912 20544
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 25136 18964 25188 18970
rect 25136 18906 25188 18912
rect 24582 18456 24638 18465
rect 24582 18391 24638 18400
rect 24596 16794 24624 18391
rect 25148 18358 25176 18906
rect 25136 18352 25188 18358
rect 25136 18294 25188 18300
rect 25044 18216 25096 18222
rect 25044 18158 25096 18164
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24872 16794 24900 17614
rect 25056 17542 25084 18158
rect 25044 17536 25096 17542
rect 25044 17478 25096 17484
rect 24584 16788 24636 16794
rect 24584 16730 24636 16736
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24492 16652 24544 16658
rect 24492 16594 24544 16600
rect 24504 12434 24532 16594
rect 25056 16572 25084 17478
rect 25136 16584 25188 16590
rect 25056 16544 25136 16572
rect 24860 16176 24912 16182
rect 24860 16118 24912 16124
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24320 12406 24532 12434
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24216 10056 24268 10062
rect 24216 9998 24268 10004
rect 24228 8430 24256 9998
rect 24216 8424 24268 8430
rect 24216 8366 24268 8372
rect 24228 5273 24256 8366
rect 24214 5264 24270 5273
rect 24214 5199 24270 5208
rect 24320 2774 24348 12406
rect 24490 11520 24546 11529
rect 24490 11455 24546 11464
rect 24504 9674 24532 11455
rect 24596 11354 24624 16050
rect 24768 14952 24820 14958
rect 24768 14894 24820 14900
rect 24676 14816 24728 14822
rect 24676 14758 24728 14764
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 24688 11150 24716 14758
rect 24780 14414 24808 14894
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24780 13394 24808 14350
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 24872 12782 24900 16118
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24964 14890 24992 16050
rect 24952 14884 25004 14890
rect 24952 14826 25004 14832
rect 25056 13258 25084 16544
rect 25136 16526 25188 16532
rect 25136 14272 25188 14278
rect 25136 14214 25188 14220
rect 25148 13326 25176 14214
rect 25136 13320 25188 13326
rect 25136 13262 25188 13268
rect 25044 13252 25096 13258
rect 25044 13194 25096 13200
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24584 10736 24636 10742
rect 24584 10678 24636 10684
rect 24412 9646 24532 9674
rect 24412 5642 24440 9646
rect 24596 9042 24624 10678
rect 25056 10470 25084 12038
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 24584 9036 24636 9042
rect 24636 8996 24716 9024
rect 24584 8978 24636 8984
rect 24688 7886 24716 8996
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24688 7546 24716 7822
rect 24780 7546 24808 8434
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24582 6896 24638 6905
rect 24582 6831 24584 6840
rect 24636 6831 24638 6840
rect 24584 6802 24636 6808
rect 24676 6724 24728 6730
rect 24676 6666 24728 6672
rect 24584 6656 24636 6662
rect 24584 6598 24636 6604
rect 24596 6118 24624 6598
rect 24492 6112 24544 6118
rect 24492 6054 24544 6060
rect 24584 6112 24636 6118
rect 24584 6054 24636 6060
rect 24400 5636 24452 5642
rect 24400 5578 24452 5584
rect 24504 5234 24532 6054
rect 24688 5778 24716 6666
rect 24872 6644 24900 7686
rect 24952 6656 25004 6662
rect 24780 6616 24952 6644
rect 24780 6458 24808 6616
rect 24952 6598 25004 6604
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 24780 6322 24900 6338
rect 24780 6316 24912 6322
rect 24780 6310 24860 6316
rect 24676 5772 24728 5778
rect 24676 5714 24728 5720
rect 24582 5672 24638 5681
rect 24582 5607 24584 5616
rect 24636 5607 24638 5616
rect 24584 5578 24636 5584
rect 24492 5228 24544 5234
rect 24492 5170 24544 5176
rect 24780 5030 24808 6310
rect 24860 6258 24912 6264
rect 24768 5024 24820 5030
rect 24768 4966 24820 4972
rect 24768 4752 24820 4758
rect 24766 4720 24768 4729
rect 24820 4720 24822 4729
rect 24766 4655 24822 4664
rect 24964 4622 24992 6394
rect 25056 6390 25084 10406
rect 25136 6792 25188 6798
rect 25134 6760 25136 6769
rect 25188 6760 25190 6769
rect 25134 6695 25190 6704
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25044 6384 25096 6390
rect 25044 6326 25096 6332
rect 25148 6089 25176 6598
rect 25134 6080 25190 6089
rect 25134 6015 25190 6024
rect 25240 5710 25268 24006
rect 25332 23118 25360 27270
rect 25872 26444 25924 26450
rect 25872 26386 25924 26392
rect 25688 26240 25740 26246
rect 25688 26182 25740 26188
rect 25596 25696 25648 25702
rect 25596 25638 25648 25644
rect 25608 24206 25636 25638
rect 25700 25226 25728 26182
rect 25884 25974 25912 26386
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 25872 25968 25924 25974
rect 25872 25910 25924 25916
rect 25884 25838 25912 25910
rect 25872 25832 25924 25838
rect 25872 25774 25924 25780
rect 26056 25832 26108 25838
rect 26056 25774 26108 25780
rect 25688 25220 25740 25226
rect 25688 25162 25740 25168
rect 25596 24200 25648 24206
rect 25596 24142 25648 24148
rect 25320 23112 25372 23118
rect 25320 23054 25372 23060
rect 25688 23112 25740 23118
rect 25688 23054 25740 23060
rect 25596 22976 25648 22982
rect 25596 22918 25648 22924
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25332 19854 25360 20742
rect 25320 19848 25372 19854
rect 25320 19790 25372 19796
rect 25504 19780 25556 19786
rect 25504 19722 25556 19728
rect 25516 19514 25544 19722
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 25320 18624 25372 18630
rect 25320 18566 25372 18572
rect 25412 18624 25464 18630
rect 25412 18566 25464 18572
rect 25332 17746 25360 18566
rect 25320 17740 25372 17746
rect 25320 17682 25372 17688
rect 25320 17536 25372 17542
rect 25320 17478 25372 17484
rect 25332 15706 25360 17478
rect 25424 17134 25452 18566
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25516 17270 25544 17614
rect 25504 17264 25556 17270
rect 25504 17206 25556 17212
rect 25412 17128 25464 17134
rect 25412 17070 25464 17076
rect 25502 17096 25558 17105
rect 25502 17031 25504 17040
rect 25556 17031 25558 17040
rect 25504 17002 25556 17008
rect 25412 16584 25464 16590
rect 25412 16526 25464 16532
rect 25424 16454 25452 16526
rect 25412 16448 25464 16454
rect 25410 16416 25412 16425
rect 25464 16416 25466 16425
rect 25410 16351 25466 16360
rect 25320 15700 25372 15706
rect 25320 15642 25372 15648
rect 25410 14512 25466 14521
rect 25410 14447 25466 14456
rect 25318 14376 25374 14385
rect 25424 14346 25452 14447
rect 25318 14311 25374 14320
rect 25412 14340 25464 14346
rect 25332 6458 25360 14311
rect 25412 14282 25464 14288
rect 25608 12434 25636 22918
rect 25700 18970 25728 23054
rect 25884 22094 25912 25774
rect 26068 24698 26096 25774
rect 26160 25158 26188 26250
rect 26240 25220 26292 25226
rect 26240 25162 26292 25168
rect 26148 25152 26200 25158
rect 26148 25094 26200 25100
rect 25976 24670 26096 24698
rect 25976 24070 26004 24670
rect 26056 24608 26108 24614
rect 26056 24550 26108 24556
rect 25964 24064 26016 24070
rect 25964 24006 26016 24012
rect 26068 23118 26096 24550
rect 26252 23322 26280 25162
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 26148 23180 26200 23186
rect 26200 23140 26280 23168
rect 26148 23122 26200 23128
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 26252 22778 26280 23140
rect 26240 22772 26292 22778
rect 26240 22714 26292 22720
rect 25884 22066 26004 22094
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25870 18864 25926 18873
rect 25870 18799 25926 18808
rect 25780 18284 25832 18290
rect 25780 18226 25832 18232
rect 25792 17814 25820 18226
rect 25780 17808 25832 17814
rect 25780 17750 25832 17756
rect 25884 17660 25912 18799
rect 25792 17632 25912 17660
rect 25688 17264 25740 17270
rect 25688 17206 25740 17212
rect 25700 16998 25728 17206
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 25700 16726 25728 16934
rect 25688 16720 25740 16726
rect 25688 16662 25740 16668
rect 25688 15428 25740 15434
rect 25688 15370 25740 15376
rect 25700 13394 25728 15370
rect 25688 13388 25740 13394
rect 25688 13330 25740 13336
rect 25792 13274 25820 17632
rect 25976 15910 26004 22066
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 26160 20942 26188 21422
rect 26148 20936 26200 20942
rect 26148 20878 26200 20884
rect 26238 18320 26294 18329
rect 26344 18290 26372 31214
rect 26436 29102 26464 35974
rect 26528 30161 26556 37742
rect 26884 36916 26936 36922
rect 26884 36858 26936 36864
rect 26896 36650 26924 36858
rect 26884 36644 26936 36650
rect 26884 36586 26936 36592
rect 27344 36372 27396 36378
rect 27344 36314 27396 36320
rect 26884 35556 26936 35562
rect 26884 35498 26936 35504
rect 26896 34542 26924 35498
rect 26884 34536 26936 34542
rect 26884 34478 26936 34484
rect 27356 33522 27384 36314
rect 27344 33516 27396 33522
rect 27344 33458 27396 33464
rect 26608 33448 26660 33454
rect 26608 33390 26660 33396
rect 26514 30152 26570 30161
rect 26514 30087 26570 30096
rect 26424 29096 26476 29102
rect 26424 29038 26476 29044
rect 26620 26926 26648 33390
rect 27356 32910 27384 33458
rect 27344 32904 27396 32910
rect 27344 32846 27396 32852
rect 27344 32496 27396 32502
rect 27344 32438 27396 32444
rect 27160 32292 27212 32298
rect 27160 32234 27212 32240
rect 27172 28694 27200 32234
rect 27160 28688 27212 28694
rect 27160 28630 27212 28636
rect 26608 26920 26660 26926
rect 26608 26862 26660 26868
rect 26792 26308 26844 26314
rect 26792 26250 26844 26256
rect 26424 24812 26476 24818
rect 26424 24754 26476 24760
rect 26436 24410 26464 24754
rect 26424 24404 26476 24410
rect 26424 24346 26476 24352
rect 26436 22778 26464 24346
rect 26698 22944 26754 22953
rect 26698 22879 26754 22888
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 26516 21956 26568 21962
rect 26516 21898 26568 21904
rect 26528 20058 26556 21898
rect 26712 21350 26740 22879
rect 26700 21344 26752 21350
rect 26700 21286 26752 21292
rect 26700 20800 26752 20806
rect 26700 20742 26752 20748
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26606 18320 26662 18329
rect 26238 18255 26294 18264
rect 26332 18284 26384 18290
rect 26148 17808 26200 17814
rect 26148 17750 26200 17756
rect 26160 17270 26188 17750
rect 26148 17264 26200 17270
rect 26148 17206 26200 17212
rect 26252 17202 26280 18255
rect 26606 18255 26662 18264
rect 26332 18226 26384 18232
rect 26330 18184 26386 18193
rect 26330 18119 26386 18128
rect 26344 18086 26372 18119
rect 26332 18080 26384 18086
rect 26332 18022 26384 18028
rect 26424 18080 26476 18086
rect 26424 18022 26476 18028
rect 26436 17202 26464 18022
rect 26240 17196 26292 17202
rect 26240 17138 26292 17144
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26148 16788 26200 16794
rect 26148 16730 26200 16736
rect 26160 15978 26188 16730
rect 26332 16652 26384 16658
rect 26332 16594 26384 16600
rect 26240 16584 26292 16590
rect 26240 16526 26292 16532
rect 26148 15972 26200 15978
rect 26148 15914 26200 15920
rect 25964 15904 26016 15910
rect 25964 15846 26016 15852
rect 25424 12406 25636 12434
rect 25700 13246 25820 13274
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25228 5704 25280 5710
rect 25228 5646 25280 5652
rect 25136 5636 25188 5642
rect 25136 5578 25188 5584
rect 25044 5092 25096 5098
rect 25044 5034 25096 5040
rect 25056 4690 25084 5034
rect 25148 4865 25176 5578
rect 25134 4856 25190 4865
rect 25134 4791 25190 4800
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 24952 4616 25004 4622
rect 24952 4558 25004 4564
rect 24584 4480 24636 4486
rect 24584 4422 24636 4428
rect 24596 4214 24624 4422
rect 25056 4282 25084 4626
rect 25136 4548 25188 4554
rect 25136 4490 25188 4496
rect 25044 4276 25096 4282
rect 25044 4218 25096 4224
rect 24584 4208 24636 4214
rect 24584 4150 24636 4156
rect 24952 4004 25004 4010
rect 24952 3946 25004 3952
rect 24964 3913 24992 3946
rect 24950 3904 25006 3913
rect 24950 3839 25006 3848
rect 24584 3664 24636 3670
rect 24584 3606 24636 3612
rect 24596 3058 24624 3606
rect 25148 3602 25176 4490
rect 25424 3942 25452 12406
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 25516 11898 25544 12174
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25596 11620 25648 11626
rect 25596 11562 25648 11568
rect 25504 11348 25556 11354
rect 25504 11290 25556 11296
rect 25516 10033 25544 11290
rect 25608 11150 25636 11562
rect 25596 11144 25648 11150
rect 25596 11086 25648 11092
rect 25502 10024 25558 10033
rect 25502 9959 25558 9968
rect 25516 9674 25544 9959
rect 25516 9646 25636 9674
rect 25504 8356 25556 8362
rect 25504 8298 25556 8304
rect 25516 7410 25544 8298
rect 25504 7404 25556 7410
rect 25504 7346 25556 7352
rect 25516 6322 25544 7346
rect 25608 6882 25636 9646
rect 25700 9586 25728 13246
rect 25872 12980 25924 12986
rect 25872 12922 25924 12928
rect 25884 11014 25912 12922
rect 26160 12850 26188 15914
rect 26252 12986 26280 16526
rect 26344 15688 26372 16594
rect 26344 15660 26556 15688
rect 26424 15564 26476 15570
rect 26424 15506 26476 15512
rect 26332 15020 26384 15026
rect 26332 14962 26384 14968
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26344 12714 26372 14962
rect 26436 14414 26464 15506
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 26528 12850 26556 15660
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 26332 12708 26384 12714
rect 26332 12650 26384 12656
rect 26620 12434 26648 18255
rect 26528 12406 26648 12434
rect 26056 12232 26108 12238
rect 26056 12174 26108 12180
rect 26068 11898 26096 12174
rect 26056 11892 26108 11898
rect 26056 11834 26108 11840
rect 26424 11212 26476 11218
rect 26424 11154 26476 11160
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 25792 10266 25820 10950
rect 25780 10260 25832 10266
rect 25780 10202 25832 10208
rect 25872 10056 25924 10062
rect 25872 9998 25924 10004
rect 25780 9716 25832 9722
rect 25780 9658 25832 9664
rect 25688 9580 25740 9586
rect 25688 9522 25740 9528
rect 25792 8072 25820 9658
rect 25884 9654 25912 9998
rect 26436 9926 26464 11154
rect 26424 9920 26476 9926
rect 26424 9862 26476 9868
rect 25872 9648 25924 9654
rect 25872 9590 25924 9596
rect 25872 8900 25924 8906
rect 25872 8842 25924 8848
rect 25884 8634 25912 8842
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 25976 8566 26004 8774
rect 26528 8634 26556 12406
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26620 9994 26648 10406
rect 26608 9988 26660 9994
rect 26608 9930 26660 9936
rect 26712 9450 26740 20742
rect 26804 14793 26832 26250
rect 26884 26240 26936 26246
rect 26884 26182 26936 26188
rect 26896 25498 26924 26182
rect 26884 25492 26936 25498
rect 26884 25434 26936 25440
rect 27252 24812 27304 24818
rect 27252 24754 27304 24760
rect 27160 24336 27212 24342
rect 27160 24278 27212 24284
rect 27068 24268 27120 24274
rect 27068 24210 27120 24216
rect 27080 23866 27108 24210
rect 27068 23860 27120 23866
rect 27068 23802 27120 23808
rect 27172 23798 27200 24278
rect 27264 23866 27292 24754
rect 27252 23860 27304 23866
rect 27252 23802 27304 23808
rect 27160 23792 27212 23798
rect 27160 23734 27212 23740
rect 27158 23216 27214 23225
rect 27158 23151 27214 23160
rect 26884 22976 26936 22982
rect 26884 22918 26936 22924
rect 26896 22030 26924 22918
rect 27068 22772 27120 22778
rect 27068 22714 27120 22720
rect 26976 22160 27028 22166
rect 26976 22102 27028 22108
rect 26884 22024 26936 22030
rect 26884 21966 26936 21972
rect 26988 20534 27016 22102
rect 26976 20528 27028 20534
rect 26976 20470 27028 20476
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 27080 18272 27108 22714
rect 27172 21690 27200 23151
rect 27252 22500 27304 22506
rect 27252 22442 27304 22448
rect 27264 21894 27292 22442
rect 27252 21888 27304 21894
rect 27252 21830 27304 21836
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 27356 21554 27384 32438
rect 27448 30598 27476 55186
rect 27528 42152 27580 42158
rect 27528 42094 27580 42100
rect 27540 38729 27568 42094
rect 27632 40934 27660 60998
rect 28264 60308 28316 60314
rect 28264 60250 28316 60256
rect 27620 40928 27672 40934
rect 27620 40870 27672 40876
rect 28276 40458 28304 60250
rect 28356 56160 28408 56166
rect 28356 56102 28408 56108
rect 28368 46034 28396 56102
rect 28356 46028 28408 46034
rect 28356 45970 28408 45976
rect 28264 40452 28316 40458
rect 28264 40394 28316 40400
rect 27526 38720 27582 38729
rect 27526 38655 27582 38664
rect 27620 34740 27672 34746
rect 27620 34682 27672 34688
rect 27632 33522 27660 34682
rect 27528 33516 27580 33522
rect 27528 33458 27580 33464
rect 27620 33516 27672 33522
rect 27620 33458 27672 33464
rect 28448 33516 28500 33522
rect 28448 33458 28500 33464
rect 27540 33046 27568 33458
rect 27528 33040 27580 33046
rect 27528 32982 27580 32988
rect 27528 32904 27580 32910
rect 27528 32846 27580 32852
rect 27540 32298 27568 32846
rect 27632 32842 27660 33458
rect 27620 32836 27672 32842
rect 27620 32778 27672 32784
rect 27528 32292 27580 32298
rect 27528 32234 27580 32240
rect 27436 30592 27488 30598
rect 27436 30534 27488 30540
rect 27712 29028 27764 29034
rect 27712 28970 27764 28976
rect 27436 26308 27488 26314
rect 27436 26250 27488 26256
rect 27448 22642 27476 26250
rect 27528 25220 27580 25226
rect 27528 25162 27580 25168
rect 27540 24834 27568 25162
rect 27540 24806 27660 24834
rect 27632 24750 27660 24806
rect 27620 24744 27672 24750
rect 27620 24686 27672 24692
rect 27620 24608 27672 24614
rect 27620 24550 27672 24556
rect 27528 24200 27580 24206
rect 27528 24142 27580 24148
rect 27540 23866 27568 24142
rect 27528 23860 27580 23866
rect 27528 23802 27580 23808
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 27448 21690 27476 22578
rect 27632 22522 27660 24550
rect 27724 22642 27752 28970
rect 28356 26444 28408 26450
rect 28356 26386 28408 26392
rect 27988 25900 28040 25906
rect 27988 25842 28040 25848
rect 27804 25696 27856 25702
rect 27804 25638 27856 25644
rect 27816 25498 27844 25638
rect 27804 25492 27856 25498
rect 27804 25434 27856 25440
rect 28000 24070 28028 25842
rect 27988 24064 28040 24070
rect 27988 24006 28040 24012
rect 28000 23730 28028 24006
rect 27896 23724 27948 23730
rect 27896 23666 27948 23672
rect 27988 23724 28040 23730
rect 27988 23666 28040 23672
rect 27908 23254 27936 23666
rect 27896 23248 27948 23254
rect 27896 23190 27948 23196
rect 28000 22642 28028 23666
rect 28264 23588 28316 23594
rect 28264 23530 28316 23536
rect 27712 22636 27764 22642
rect 27988 22636 28040 22642
rect 27764 22596 27844 22624
rect 27712 22578 27764 22584
rect 27632 22494 27752 22522
rect 27526 22128 27582 22137
rect 27724 22094 27752 22494
rect 27816 22137 27844 22596
rect 27988 22578 28040 22584
rect 28000 22166 28028 22578
rect 28276 22522 28304 23530
rect 28368 22642 28396 26386
rect 28460 25974 28488 33458
rect 28552 30734 28580 60998
rect 29656 60722 29684 63294
rect 30286 63200 30342 64000
rect 31022 63200 31078 64000
rect 31758 63200 31814 64000
rect 32494 63200 32550 64000
rect 33230 63200 33286 64000
rect 33966 63200 34022 64000
rect 34702 63200 34758 64000
rect 35438 63322 35494 64000
rect 36174 63322 36230 64000
rect 36910 63322 36966 64000
rect 35438 63294 35848 63322
rect 35438 63200 35494 63294
rect 30012 61056 30064 61062
rect 30012 60998 30064 61004
rect 29644 60716 29696 60722
rect 29644 60658 29696 60664
rect 29828 60512 29880 60518
rect 29828 60454 29880 60460
rect 29552 56500 29604 56506
rect 29552 56442 29604 56448
rect 29460 56364 29512 56370
rect 29460 56306 29512 56312
rect 29472 55962 29500 56306
rect 29564 56234 29592 56442
rect 29644 56364 29696 56370
rect 29644 56306 29696 56312
rect 29552 56228 29604 56234
rect 29552 56170 29604 56176
rect 29656 56166 29684 56306
rect 29644 56160 29696 56166
rect 29644 56102 29696 56108
rect 29656 55962 29684 56102
rect 29460 55956 29512 55962
rect 29460 55898 29512 55904
rect 29644 55956 29696 55962
rect 29644 55898 29696 55904
rect 29644 39296 29696 39302
rect 29644 39238 29696 39244
rect 29552 33312 29604 33318
rect 29552 33254 29604 33260
rect 28540 30728 28592 30734
rect 28540 30670 28592 30676
rect 28448 25968 28500 25974
rect 28448 25910 28500 25916
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 28184 22494 28304 22522
rect 27988 22160 28040 22166
rect 27526 22063 27582 22072
rect 27632 22066 27752 22094
rect 27802 22128 27858 22137
rect 27988 22102 28040 22108
rect 27540 22001 27568 22063
rect 27526 21992 27582 22001
rect 27526 21927 27582 21936
rect 27436 21684 27488 21690
rect 27436 21626 27488 21632
rect 27632 21554 27660 22066
rect 27802 22063 27858 22072
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 27620 21548 27672 21554
rect 27620 21490 27672 21496
rect 27252 21072 27304 21078
rect 27252 21014 27304 21020
rect 27264 20534 27292 21014
rect 27356 20806 27384 21490
rect 27712 21344 27764 21350
rect 27712 21286 27764 21292
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 27724 20806 27752 21286
rect 27816 21078 27844 21286
rect 27804 21072 27856 21078
rect 27804 21014 27856 21020
rect 27802 20904 27858 20913
rect 27802 20839 27858 20848
rect 27344 20800 27396 20806
rect 27344 20742 27396 20748
rect 27712 20800 27764 20806
rect 27712 20742 27764 20748
rect 27356 20602 27752 20618
rect 27344 20596 27764 20602
rect 27396 20590 27712 20596
rect 27344 20538 27396 20544
rect 27712 20538 27764 20544
rect 27252 20528 27304 20534
rect 27252 20470 27304 20476
rect 27436 20528 27488 20534
rect 27436 20470 27488 20476
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27356 19990 27384 20402
rect 27344 19984 27396 19990
rect 27344 19926 27396 19932
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27160 19168 27212 19174
rect 27160 19110 27212 19116
rect 27172 18766 27200 19110
rect 27356 18834 27384 19314
rect 27448 19310 27476 20470
rect 27528 20460 27580 20466
rect 27528 20402 27580 20408
rect 27540 19514 27568 20402
rect 27620 20324 27672 20330
rect 27620 20266 27672 20272
rect 27712 20324 27764 20330
rect 27712 20266 27764 20272
rect 27528 19508 27580 19514
rect 27528 19450 27580 19456
rect 27632 19310 27660 20266
rect 27724 19922 27752 20266
rect 27712 19916 27764 19922
rect 27712 19858 27764 19864
rect 27816 19802 27844 20839
rect 27896 19984 27948 19990
rect 27896 19926 27948 19932
rect 27724 19774 27844 19802
rect 27436 19304 27488 19310
rect 27620 19304 27672 19310
rect 27488 19264 27568 19292
rect 27436 19246 27488 19252
rect 27344 18828 27396 18834
rect 27344 18770 27396 18776
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 27540 18698 27568 19264
rect 27618 19272 27620 19281
rect 27672 19272 27674 19281
rect 27618 19207 27674 19216
rect 27528 18692 27580 18698
rect 27528 18634 27580 18640
rect 27436 18420 27488 18426
rect 27436 18362 27488 18368
rect 27160 18284 27212 18290
rect 27080 18244 27160 18272
rect 26884 17128 26936 17134
rect 26884 17070 26936 17076
rect 26896 16726 26924 17070
rect 26884 16720 26936 16726
rect 26884 16662 26936 16668
rect 26884 16584 26936 16590
rect 26884 16526 26936 16532
rect 26896 16250 26924 16526
rect 26884 16244 26936 16250
rect 26884 16186 26936 16192
rect 26884 15496 26936 15502
rect 26884 15438 26936 15444
rect 26896 15366 26924 15438
rect 26884 15360 26936 15366
rect 26884 15302 26936 15308
rect 26790 14784 26846 14793
rect 26790 14719 26846 14728
rect 26804 12434 26832 14719
rect 26896 14074 26924 15302
rect 26988 15094 27016 18226
rect 27080 17270 27108 18244
rect 27160 18226 27212 18232
rect 27172 18057 27200 18226
rect 27158 18048 27214 18057
rect 27158 17983 27214 17992
rect 27068 17264 27120 17270
rect 27068 17206 27120 17212
rect 27448 16674 27476 18362
rect 27724 18358 27752 19774
rect 27802 19408 27858 19417
rect 27802 19343 27858 19352
rect 27712 18352 27764 18358
rect 27712 18294 27764 18300
rect 27448 16646 27568 16674
rect 27436 16448 27488 16454
rect 27436 16390 27488 16396
rect 27068 16040 27120 16046
rect 27068 15982 27120 15988
rect 26976 15088 27028 15094
rect 26976 15030 27028 15036
rect 27080 14414 27108 15982
rect 27160 15020 27212 15026
rect 27160 14962 27212 14968
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 27172 14278 27200 14962
rect 27160 14272 27212 14278
rect 27160 14214 27212 14220
rect 27344 14272 27396 14278
rect 27344 14214 27396 14220
rect 26884 14068 26936 14074
rect 26884 14010 26936 14016
rect 27252 14000 27304 14006
rect 27252 13942 27304 13948
rect 27264 13394 27292 13942
rect 27252 13388 27304 13394
rect 27252 13330 27304 13336
rect 27068 12844 27120 12850
rect 27068 12786 27120 12792
rect 26804 12406 26924 12434
rect 26792 10464 26844 10470
rect 26790 10432 26792 10441
rect 26844 10432 26846 10441
rect 26790 10367 26846 10376
rect 26700 9444 26752 9450
rect 26700 9386 26752 9392
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 25964 8560 26016 8566
rect 25964 8502 26016 8508
rect 26424 8424 26476 8430
rect 26054 8392 26110 8401
rect 26424 8366 26476 8372
rect 26054 8327 26110 8336
rect 25792 8044 25912 8072
rect 25780 7812 25832 7818
rect 25780 7754 25832 7760
rect 25608 6854 25728 6882
rect 25596 6724 25648 6730
rect 25596 6666 25648 6672
rect 25608 6390 25636 6666
rect 25596 6384 25648 6390
rect 25596 6326 25648 6332
rect 25504 6316 25556 6322
rect 25504 6258 25556 6264
rect 25700 6254 25728 6854
rect 25792 6458 25820 7754
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 25594 5808 25650 5817
rect 25594 5743 25596 5752
rect 25648 5743 25650 5752
rect 25596 5714 25648 5720
rect 25780 5704 25832 5710
rect 25778 5672 25780 5681
rect 25832 5672 25834 5681
rect 25778 5607 25834 5616
rect 25884 5574 25912 8044
rect 26068 6322 26096 8327
rect 26436 7818 26464 8366
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26424 7812 26476 7818
rect 26424 7754 26476 7760
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 26160 6458 26188 7686
rect 26148 6452 26200 6458
rect 26148 6394 26200 6400
rect 26056 6316 26108 6322
rect 26056 6258 26108 6264
rect 26436 6254 26464 7754
rect 26804 7002 26832 8230
rect 26608 6996 26660 7002
rect 26608 6938 26660 6944
rect 26792 6996 26844 7002
rect 26792 6938 26844 6944
rect 26514 6488 26570 6497
rect 26514 6423 26570 6432
rect 25964 6248 26016 6254
rect 25964 6190 26016 6196
rect 26424 6248 26476 6254
rect 26424 6190 26476 6196
rect 25976 5930 26004 6190
rect 25976 5914 26372 5930
rect 25976 5908 26384 5914
rect 25976 5902 26332 5908
rect 26332 5850 26384 5856
rect 25964 5704 26016 5710
rect 25964 5646 26016 5652
rect 25872 5568 25924 5574
rect 25872 5510 25924 5516
rect 25504 5296 25556 5302
rect 25872 5296 25924 5302
rect 25556 5256 25872 5284
rect 25504 5238 25556 5244
rect 25872 5238 25924 5244
rect 25504 4072 25556 4078
rect 25504 4014 25556 4020
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 25136 3596 25188 3602
rect 25136 3538 25188 3544
rect 24676 3460 24728 3466
rect 24676 3402 24728 3408
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24400 2848 24452 2854
rect 24400 2790 24452 2796
rect 23584 2746 23888 2774
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 23480 2372 23532 2378
rect 23480 2314 23532 2320
rect 23492 1170 23520 2314
rect 23492 1142 23612 1170
rect 23584 800 23612 1142
rect 23860 800 23888 2746
rect 24044 2746 24164 2774
rect 24228 2746 24348 2774
rect 24044 2106 24072 2746
rect 24228 2582 24256 2746
rect 24216 2576 24268 2582
rect 24216 2518 24268 2524
rect 24124 2304 24176 2310
rect 24124 2246 24176 2252
rect 24032 2100 24084 2106
rect 24032 2042 24084 2048
rect 24136 800 24164 2246
rect 24412 800 24440 2790
rect 24688 800 24716 3402
rect 24872 2922 24900 3538
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 24952 2916 25004 2922
rect 24952 2858 25004 2864
rect 24964 2650 24992 2858
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 24952 2508 25004 2514
rect 24952 2450 25004 2456
rect 24964 800 24992 2450
rect 25228 2304 25280 2310
rect 25228 2246 25280 2252
rect 25240 800 25268 2246
rect 25516 800 25544 4014
rect 25976 3641 26004 5646
rect 26436 4690 26464 6190
rect 26528 5166 26556 6423
rect 26620 5166 26648 6938
rect 26516 5160 26568 5166
rect 26516 5102 26568 5108
rect 26608 5160 26660 5166
rect 26608 5102 26660 5108
rect 26896 4690 26924 12406
rect 27080 10713 27108 12786
rect 27160 12300 27212 12306
rect 27160 12242 27212 12248
rect 27066 10704 27122 10713
rect 27066 10639 27122 10648
rect 26976 10532 27028 10538
rect 26976 10474 27028 10480
rect 26988 10441 27016 10474
rect 26974 10432 27030 10441
rect 26974 10367 27030 10376
rect 27080 9518 27108 10639
rect 27068 9512 27120 9518
rect 27068 9454 27120 9460
rect 27172 8022 27200 12242
rect 27264 11762 27292 13330
rect 27356 12850 27384 14214
rect 27448 13938 27476 16390
rect 27436 13932 27488 13938
rect 27436 13874 27488 13880
rect 27344 12844 27396 12850
rect 27344 12786 27396 12792
rect 27540 12434 27568 16646
rect 27356 12406 27568 12434
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 27160 8016 27212 8022
rect 27160 7958 27212 7964
rect 27356 7562 27384 12406
rect 27436 10600 27488 10606
rect 27436 10542 27488 10548
rect 27448 9722 27476 10542
rect 27620 10056 27672 10062
rect 27672 10016 27752 10044
rect 27620 9998 27672 10004
rect 27436 9716 27488 9722
rect 27436 9658 27488 9664
rect 27416 9580 27468 9586
rect 27468 9528 27476 9568
rect 27416 9522 27476 9528
rect 27448 9489 27476 9522
rect 27434 9480 27490 9489
rect 27724 9450 27752 10016
rect 27434 9415 27490 9424
rect 27620 9444 27672 9450
rect 27620 9386 27672 9392
rect 27712 9444 27764 9450
rect 27712 9386 27764 9392
rect 27528 8016 27580 8022
rect 27528 7958 27580 7964
rect 27080 7534 27384 7562
rect 26424 4684 26476 4690
rect 26424 4626 26476 4632
rect 26884 4684 26936 4690
rect 26884 4626 26936 4632
rect 26436 4146 26464 4626
rect 26424 4140 26476 4146
rect 26424 4082 26476 4088
rect 26988 4078 27016 4109
rect 26884 4072 26936 4078
rect 26976 4072 27028 4078
rect 26884 4014 26936 4020
rect 26974 4040 26976 4049
rect 27028 4040 27030 4049
rect 25962 3632 26018 3641
rect 26896 3602 26924 4014
rect 26974 3975 27030 3984
rect 26988 3670 27016 3975
rect 26976 3664 27028 3670
rect 26976 3606 27028 3612
rect 25962 3567 26018 3576
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 26056 2984 26108 2990
rect 26056 2926 26108 2932
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 25780 2372 25832 2378
rect 25780 2314 25832 2320
rect 25792 800 25820 2314
rect 26068 800 26096 2926
rect 26436 2774 26464 2926
rect 26344 2746 26464 2774
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 26252 1698 26280 2382
rect 26240 1692 26292 1698
rect 26240 1634 26292 1640
rect 26344 800 26372 2746
rect 27080 2650 27108 7534
rect 27160 7404 27212 7410
rect 27160 7346 27212 7352
rect 27172 7313 27200 7346
rect 27158 7304 27214 7313
rect 27158 7239 27214 7248
rect 27160 6724 27212 6730
rect 27160 6666 27212 6672
rect 27172 6458 27200 6666
rect 27160 6452 27212 6458
rect 27160 6394 27212 6400
rect 27540 6322 27568 7958
rect 27632 6866 27660 9386
rect 27620 6860 27672 6866
rect 27620 6802 27672 6808
rect 27620 6656 27672 6662
rect 27620 6598 27672 6604
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27632 6254 27660 6598
rect 27724 6497 27752 9386
rect 27816 9178 27844 19343
rect 27908 19242 27936 19926
rect 27896 19236 27948 19242
rect 27896 19178 27948 19184
rect 27908 17610 27936 19178
rect 28078 18864 28134 18873
rect 28078 18799 28080 18808
rect 28132 18799 28134 18808
rect 28080 18770 28132 18776
rect 28080 18624 28132 18630
rect 28080 18566 28132 18572
rect 28092 18290 28120 18566
rect 28080 18284 28132 18290
rect 28080 18226 28132 18232
rect 27988 17740 28040 17746
rect 27988 17682 28040 17688
rect 27896 17604 27948 17610
rect 27896 17546 27948 17552
rect 27896 12096 27948 12102
rect 27896 12038 27948 12044
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 27710 6488 27766 6497
rect 27710 6423 27766 6432
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 27620 5704 27672 5710
rect 27620 5646 27672 5652
rect 27252 5024 27304 5030
rect 27252 4966 27304 4972
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 27172 3534 27200 3878
rect 27160 3528 27212 3534
rect 27160 3470 27212 3476
rect 27264 2774 27292 4966
rect 27632 4622 27660 5646
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 27620 4616 27672 4622
rect 27620 4558 27672 4564
rect 27172 2746 27292 2774
rect 27068 2644 27120 2650
rect 27068 2586 27120 2592
rect 26608 2372 26660 2378
rect 26608 2314 26660 2320
rect 26884 2372 26936 2378
rect 26884 2314 26936 2320
rect 26620 800 26648 2314
rect 26896 800 26924 2314
rect 27172 800 27200 2746
rect 27448 800 27476 4558
rect 27632 3398 27660 4558
rect 27620 3392 27672 3398
rect 27620 3334 27672 3340
rect 27712 2916 27764 2922
rect 27712 2858 27764 2864
rect 27724 800 27752 2858
rect 27908 2582 27936 12038
rect 28000 2938 28028 17682
rect 28080 13728 28132 13734
rect 28080 13670 28132 13676
rect 28092 12850 28120 13670
rect 28080 12844 28132 12850
rect 28080 12786 28132 12792
rect 28184 12170 28212 22494
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28276 19145 28304 19314
rect 28262 19136 28318 19145
rect 28262 19071 28318 19080
rect 28264 18624 28316 18630
rect 28264 18566 28316 18572
rect 28276 16425 28304 18566
rect 28368 17513 28396 20878
rect 28460 20806 28488 25910
rect 29092 25832 29144 25838
rect 29092 25774 29144 25780
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 28540 25152 28592 25158
rect 28540 25094 28592 25100
rect 28552 23118 28580 25094
rect 28908 24744 28960 24750
rect 28908 24686 28960 24692
rect 28920 24614 28948 24686
rect 28908 24608 28960 24614
rect 28908 24550 28960 24556
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28540 22636 28592 22642
rect 28540 22578 28592 22584
rect 28552 20942 28580 22578
rect 28920 21486 28948 24550
rect 29012 24410 29040 25230
rect 29104 25226 29132 25774
rect 29460 25288 29512 25294
rect 29460 25230 29512 25236
rect 29092 25220 29144 25226
rect 29092 25162 29144 25168
rect 29104 24614 29132 25162
rect 29092 24608 29144 24614
rect 29092 24550 29144 24556
rect 29000 24404 29052 24410
rect 29000 24346 29052 24352
rect 29012 23730 29040 24346
rect 29000 23724 29052 23730
rect 29000 23666 29052 23672
rect 29104 23526 29132 24550
rect 29092 23520 29144 23526
rect 29092 23462 29144 23468
rect 29368 22772 29420 22778
rect 29368 22714 29420 22720
rect 29000 22704 29052 22710
rect 29000 22646 29052 22652
rect 28908 21480 28960 21486
rect 28908 21422 28960 21428
rect 28540 20936 28592 20942
rect 28816 20936 28868 20942
rect 28592 20896 28672 20924
rect 28540 20878 28592 20884
rect 28448 20800 28500 20806
rect 28448 20742 28500 20748
rect 28540 20528 28592 20534
rect 28540 20470 28592 20476
rect 28552 20058 28580 20470
rect 28644 20330 28672 20896
rect 28814 20904 28816 20913
rect 28868 20904 28870 20913
rect 28814 20839 28870 20848
rect 28816 20392 28868 20398
rect 28816 20334 28868 20340
rect 28632 20324 28684 20330
rect 28632 20266 28684 20272
rect 28540 20052 28592 20058
rect 28540 19994 28592 20000
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28460 18601 28488 19790
rect 28538 19544 28594 19553
rect 28538 19479 28540 19488
rect 28592 19479 28594 19488
rect 28540 19450 28592 19456
rect 28538 19408 28594 19417
rect 28538 19343 28540 19352
rect 28592 19343 28594 19352
rect 28540 19314 28592 19320
rect 28644 19242 28672 20266
rect 28828 19854 28856 20334
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28724 19712 28776 19718
rect 28724 19654 28776 19660
rect 28632 19236 28684 19242
rect 28632 19178 28684 19184
rect 28632 18964 28684 18970
rect 28632 18906 28684 18912
rect 28540 18828 28592 18834
rect 28540 18770 28592 18776
rect 28446 18592 28502 18601
rect 28446 18527 28502 18536
rect 28354 17504 28410 17513
rect 28354 17439 28410 17448
rect 28262 16416 28318 16425
rect 28262 16351 28318 16360
rect 28172 12164 28224 12170
rect 28172 12106 28224 12112
rect 28460 12102 28488 18527
rect 28552 18057 28580 18770
rect 28538 18048 28594 18057
rect 28538 17983 28594 17992
rect 28552 16726 28580 17983
rect 28540 16720 28592 16726
rect 28540 16662 28592 16668
rect 28644 14074 28672 18906
rect 28736 18306 28764 19654
rect 28816 18964 28868 18970
rect 28816 18906 28868 18912
rect 28828 18465 28856 18906
rect 28814 18456 28870 18465
rect 28814 18391 28870 18400
rect 28920 18358 28948 21422
rect 29012 19378 29040 22646
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 29182 19544 29238 19553
rect 29182 19479 29238 19488
rect 29090 19408 29146 19417
rect 29000 19372 29052 19378
rect 29090 19343 29146 19352
rect 29000 19314 29052 19320
rect 29104 19242 29132 19343
rect 29092 19236 29144 19242
rect 29092 19178 29144 19184
rect 28908 18352 28960 18358
rect 28736 18290 28856 18306
rect 28908 18294 28960 18300
rect 28736 18284 28868 18290
rect 28736 18278 28816 18284
rect 28816 18226 28868 18232
rect 28920 17270 28948 18294
rect 29000 18216 29052 18222
rect 28998 18184 29000 18193
rect 29052 18184 29054 18193
rect 28998 18119 29054 18128
rect 29196 18086 29224 19479
rect 29184 18080 29236 18086
rect 29184 18022 29236 18028
rect 29196 17678 29224 18022
rect 29184 17672 29236 17678
rect 29184 17614 29236 17620
rect 29092 17604 29144 17610
rect 29092 17546 29144 17552
rect 28908 17264 28960 17270
rect 28908 17206 28960 17212
rect 28920 16114 28948 17206
rect 28908 16108 28960 16114
rect 28908 16050 28960 16056
rect 28632 14068 28684 14074
rect 28632 14010 28684 14016
rect 28920 14006 28948 16050
rect 29104 15450 29132 17546
rect 29196 17105 29224 17614
rect 29182 17096 29238 17105
rect 29182 17031 29238 17040
rect 29104 15422 29224 15450
rect 29288 15434 29316 21966
rect 29380 21146 29408 22714
rect 29472 21146 29500 25230
rect 29564 22094 29592 33254
rect 29656 24274 29684 39238
rect 29840 31142 29868 60454
rect 29920 57452 29972 57458
rect 29920 57394 29972 57400
rect 29932 56846 29960 57394
rect 29920 56840 29972 56846
rect 29920 56782 29972 56788
rect 29932 56370 29960 56782
rect 29920 56364 29972 56370
rect 29920 56306 29972 56312
rect 29828 31136 29880 31142
rect 29828 31078 29880 31084
rect 29736 30660 29788 30666
rect 29736 30602 29788 30608
rect 29748 24342 29776 30602
rect 29828 25968 29880 25974
rect 29828 25910 29880 25916
rect 29840 25294 29868 25910
rect 29828 25288 29880 25294
rect 29880 25248 29960 25276
rect 29828 25230 29880 25236
rect 29932 24886 29960 25248
rect 29920 24880 29972 24886
rect 29920 24822 29972 24828
rect 29828 24812 29880 24818
rect 29828 24754 29880 24760
rect 29736 24336 29788 24342
rect 29736 24278 29788 24284
rect 29644 24268 29696 24274
rect 29644 24210 29696 24216
rect 29656 23118 29684 24210
rect 29736 23656 29788 23662
rect 29736 23598 29788 23604
rect 29644 23112 29696 23118
rect 29644 23054 29696 23060
rect 29642 22944 29698 22953
rect 29642 22879 29698 22888
rect 29656 22642 29684 22879
rect 29644 22636 29696 22642
rect 29644 22578 29696 22584
rect 29748 22098 29776 23598
rect 29840 23322 29868 24754
rect 30024 24410 30052 60998
rect 30300 60722 30328 63200
rect 31036 61198 31064 63200
rect 31772 61198 31800 63200
rect 32508 61198 32536 63200
rect 33244 61198 33272 63200
rect 31024 61192 31076 61198
rect 31024 61134 31076 61140
rect 31760 61192 31812 61198
rect 31760 61134 31812 61140
rect 32496 61192 32548 61198
rect 32496 61134 32548 61140
rect 33232 61192 33284 61198
rect 33232 61134 33284 61140
rect 31668 61124 31720 61130
rect 31668 61066 31720 61072
rect 31024 61056 31076 61062
rect 31024 60998 31076 61004
rect 30288 60716 30340 60722
rect 30288 60658 30340 60664
rect 30564 60512 30616 60518
rect 30564 60454 30616 60460
rect 30380 57248 30432 57254
rect 30380 57190 30432 57196
rect 30392 27878 30420 57190
rect 30472 56160 30524 56166
rect 30472 56102 30524 56108
rect 30484 30802 30512 56102
rect 30576 42838 30604 60454
rect 30748 57928 30800 57934
rect 30748 57870 30800 57876
rect 30760 57458 30788 57870
rect 31036 57458 31064 60998
rect 31680 59430 31708 61066
rect 31944 61056 31996 61062
rect 31944 60998 31996 61004
rect 33232 61056 33284 61062
rect 33232 60998 33284 61004
rect 33324 61056 33376 61062
rect 33324 60998 33376 61004
rect 31668 59424 31720 59430
rect 31668 59366 31720 59372
rect 31956 57934 31984 60998
rect 33244 60761 33272 60998
rect 33336 60897 33364 60998
rect 33322 60888 33378 60897
rect 33322 60823 33378 60832
rect 33980 60790 34008 63200
rect 34716 61198 34744 63200
rect 35820 62098 35848 63294
rect 36174 63294 36400 63322
rect 36174 63200 36230 63294
rect 35820 62070 35940 62098
rect 34934 61500 35242 61509
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61435 35242 61444
rect 35912 61198 35940 62070
rect 34704 61192 34756 61198
rect 34704 61134 34756 61140
rect 35900 61192 35952 61198
rect 35900 61134 35952 61140
rect 35072 61056 35124 61062
rect 35072 60998 35124 61004
rect 35992 61056 36044 61062
rect 35992 60998 36044 61004
rect 33968 60784 34020 60790
rect 33230 60752 33286 60761
rect 35084 60761 35112 60998
rect 33968 60726 34020 60732
rect 35070 60752 35126 60761
rect 33230 60687 33286 60696
rect 35070 60687 35126 60696
rect 34244 60512 34296 60518
rect 34244 60454 34296 60460
rect 33692 59424 33744 59430
rect 33692 59366 33744 59372
rect 31852 57928 31904 57934
rect 31852 57870 31904 57876
rect 31944 57928 31996 57934
rect 31944 57870 31996 57876
rect 32220 57928 32272 57934
rect 32220 57870 32272 57876
rect 32496 57928 32548 57934
rect 32496 57870 32548 57876
rect 32680 57928 32732 57934
rect 32680 57870 32732 57876
rect 31484 57792 31536 57798
rect 31484 57734 31536 57740
rect 30748 57452 30800 57458
rect 30748 57394 30800 57400
rect 31024 57452 31076 57458
rect 31024 57394 31076 57400
rect 31116 57452 31168 57458
rect 31116 57394 31168 57400
rect 31392 57452 31444 57458
rect 31392 57394 31444 57400
rect 30564 42832 30616 42838
rect 30564 42774 30616 42780
rect 31128 31210 31156 57394
rect 31404 57254 31432 57394
rect 31392 57248 31444 57254
rect 31392 57190 31444 57196
rect 31404 55962 31432 57190
rect 31392 55956 31444 55962
rect 31392 55898 31444 55904
rect 31496 44946 31524 57734
rect 31576 57452 31628 57458
rect 31576 57394 31628 57400
rect 31588 57050 31616 57394
rect 31576 57044 31628 57050
rect 31576 56986 31628 56992
rect 31484 44940 31536 44946
rect 31484 44882 31536 44888
rect 31864 42702 31892 57870
rect 32232 57526 32260 57870
rect 32220 57520 32272 57526
rect 32220 57462 32272 57468
rect 32508 57254 32536 57870
rect 32496 57248 32548 57254
rect 32496 57190 32548 57196
rect 32692 56914 32720 57870
rect 32680 56908 32732 56914
rect 32680 56850 32732 56856
rect 33600 56364 33652 56370
rect 33600 56306 33652 56312
rect 33612 55894 33640 56306
rect 33600 55888 33652 55894
rect 33600 55830 33652 55836
rect 32220 42832 32272 42838
rect 32220 42774 32272 42780
rect 31852 42696 31904 42702
rect 31852 42638 31904 42644
rect 31760 42628 31812 42634
rect 31760 42570 31812 42576
rect 31772 39302 31800 42570
rect 31864 41478 31892 42638
rect 31852 41472 31904 41478
rect 31852 41414 31904 41420
rect 31760 39296 31812 39302
rect 31760 39238 31812 39244
rect 32128 33516 32180 33522
rect 32128 33458 32180 33464
rect 31760 31748 31812 31754
rect 31760 31690 31812 31696
rect 31116 31204 31168 31210
rect 31116 31146 31168 31152
rect 31128 30802 31156 31146
rect 30472 30796 30524 30802
rect 30472 30738 30524 30744
rect 31116 30796 31168 30802
rect 31116 30738 31168 30744
rect 31772 30734 31800 31690
rect 32036 31680 32088 31686
rect 32036 31622 32088 31628
rect 32048 31346 32076 31622
rect 32036 31340 32088 31346
rect 32036 31282 32088 31288
rect 31760 30728 31812 30734
rect 31760 30670 31812 30676
rect 31300 29164 31352 29170
rect 31300 29106 31352 29112
rect 31024 29096 31076 29102
rect 31024 29038 31076 29044
rect 30380 27872 30432 27878
rect 30380 27814 30432 27820
rect 30196 25356 30248 25362
rect 30196 25298 30248 25304
rect 30104 25152 30156 25158
rect 30104 25094 30156 25100
rect 30012 24404 30064 24410
rect 30012 24346 30064 24352
rect 29920 24336 29972 24342
rect 29920 24278 29972 24284
rect 29932 23866 29960 24278
rect 29920 23860 29972 23866
rect 29920 23802 29972 23808
rect 30116 23798 30144 25094
rect 30104 23792 30156 23798
rect 30104 23734 30156 23740
rect 30104 23656 30156 23662
rect 30104 23598 30156 23604
rect 29828 23316 29880 23322
rect 29828 23258 29880 23264
rect 30116 23254 30144 23598
rect 29920 23248 29972 23254
rect 29920 23190 29972 23196
rect 30104 23248 30156 23254
rect 30104 23190 30156 23196
rect 29932 23089 29960 23190
rect 30208 23118 30236 25298
rect 30472 24608 30524 24614
rect 30840 24608 30892 24614
rect 30524 24556 30604 24562
rect 30472 24550 30604 24556
rect 30840 24550 30892 24556
rect 30484 24534 30604 24550
rect 30196 23112 30248 23118
rect 29918 23080 29974 23089
rect 30380 23112 30432 23118
rect 30196 23054 30248 23060
rect 30378 23080 30380 23089
rect 30432 23080 30434 23089
rect 29918 23015 29974 23024
rect 30378 23015 30434 23024
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 30392 22506 30420 22578
rect 30380 22500 30432 22506
rect 30380 22442 30432 22448
rect 30472 22500 30524 22506
rect 30472 22442 30524 22448
rect 29564 22066 29684 22094
rect 29368 21140 29420 21146
rect 29368 21082 29420 21088
rect 29460 21140 29512 21146
rect 29460 21082 29512 21088
rect 29472 20466 29500 21082
rect 29460 20460 29512 20466
rect 29460 20402 29512 20408
rect 29472 19922 29500 20402
rect 29460 19916 29512 19922
rect 29460 19858 29512 19864
rect 29458 19544 29514 19553
rect 29458 19479 29514 19488
rect 29472 19378 29500 19479
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29458 17640 29514 17649
rect 29458 17575 29460 17584
rect 29512 17575 29514 17584
rect 29460 17546 29512 17552
rect 29460 17264 29512 17270
rect 29460 17206 29512 17212
rect 29368 16720 29420 16726
rect 29366 16688 29368 16697
rect 29420 16688 29422 16697
rect 29366 16623 29422 16632
rect 29472 15706 29500 17206
rect 29552 16992 29604 16998
rect 29552 16934 29604 16940
rect 29564 16182 29592 16934
rect 29552 16176 29604 16182
rect 29552 16118 29604 16124
rect 29460 15700 29512 15706
rect 29460 15642 29512 15648
rect 29092 15360 29144 15366
rect 29092 15302 29144 15308
rect 29104 14414 29132 15302
rect 29196 14414 29224 15422
rect 29276 15428 29328 15434
rect 29276 15370 29328 15376
rect 29276 14476 29328 14482
rect 29276 14418 29328 14424
rect 29092 14408 29144 14414
rect 29092 14350 29144 14356
rect 29184 14408 29236 14414
rect 29184 14350 29236 14356
rect 28908 14000 28960 14006
rect 28908 13942 28960 13948
rect 28724 13864 28776 13870
rect 28724 13806 28776 13812
rect 28736 13190 28764 13806
rect 29000 13728 29052 13734
rect 29000 13670 29052 13676
rect 29012 13326 29040 13670
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 29104 12918 29132 14350
rect 29092 12912 29144 12918
rect 29092 12854 29144 12860
rect 29000 12708 29052 12714
rect 29000 12650 29052 12656
rect 28448 12096 28500 12102
rect 28448 12038 28500 12044
rect 28172 11756 28224 11762
rect 28172 11698 28224 11704
rect 28184 10538 28212 11698
rect 28448 11620 28500 11626
rect 28448 11562 28500 11568
rect 28460 11150 28488 11562
rect 29012 11370 29040 12650
rect 29092 12164 29144 12170
rect 29092 12106 29144 12112
rect 28828 11342 29040 11370
rect 28448 11144 28500 11150
rect 28828 11098 28856 11342
rect 29000 11212 29052 11218
rect 29000 11154 29052 11160
rect 28448 11086 28500 11092
rect 28264 11076 28316 11082
rect 28264 11018 28316 11024
rect 28736 11070 28856 11098
rect 28172 10532 28224 10538
rect 28172 10474 28224 10480
rect 28184 9586 28212 10474
rect 28172 9580 28224 9586
rect 28172 9522 28224 9528
rect 28170 9480 28226 9489
rect 28170 9415 28226 9424
rect 28184 9382 28212 9415
rect 28080 9376 28132 9382
rect 28080 9318 28132 9324
rect 28172 9376 28224 9382
rect 28172 9318 28224 9324
rect 28092 9178 28120 9318
rect 28080 9172 28132 9178
rect 28080 9114 28132 9120
rect 28080 8492 28132 8498
rect 28080 8434 28132 8440
rect 28092 7750 28120 8434
rect 28080 7744 28132 7750
rect 28080 7686 28132 7692
rect 28092 7410 28120 7686
rect 28080 7404 28132 7410
rect 28080 7346 28132 7352
rect 28172 6860 28224 6866
rect 28172 6802 28224 6808
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 28092 6322 28120 6734
rect 28080 6316 28132 6322
rect 28080 6258 28132 6264
rect 28092 5234 28120 6258
rect 28184 5846 28212 6802
rect 28276 6458 28304 11018
rect 28356 11008 28408 11014
rect 28356 10950 28408 10956
rect 28368 10674 28396 10950
rect 28540 10804 28592 10810
rect 28540 10746 28592 10752
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 28552 9926 28580 10746
rect 28632 10736 28684 10742
rect 28632 10678 28684 10684
rect 28644 10266 28672 10678
rect 28632 10260 28684 10266
rect 28632 10202 28684 10208
rect 28540 9920 28592 9926
rect 28540 9862 28592 9868
rect 28356 8288 28408 8294
rect 28356 8230 28408 8236
rect 28264 6452 28316 6458
rect 28264 6394 28316 6400
rect 28172 5840 28224 5846
rect 28172 5782 28224 5788
rect 28368 5710 28396 8230
rect 28736 7818 28764 11070
rect 28724 7812 28776 7818
rect 28724 7754 28776 7760
rect 28540 7336 28592 7342
rect 28540 7278 28592 7284
rect 28632 7336 28684 7342
rect 28632 7278 28684 7284
rect 28356 5704 28408 5710
rect 28356 5646 28408 5652
rect 28356 5568 28408 5574
rect 28356 5510 28408 5516
rect 28368 5234 28396 5510
rect 28080 5228 28132 5234
rect 28080 5170 28132 5176
rect 28356 5228 28408 5234
rect 28356 5170 28408 5176
rect 28092 3058 28120 5170
rect 28552 4554 28580 7278
rect 28644 7041 28672 7278
rect 28630 7032 28686 7041
rect 28630 6967 28686 6976
rect 28644 6798 28672 6967
rect 28632 6792 28684 6798
rect 28632 6734 28684 6740
rect 28632 5772 28684 5778
rect 28632 5714 28684 5720
rect 28644 5681 28672 5714
rect 28630 5672 28686 5681
rect 28630 5607 28686 5616
rect 28448 4548 28500 4554
rect 28448 4490 28500 4496
rect 28540 4548 28592 4554
rect 28540 4490 28592 4496
rect 28264 4480 28316 4486
rect 28264 4422 28316 4428
rect 28172 3528 28224 3534
rect 28172 3470 28224 3476
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 28000 2910 28120 2938
rect 27988 2848 28040 2854
rect 27988 2790 28040 2796
rect 27896 2576 27948 2582
rect 27896 2518 27948 2524
rect 28000 800 28028 2790
rect 28092 2514 28120 2910
rect 28080 2508 28132 2514
rect 28080 2450 28132 2456
rect 28184 2446 28212 3470
rect 28172 2440 28224 2446
rect 28172 2382 28224 2388
rect 28276 800 28304 4422
rect 28356 3460 28408 3466
rect 28356 3402 28408 3408
rect 28368 1970 28396 3402
rect 28460 2774 28488 4490
rect 28552 4146 28580 4490
rect 28736 4146 28764 7754
rect 28908 6656 28960 6662
rect 28908 6598 28960 6604
rect 28920 6254 28948 6598
rect 29012 6458 29040 11154
rect 29104 11014 29132 12106
rect 29288 11762 29316 14418
rect 29276 11756 29328 11762
rect 29276 11698 29328 11704
rect 29472 11082 29500 15642
rect 29460 11076 29512 11082
rect 29460 11018 29512 11024
rect 29092 11008 29144 11014
rect 29092 10950 29144 10956
rect 29104 10470 29132 10950
rect 29274 10704 29330 10713
rect 29274 10639 29276 10648
rect 29328 10639 29330 10648
rect 29460 10668 29512 10674
rect 29276 10610 29328 10616
rect 29460 10610 29512 10616
rect 29092 10464 29144 10470
rect 29092 10406 29144 10412
rect 29368 10464 29420 10470
rect 29368 10406 29420 10412
rect 29104 9926 29132 10406
rect 29184 10192 29236 10198
rect 29184 10134 29236 10140
rect 29092 9920 29144 9926
rect 29092 9862 29144 9868
rect 29196 9761 29224 10134
rect 29182 9752 29238 9761
rect 29238 9710 29316 9738
rect 29182 9687 29238 9696
rect 29184 8356 29236 8362
rect 29184 8298 29236 8304
rect 29196 6866 29224 8298
rect 29184 6860 29236 6866
rect 29184 6802 29236 6808
rect 29288 6746 29316 9710
rect 29380 9654 29408 10406
rect 29472 9926 29500 10610
rect 29656 9994 29684 22066
rect 29736 22092 29788 22098
rect 29736 22034 29788 22040
rect 30012 22024 30064 22030
rect 30010 21992 30012 22001
rect 30064 21992 30066 22001
rect 30010 21927 30066 21936
rect 29828 21888 29880 21894
rect 29828 21830 29880 21836
rect 30196 21888 30248 21894
rect 30196 21830 30248 21836
rect 29840 21622 29868 21830
rect 29736 21616 29788 21622
rect 29736 21558 29788 21564
rect 29828 21616 29880 21622
rect 29828 21558 29880 21564
rect 29748 21162 29776 21558
rect 30208 21554 30236 21830
rect 30196 21548 30248 21554
rect 30196 21490 30248 21496
rect 30380 21412 30432 21418
rect 30380 21354 30432 21360
rect 29748 21146 29960 21162
rect 29748 21140 29972 21146
rect 29748 21134 29920 21140
rect 29920 21082 29972 21088
rect 30392 20942 30420 21354
rect 30380 20936 30432 20942
rect 30380 20878 30432 20884
rect 30484 20874 30512 22442
rect 30472 20868 30524 20874
rect 30472 20810 30524 20816
rect 30380 20528 30432 20534
rect 30576 20482 30604 24534
rect 30748 24404 30800 24410
rect 30748 24346 30800 24352
rect 30656 22092 30708 22098
rect 30656 22034 30708 22040
rect 30668 21690 30696 22034
rect 30656 21684 30708 21690
rect 30656 21626 30708 21632
rect 30380 20470 30432 20476
rect 29736 19780 29788 19786
rect 29736 19722 29788 19728
rect 29748 18426 29776 19722
rect 29828 19712 29880 19718
rect 29828 19654 29880 19660
rect 29840 19378 29868 19654
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 30392 18986 30420 20470
rect 30484 20454 30604 20482
rect 30484 19922 30512 20454
rect 30564 20324 30616 20330
rect 30564 20266 30616 20272
rect 30472 19916 30524 19922
rect 30472 19858 30524 19864
rect 30484 19174 30512 19858
rect 30472 19168 30524 19174
rect 30576 19145 30604 20266
rect 30760 19854 30788 24346
rect 30852 22642 30880 24550
rect 30932 24404 30984 24410
rect 30932 24346 30984 24352
rect 30944 23594 30972 24346
rect 30932 23588 30984 23594
rect 30932 23530 30984 23536
rect 31036 23474 31064 29038
rect 31116 24132 31168 24138
rect 31116 24074 31168 24080
rect 31128 23866 31156 24074
rect 31116 23860 31168 23866
rect 31116 23802 31168 23808
rect 31312 23730 31340 29106
rect 31852 28484 31904 28490
rect 31852 28426 31904 28432
rect 31864 28218 31892 28426
rect 31852 28212 31904 28218
rect 31852 28154 31904 28160
rect 31944 27532 31996 27538
rect 31944 27474 31996 27480
rect 31576 25696 31628 25702
rect 31576 25638 31628 25644
rect 31392 24880 31444 24886
rect 31392 24822 31444 24828
rect 31300 23724 31352 23730
rect 30944 23446 31064 23474
rect 31220 23684 31300 23712
rect 30840 22636 30892 22642
rect 30840 22578 30892 22584
rect 30944 22094 30972 23446
rect 31024 23112 31076 23118
rect 31024 23054 31076 23060
rect 31036 22778 31064 23054
rect 31024 22772 31076 22778
rect 31076 22732 31156 22760
rect 31024 22714 31076 22720
rect 31128 22098 31156 22732
rect 30852 22066 30972 22094
rect 31116 22092 31168 22098
rect 30852 20534 30880 22066
rect 31116 22034 31168 22040
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 30840 20528 30892 20534
rect 30840 20470 30892 20476
rect 30840 20392 30892 20398
rect 30840 20334 30892 20340
rect 30748 19848 30800 19854
rect 30748 19790 30800 19796
rect 30656 19712 30708 19718
rect 30656 19654 30708 19660
rect 30668 19310 30696 19654
rect 30656 19304 30708 19310
rect 30656 19246 30708 19252
rect 30472 19110 30524 19116
rect 30562 19136 30618 19145
rect 30562 19071 30618 19080
rect 30392 18958 30512 18986
rect 30484 18834 30512 18958
rect 30472 18828 30524 18834
rect 30472 18770 30524 18776
rect 30380 18760 30432 18766
rect 30380 18702 30432 18708
rect 30012 18692 30064 18698
rect 30012 18634 30064 18640
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 29734 17776 29790 17785
rect 29734 17711 29790 17720
rect 29748 17134 29776 17711
rect 30024 17649 30052 18634
rect 30392 18442 30420 18702
rect 30484 18578 30512 18770
rect 30576 18766 30604 19071
rect 30746 19000 30802 19009
rect 30746 18935 30802 18944
rect 30760 18834 30788 18935
rect 30852 18902 30880 20334
rect 30840 18896 30892 18902
rect 30840 18838 30892 18844
rect 30748 18828 30800 18834
rect 30748 18770 30800 18776
rect 30564 18760 30616 18766
rect 30944 18714 30972 21966
rect 31024 21140 31076 21146
rect 31024 21082 31076 21088
rect 31036 18766 31064 21082
rect 31116 19848 31168 19854
rect 31116 19790 31168 19796
rect 31128 19718 31156 19790
rect 31116 19712 31168 19718
rect 31116 19654 31168 19660
rect 31116 19236 31168 19242
rect 31116 19178 31168 19184
rect 30564 18702 30616 18708
rect 30668 18686 30972 18714
rect 31024 18760 31076 18766
rect 31024 18702 31076 18708
rect 30484 18550 30604 18578
rect 30392 18414 30512 18442
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 30104 17808 30156 17814
rect 30288 17808 30340 17814
rect 30156 17768 30236 17796
rect 30104 17750 30156 17756
rect 30010 17640 30066 17649
rect 30208 17610 30236 17768
rect 30288 17750 30340 17756
rect 30010 17575 30066 17584
rect 30196 17604 30248 17610
rect 30196 17546 30248 17552
rect 30104 17536 30156 17542
rect 30104 17478 30156 17484
rect 30116 17377 30144 17478
rect 30102 17368 30158 17377
rect 30102 17303 30158 17312
rect 30196 17332 30248 17338
rect 30196 17274 30248 17280
rect 29828 17196 29880 17202
rect 29880 17156 29960 17184
rect 29828 17138 29880 17144
rect 29736 17128 29788 17134
rect 29736 17070 29788 17076
rect 29736 16992 29788 16998
rect 29736 16934 29788 16940
rect 29748 16590 29776 16934
rect 29828 16652 29880 16658
rect 29828 16594 29880 16600
rect 29736 16584 29788 16590
rect 29736 16526 29788 16532
rect 29736 15496 29788 15502
rect 29736 15438 29788 15444
rect 29748 14822 29776 15438
rect 29840 15026 29868 16594
rect 29932 15502 29960 17156
rect 30208 17066 30236 17274
rect 30196 17060 30248 17066
rect 30196 17002 30248 17008
rect 30300 16969 30328 17750
rect 30392 17542 30420 18226
rect 30484 18057 30512 18414
rect 30576 18068 30604 18550
rect 30668 18222 30696 18686
rect 30746 18456 30802 18465
rect 30746 18391 30802 18400
rect 30760 18222 30788 18391
rect 31024 18352 31076 18358
rect 31024 18294 31076 18300
rect 30656 18216 30708 18222
rect 30656 18158 30708 18164
rect 30748 18216 30800 18222
rect 30748 18158 30800 18164
rect 30838 18184 30894 18193
rect 30838 18119 30894 18128
rect 30748 18080 30800 18086
rect 30470 18048 30526 18057
rect 30576 18040 30696 18068
rect 30470 17983 30526 17992
rect 30380 17536 30432 17542
rect 30380 17478 30432 17484
rect 30380 17332 30432 17338
rect 30380 17274 30432 17280
rect 30286 16960 30342 16969
rect 30286 16895 30342 16904
rect 30392 16776 30420 17274
rect 30484 17202 30512 17983
rect 30562 17912 30618 17921
rect 30562 17847 30618 17856
rect 30576 17678 30604 17847
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 30564 17332 30616 17338
rect 30564 17274 30616 17280
rect 30472 17196 30524 17202
rect 30472 17138 30524 17144
rect 30472 16788 30524 16794
rect 30392 16748 30472 16776
rect 30472 16730 30524 16736
rect 30576 16522 30604 17274
rect 30564 16516 30616 16522
rect 30564 16458 30616 16464
rect 29920 15496 29972 15502
rect 29920 15438 29972 15444
rect 29828 15020 29880 15026
rect 29828 14962 29880 14968
rect 29736 14816 29788 14822
rect 29736 14758 29788 14764
rect 29748 14346 29776 14758
rect 29736 14340 29788 14346
rect 29736 14282 29788 14288
rect 29736 12096 29788 12102
rect 29736 12038 29788 12044
rect 29748 11830 29776 12038
rect 29736 11824 29788 11830
rect 29736 11766 29788 11772
rect 29828 11824 29880 11830
rect 29828 11766 29880 11772
rect 29736 10464 29788 10470
rect 29736 10406 29788 10412
rect 29748 10062 29776 10406
rect 29736 10056 29788 10062
rect 29736 9998 29788 10004
rect 29644 9988 29696 9994
rect 29644 9930 29696 9936
rect 29460 9920 29512 9926
rect 29460 9862 29512 9868
rect 29368 9648 29420 9654
rect 29368 9590 29420 9596
rect 29472 9586 29500 9862
rect 29552 9648 29604 9654
rect 29552 9590 29604 9596
rect 29460 9580 29512 9586
rect 29460 9522 29512 9528
rect 29564 9466 29592 9590
rect 29472 9438 29592 9466
rect 29472 8498 29500 9438
rect 29552 9376 29604 9382
rect 29552 9318 29604 9324
rect 29460 8492 29512 8498
rect 29460 8434 29512 8440
rect 29460 7744 29512 7750
rect 29460 7686 29512 7692
rect 29196 6718 29316 6746
rect 29000 6452 29052 6458
rect 29000 6394 29052 6400
rect 28908 6248 28960 6254
rect 28908 6190 28960 6196
rect 29000 5840 29052 5846
rect 29000 5782 29052 5788
rect 28908 5636 28960 5642
rect 28908 5578 28960 5584
rect 28816 5568 28868 5574
rect 28816 5510 28868 5516
rect 28540 4140 28592 4146
rect 28540 4082 28592 4088
rect 28724 4140 28776 4146
rect 28724 4082 28776 4088
rect 28540 3936 28592 3942
rect 28540 3878 28592 3884
rect 28552 3534 28580 3878
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 28460 2746 28580 2774
rect 28356 1964 28408 1970
rect 28356 1906 28408 1912
rect 28552 800 28580 2746
rect 28828 800 28856 5510
rect 28920 4622 28948 5578
rect 29012 5370 29040 5782
rect 29000 5364 29052 5370
rect 29000 5306 29052 5312
rect 29092 5092 29144 5098
rect 29092 5034 29144 5040
rect 29104 4758 29132 5034
rect 29092 4752 29144 4758
rect 29092 4694 29144 4700
rect 28908 4616 28960 4622
rect 28908 4558 28960 4564
rect 29000 4480 29052 4486
rect 29000 4422 29052 4428
rect 29092 4480 29144 4486
rect 29092 4422 29144 4428
rect 28906 3496 28962 3505
rect 28906 3431 28908 3440
rect 28960 3431 28962 3440
rect 28908 3402 28960 3408
rect 29012 2774 29040 4422
rect 29104 4214 29132 4422
rect 29092 4208 29144 4214
rect 29092 4150 29144 4156
rect 29012 2746 29132 2774
rect 29104 800 29132 2746
rect 29196 2514 29224 6718
rect 29472 5370 29500 7686
rect 29460 5364 29512 5370
rect 29460 5306 29512 5312
rect 29564 5166 29592 9318
rect 29736 8900 29788 8906
rect 29736 8842 29788 8848
rect 29748 8634 29776 8842
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 29552 5160 29604 5166
rect 29552 5102 29604 5108
rect 29564 4282 29592 5102
rect 29552 4276 29604 4282
rect 29552 4218 29604 4224
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 29276 3936 29328 3942
rect 29276 3878 29328 3884
rect 29288 3126 29316 3878
rect 29368 3596 29420 3602
rect 29368 3538 29420 3544
rect 29276 3120 29328 3126
rect 29276 3062 29328 3068
rect 29184 2508 29236 2514
rect 29184 2450 29236 2456
rect 29380 800 29408 3538
rect 29748 3534 29776 4014
rect 29840 3670 29868 11766
rect 29932 7478 29960 15438
rect 30104 15428 30156 15434
rect 30104 15370 30156 15376
rect 30012 14408 30064 14414
rect 30012 14350 30064 14356
rect 30024 13870 30052 14350
rect 30012 13864 30064 13870
rect 30012 13806 30064 13812
rect 30116 12238 30144 15370
rect 30196 15088 30248 15094
rect 30196 15030 30248 15036
rect 30208 14482 30236 15030
rect 30288 15020 30340 15026
rect 30288 14962 30340 14968
rect 30196 14476 30248 14482
rect 30196 14418 30248 14424
rect 30196 13796 30248 13802
rect 30196 13738 30248 13744
rect 30208 13138 30236 13738
rect 30300 13326 30328 14962
rect 30288 13320 30340 13326
rect 30288 13262 30340 13268
rect 30208 13110 30328 13138
rect 30196 12776 30248 12782
rect 30196 12718 30248 12724
rect 30208 12374 30236 12718
rect 30196 12368 30248 12374
rect 30196 12310 30248 12316
rect 30300 12306 30328 13110
rect 30576 12730 30604 16458
rect 30668 14618 30696 18040
rect 30748 18022 30800 18028
rect 30760 17746 30788 18022
rect 30748 17740 30800 17746
rect 30748 17682 30800 17688
rect 30852 17678 30880 18119
rect 31036 17921 31064 18294
rect 31128 18290 31156 19178
rect 31116 18284 31168 18290
rect 31116 18226 31168 18232
rect 31022 17912 31078 17921
rect 31022 17847 31078 17856
rect 30840 17672 30892 17678
rect 30840 17614 30892 17620
rect 30746 17368 30802 17377
rect 30746 17303 30802 17312
rect 30760 16454 30788 17303
rect 30748 16448 30800 16454
rect 30748 16390 30800 16396
rect 30656 14612 30708 14618
rect 30656 14554 30708 14560
rect 30852 14074 30880 17614
rect 30932 17128 30984 17134
rect 30932 17070 30984 17076
rect 30944 16697 30972 17070
rect 31036 16998 31064 17847
rect 31116 17672 31168 17678
rect 31116 17614 31168 17620
rect 31128 17066 31156 17614
rect 31116 17060 31168 17066
rect 31116 17002 31168 17008
rect 31024 16992 31076 16998
rect 31024 16934 31076 16940
rect 30930 16688 30986 16697
rect 30930 16623 30986 16632
rect 31036 16046 31064 16934
rect 31128 16561 31156 17002
rect 31114 16552 31170 16561
rect 31114 16487 31170 16496
rect 31024 16040 31076 16046
rect 31024 15982 31076 15988
rect 30932 14476 30984 14482
rect 30932 14418 30984 14424
rect 30840 14068 30892 14074
rect 30840 14010 30892 14016
rect 30746 13968 30802 13977
rect 30944 13938 30972 14418
rect 31036 14414 31064 15982
rect 31116 15020 31168 15026
rect 31116 14962 31168 14968
rect 31128 14618 31156 14962
rect 31116 14612 31168 14618
rect 31116 14554 31168 14560
rect 31024 14408 31076 14414
rect 31024 14350 31076 14356
rect 30746 13903 30802 13912
rect 30932 13932 30984 13938
rect 30760 13870 30788 13903
rect 30932 13874 30984 13880
rect 30748 13864 30800 13870
rect 30748 13806 30800 13812
rect 31116 13796 31168 13802
rect 31116 13738 31168 13744
rect 31128 13462 31156 13738
rect 31116 13456 31168 13462
rect 31116 13398 31168 13404
rect 30840 13252 30892 13258
rect 30840 13194 30892 13200
rect 30852 12986 30880 13194
rect 31116 13184 31168 13190
rect 31116 13126 31168 13132
rect 30840 12980 30892 12986
rect 30840 12922 30892 12928
rect 31128 12782 31156 13126
rect 31220 12986 31248 23684
rect 31300 23666 31352 23672
rect 31404 21554 31432 24822
rect 31588 23730 31616 25638
rect 31668 24744 31720 24750
rect 31668 24686 31720 24692
rect 31852 24744 31904 24750
rect 31852 24686 31904 24692
rect 31576 23724 31628 23730
rect 31576 23666 31628 23672
rect 31680 23526 31708 24686
rect 31760 23724 31812 23730
rect 31760 23666 31812 23672
rect 31668 23520 31720 23526
rect 31668 23462 31720 23468
rect 31484 22160 31536 22166
rect 31484 22102 31536 22108
rect 31392 21548 31444 21554
rect 31392 21490 31444 21496
rect 31300 21412 31352 21418
rect 31300 21354 31352 21360
rect 31312 21146 31340 21354
rect 31404 21146 31432 21490
rect 31300 21140 31352 21146
rect 31300 21082 31352 21088
rect 31392 21140 31444 21146
rect 31392 21082 31444 21088
rect 31392 19780 31444 19786
rect 31392 19722 31444 19728
rect 31300 19304 31352 19310
rect 31298 19272 31300 19281
rect 31352 19272 31354 19281
rect 31298 19207 31354 19216
rect 31298 18728 31354 18737
rect 31298 18663 31354 18672
rect 31312 18630 31340 18663
rect 31300 18624 31352 18630
rect 31300 18566 31352 18572
rect 31300 14476 31352 14482
rect 31300 14418 31352 14424
rect 31208 12980 31260 12986
rect 31208 12922 31260 12928
rect 31208 12844 31260 12850
rect 31312 12832 31340 14418
rect 31260 12804 31340 12832
rect 31208 12786 31260 12792
rect 31116 12776 31168 12782
rect 30576 12702 30788 12730
rect 31116 12718 31168 12724
rect 30656 12640 30708 12646
rect 30656 12582 30708 12588
rect 30288 12300 30340 12306
rect 30288 12242 30340 12248
rect 30104 12232 30156 12238
rect 30104 12174 30156 12180
rect 30196 12096 30248 12102
rect 30196 12038 30248 12044
rect 30288 12096 30340 12102
rect 30288 12038 30340 12044
rect 30104 11756 30156 11762
rect 30104 11698 30156 11704
rect 30010 9752 30066 9761
rect 30010 9687 30066 9696
rect 30024 9654 30052 9687
rect 30012 9648 30064 9654
rect 30012 9590 30064 9596
rect 30116 9586 30144 11698
rect 30208 11558 30236 12038
rect 30300 11830 30328 12038
rect 30288 11824 30340 11830
rect 30288 11766 30340 11772
rect 30196 11552 30248 11558
rect 30196 11494 30248 11500
rect 30562 10432 30618 10441
rect 30562 10367 30618 10376
rect 30472 10260 30524 10266
rect 30472 10202 30524 10208
rect 30484 10130 30512 10202
rect 30472 10124 30524 10130
rect 30472 10066 30524 10072
rect 30380 10056 30432 10062
rect 30380 9998 30432 10004
rect 30392 9722 30420 9998
rect 30380 9716 30432 9722
rect 30380 9658 30432 9664
rect 30378 9616 30434 9625
rect 30104 9580 30156 9586
rect 30104 9522 30156 9528
rect 30196 9580 30248 9586
rect 30378 9551 30434 9560
rect 30196 9522 30248 9528
rect 30116 9450 30144 9522
rect 30104 9444 30156 9450
rect 30104 9386 30156 9392
rect 30012 8560 30064 8566
rect 30012 8502 30064 8508
rect 29920 7472 29972 7478
rect 29920 7414 29972 7420
rect 30024 6458 30052 8502
rect 30012 6452 30064 6458
rect 30012 6394 30064 6400
rect 30104 6180 30156 6186
rect 30104 6122 30156 6128
rect 30116 4622 30144 6122
rect 30104 4616 30156 4622
rect 30104 4558 30156 4564
rect 30012 4548 30064 4554
rect 30012 4490 30064 4496
rect 30024 4146 30052 4490
rect 30208 4282 30236 9522
rect 30288 9512 30340 9518
rect 30286 9480 30288 9489
rect 30340 9480 30342 9489
rect 30286 9415 30342 9424
rect 30392 9178 30420 9551
rect 30380 9172 30432 9178
rect 30380 9114 30432 9120
rect 30472 9172 30524 9178
rect 30472 9114 30524 9120
rect 30392 8430 30420 9114
rect 30484 8974 30512 9114
rect 30472 8968 30524 8974
rect 30472 8910 30524 8916
rect 30484 8498 30512 8910
rect 30472 8492 30524 8498
rect 30472 8434 30524 8440
rect 30380 8424 30432 8430
rect 30380 8366 30432 8372
rect 30484 7954 30512 8434
rect 30472 7948 30524 7954
rect 30472 7890 30524 7896
rect 30576 6798 30604 10367
rect 30668 7698 30696 12582
rect 30760 10198 30788 12702
rect 31114 10704 31170 10713
rect 30932 10668 30984 10674
rect 31312 10690 31340 12804
rect 31170 10662 31340 10690
rect 31114 10639 31170 10648
rect 30932 10610 30984 10616
rect 30748 10192 30800 10198
rect 30748 10134 30800 10140
rect 30760 8634 30788 10134
rect 30944 10130 30972 10610
rect 30932 10124 30984 10130
rect 30932 10066 30984 10072
rect 30748 8628 30800 8634
rect 30748 8570 30800 8576
rect 30748 8492 30800 8498
rect 30748 8434 30800 8440
rect 30760 7886 30788 8434
rect 30748 7880 30800 7886
rect 30748 7822 30800 7828
rect 30840 7880 30892 7886
rect 30840 7822 30892 7828
rect 30668 7670 30788 7698
rect 30380 6792 30432 6798
rect 30380 6734 30432 6740
rect 30564 6792 30616 6798
rect 30564 6734 30616 6740
rect 30392 6338 30420 6734
rect 30300 6310 30420 6338
rect 30300 5710 30328 6310
rect 30288 5704 30340 5710
rect 30288 5646 30340 5652
rect 30472 5704 30524 5710
rect 30472 5646 30524 5652
rect 30484 5370 30512 5646
rect 30656 5568 30708 5574
rect 30656 5510 30708 5516
rect 30472 5364 30524 5370
rect 30472 5306 30524 5312
rect 30564 5228 30616 5234
rect 30564 5170 30616 5176
rect 30576 4826 30604 5170
rect 30564 4820 30616 4826
rect 30564 4762 30616 4768
rect 30668 4554 30696 5510
rect 30656 4548 30708 4554
rect 30656 4490 30708 4496
rect 30196 4276 30248 4282
rect 30196 4218 30248 4224
rect 30104 4208 30156 4214
rect 30104 4150 30156 4156
rect 30012 4140 30064 4146
rect 30012 4082 30064 4088
rect 29828 3664 29880 3670
rect 29828 3606 29880 3612
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 29748 2922 29776 3470
rect 29736 2916 29788 2922
rect 29736 2858 29788 2864
rect 30116 2446 30144 4150
rect 30288 3936 30340 3942
rect 30288 3878 30340 3884
rect 30300 3534 30328 3878
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 30196 3460 30248 3466
rect 30196 3402 30248 3408
rect 30104 2440 30156 2446
rect 30104 2382 30156 2388
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 29656 800 29684 2246
rect 29932 800 29960 2314
rect 30208 800 30236 3402
rect 30760 3126 30788 7670
rect 30852 7206 30880 7822
rect 30944 7546 30972 10066
rect 31128 9586 31156 10639
rect 31208 10056 31260 10062
rect 31208 9998 31260 10004
rect 31220 9722 31248 9998
rect 31300 9920 31352 9926
rect 31300 9862 31352 9868
rect 31208 9716 31260 9722
rect 31208 9658 31260 9664
rect 31208 9586 31260 9592
rect 31116 9580 31168 9586
rect 31208 9528 31260 9534
rect 31116 9522 31168 9528
rect 31220 9489 31248 9528
rect 31206 9480 31262 9489
rect 31206 9415 31262 9424
rect 31312 8974 31340 9862
rect 31404 9722 31432 19722
rect 31496 17202 31524 22102
rect 31680 22094 31708 23462
rect 31772 23186 31800 23666
rect 31864 23662 31892 24686
rect 31852 23656 31904 23662
rect 31852 23598 31904 23604
rect 31760 23180 31812 23186
rect 31760 23122 31812 23128
rect 31588 22066 31708 22094
rect 31588 22030 31616 22066
rect 31576 22024 31628 22030
rect 31576 21966 31628 21972
rect 31772 21962 31800 23122
rect 31760 21956 31812 21962
rect 31760 21898 31812 21904
rect 31576 21548 31628 21554
rect 31576 21490 31628 21496
rect 31588 21418 31616 21490
rect 31576 21412 31628 21418
rect 31576 21354 31628 21360
rect 31760 21140 31812 21146
rect 31760 21082 31812 21088
rect 31576 20460 31628 20466
rect 31576 20402 31628 20408
rect 31588 18766 31616 20402
rect 31576 18760 31628 18766
rect 31628 18720 31708 18748
rect 31576 18702 31628 18708
rect 31576 18624 31628 18630
rect 31574 18592 31576 18601
rect 31628 18592 31630 18601
rect 31574 18527 31630 18536
rect 31680 18358 31708 18720
rect 31772 18358 31800 21082
rect 31852 20052 31904 20058
rect 31852 19994 31904 20000
rect 31668 18352 31720 18358
rect 31668 18294 31720 18300
rect 31760 18352 31812 18358
rect 31760 18294 31812 18300
rect 31576 17672 31628 17678
rect 31576 17614 31628 17620
rect 31484 17196 31536 17202
rect 31484 17138 31536 17144
rect 31588 17082 31616 17614
rect 31760 17536 31812 17542
rect 31760 17478 31812 17484
rect 31668 17264 31720 17270
rect 31668 17206 31720 17212
rect 31496 17054 31616 17082
rect 31496 14618 31524 17054
rect 31574 16688 31630 16697
rect 31574 16623 31630 16632
rect 31588 16590 31616 16623
rect 31576 16584 31628 16590
rect 31576 16526 31628 16532
rect 31484 14612 31536 14618
rect 31484 14554 31536 14560
rect 31484 14408 31536 14414
rect 31482 14376 31484 14385
rect 31536 14376 31538 14385
rect 31482 14311 31538 14320
rect 31588 13025 31616 16526
rect 31680 14278 31708 17206
rect 31772 16658 31800 17478
rect 31864 17338 31892 19994
rect 31956 17610 31984 27474
rect 32140 23662 32168 33458
rect 32128 23656 32180 23662
rect 32128 23598 32180 23604
rect 32034 20632 32090 20641
rect 32034 20567 32090 20576
rect 32048 19009 32076 20567
rect 32034 19000 32090 19009
rect 32034 18935 32090 18944
rect 32232 18698 32260 42774
rect 32772 42084 32824 42090
rect 32772 42026 32824 42032
rect 32404 41472 32456 41478
rect 32404 41414 32456 41420
rect 32416 31482 32444 41414
rect 32784 33522 32812 42026
rect 32956 36304 33008 36310
rect 32956 36246 33008 36252
rect 32968 34406 32996 36246
rect 32956 34400 33008 34406
rect 32956 34342 33008 34348
rect 32864 33652 32916 33658
rect 32864 33594 32916 33600
rect 32772 33516 32824 33522
rect 32772 33458 32824 33464
rect 32876 33386 32904 33594
rect 32968 33522 32996 34342
rect 32956 33516 33008 33522
rect 32956 33458 33008 33464
rect 33048 33516 33100 33522
rect 33048 33458 33100 33464
rect 32772 33380 32824 33386
rect 32772 33322 32824 33328
rect 32864 33380 32916 33386
rect 32864 33322 32916 33328
rect 32784 33046 32812 33322
rect 32772 33040 32824 33046
rect 33060 32994 33088 33458
rect 33416 33312 33468 33318
rect 33416 33254 33468 33260
rect 32772 32982 32824 32988
rect 32968 32966 33088 32994
rect 32404 31476 32456 31482
rect 32404 31418 32456 31424
rect 32864 29300 32916 29306
rect 32864 29242 32916 29248
rect 32876 27538 32904 29242
rect 32968 29034 32996 32966
rect 33428 32910 33456 33254
rect 33508 33108 33560 33114
rect 33508 33050 33560 33056
rect 33048 32904 33100 32910
rect 33048 32846 33100 32852
rect 33416 32904 33468 32910
rect 33416 32846 33468 32852
rect 33060 31686 33088 32846
rect 33520 32434 33548 33050
rect 33508 32428 33560 32434
rect 33508 32370 33560 32376
rect 33508 32292 33560 32298
rect 33508 32234 33560 32240
rect 33520 31958 33548 32234
rect 33508 31952 33560 31958
rect 33508 31894 33560 31900
rect 33520 31754 33548 31894
rect 33508 31748 33560 31754
rect 33508 31690 33560 31696
rect 33048 31680 33100 31686
rect 33048 31622 33100 31628
rect 33140 31272 33192 31278
rect 33140 31214 33192 31220
rect 33152 29073 33180 31214
rect 33138 29064 33194 29073
rect 32956 29028 33008 29034
rect 33138 28999 33194 29008
rect 32956 28970 33008 28976
rect 33048 27872 33100 27878
rect 33048 27814 33100 27820
rect 32864 27532 32916 27538
rect 32864 27474 32916 27480
rect 32588 24812 32640 24818
rect 32588 24754 32640 24760
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 32600 24721 32628 24754
rect 32586 24712 32642 24721
rect 32586 24647 32588 24656
rect 32640 24647 32642 24656
rect 32588 24618 32640 24624
rect 32312 24608 32364 24614
rect 32600 24587 32628 24618
rect 32312 24550 32364 24556
rect 32324 24138 32352 24550
rect 32312 24132 32364 24138
rect 32312 24074 32364 24080
rect 32680 24064 32732 24070
rect 32680 24006 32732 24012
rect 32692 23798 32720 24006
rect 32680 23792 32732 23798
rect 32680 23734 32732 23740
rect 32692 23594 32720 23734
rect 32876 23730 32904 24754
rect 33060 24750 33088 27814
rect 33048 24744 33100 24750
rect 33048 24686 33100 24692
rect 32864 23724 32916 23730
rect 32864 23666 32916 23672
rect 32680 23588 32732 23594
rect 32680 23530 32732 23536
rect 33140 22500 33192 22506
rect 33140 22442 33192 22448
rect 33152 22166 33180 22442
rect 33140 22160 33192 22166
rect 33140 22102 33192 22108
rect 33520 22094 33548 31690
rect 33600 31680 33652 31686
rect 33600 31622 33652 31628
rect 33612 31346 33640 31622
rect 33600 31340 33652 31346
rect 33600 31282 33652 31288
rect 33598 22808 33654 22817
rect 33598 22743 33654 22752
rect 33612 22574 33640 22743
rect 33600 22568 33652 22574
rect 33600 22510 33652 22516
rect 33244 22066 33548 22094
rect 32312 21004 32364 21010
rect 32312 20946 32364 20952
rect 32324 20058 32352 20946
rect 32680 20800 32732 20806
rect 32680 20742 32732 20748
rect 32692 20534 32720 20742
rect 32496 20528 32548 20534
rect 32496 20470 32548 20476
rect 32680 20528 32732 20534
rect 32680 20470 32732 20476
rect 32312 20052 32364 20058
rect 32312 19994 32364 20000
rect 32220 18692 32272 18698
rect 32220 18634 32272 18640
rect 32312 18352 32364 18358
rect 32312 18294 32364 18300
rect 32034 17912 32090 17921
rect 32034 17847 32090 17856
rect 32048 17678 32076 17847
rect 32036 17672 32088 17678
rect 32036 17614 32088 17620
rect 32126 17640 32182 17649
rect 31944 17604 31996 17610
rect 32126 17575 32182 17584
rect 31944 17546 31996 17552
rect 31852 17332 31904 17338
rect 31852 17274 31904 17280
rect 31864 16998 31892 17274
rect 31944 17196 31996 17202
rect 31944 17138 31996 17144
rect 31956 17105 31984 17138
rect 32140 17134 32168 17575
rect 32324 17202 32352 18294
rect 32312 17196 32364 17202
rect 32364 17156 32444 17184
rect 32312 17138 32364 17144
rect 32128 17128 32180 17134
rect 31942 17096 31998 17105
rect 32128 17070 32180 17076
rect 31942 17031 31998 17040
rect 31852 16992 31904 16998
rect 31852 16934 31904 16940
rect 32312 16992 32364 16998
rect 32312 16934 32364 16940
rect 32324 16658 32352 16934
rect 31760 16652 31812 16658
rect 31760 16594 31812 16600
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32036 16584 32088 16590
rect 31772 16532 32036 16538
rect 31772 16526 32088 16532
rect 31772 16510 32076 16526
rect 32416 16522 32444 17156
rect 32508 16833 32536 20470
rect 32586 19544 32642 19553
rect 32586 19479 32642 19488
rect 32600 19378 32628 19479
rect 32588 19372 32640 19378
rect 32588 19314 32640 19320
rect 32600 18358 32628 19314
rect 32772 19168 32824 19174
rect 32772 19110 32824 19116
rect 32784 18766 32812 19110
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32864 18760 32916 18766
rect 32864 18702 32916 18708
rect 32588 18352 32640 18358
rect 32588 18294 32640 18300
rect 32680 18148 32732 18154
rect 32680 18090 32732 18096
rect 32692 18057 32720 18090
rect 32772 18080 32824 18086
rect 32678 18048 32734 18057
rect 32876 18057 32904 18702
rect 33138 18456 33194 18465
rect 33138 18391 33194 18400
rect 33152 18290 33180 18391
rect 33140 18284 33192 18290
rect 33140 18226 33192 18232
rect 32772 18022 32824 18028
rect 32862 18048 32918 18057
rect 32678 17983 32734 17992
rect 32784 17814 32812 18022
rect 32862 17983 32918 17992
rect 33138 17912 33194 17921
rect 33048 17876 33100 17882
rect 33138 17847 33194 17856
rect 33048 17818 33100 17824
rect 32772 17808 32824 17814
rect 32772 17750 32824 17756
rect 32864 17672 32916 17678
rect 32864 17614 32916 17620
rect 32588 17604 32640 17610
rect 32588 17546 32640 17552
rect 32494 16824 32550 16833
rect 32494 16759 32550 16768
rect 32404 16516 32456 16522
rect 31772 14346 31800 16510
rect 32404 16458 32456 16464
rect 32508 15314 32536 16759
rect 32600 16250 32628 17546
rect 32772 17536 32824 17542
rect 32772 17478 32824 17484
rect 32784 17202 32812 17478
rect 32772 17196 32824 17202
rect 32772 17138 32824 17144
rect 32588 16244 32640 16250
rect 32588 16186 32640 16192
rect 32772 16108 32824 16114
rect 32772 16050 32824 16056
rect 32508 15286 32628 15314
rect 32404 15156 32456 15162
rect 32404 15098 32456 15104
rect 31760 14340 31812 14346
rect 31760 14282 31812 14288
rect 31668 14272 31720 14278
rect 31668 14214 31720 14220
rect 32312 14068 32364 14074
rect 32312 14010 32364 14016
rect 32324 13977 32352 14010
rect 32310 13968 32366 13977
rect 32128 13932 32180 13938
rect 32416 13938 32444 15098
rect 32496 14816 32548 14822
rect 32496 14758 32548 14764
rect 32508 14414 32536 14758
rect 32496 14408 32548 14414
rect 32496 14350 32548 14356
rect 32600 14260 32628 15286
rect 32508 14232 32628 14260
rect 32310 13903 32366 13912
rect 32404 13932 32456 13938
rect 32128 13874 32180 13880
rect 32404 13874 32456 13880
rect 31668 13796 31720 13802
rect 31668 13738 31720 13744
rect 31574 13016 31630 13025
rect 31574 12951 31630 12960
rect 31484 12708 31536 12714
rect 31484 12650 31536 12656
rect 31496 10441 31524 12650
rect 31680 12646 31708 13738
rect 31852 13728 31904 13734
rect 31852 13670 31904 13676
rect 31864 13326 31892 13670
rect 31852 13320 31904 13326
rect 31852 13262 31904 13268
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31760 13252 31812 13258
rect 31760 13194 31812 13200
rect 31668 12640 31720 12646
rect 31668 12582 31720 12588
rect 31482 10432 31538 10441
rect 31482 10367 31538 10376
rect 31392 9716 31444 9722
rect 31392 9658 31444 9664
rect 31496 9586 31524 10367
rect 31668 10260 31720 10266
rect 31668 10202 31720 10208
rect 31680 10130 31708 10202
rect 31668 10124 31720 10130
rect 31668 10066 31720 10072
rect 31484 9580 31536 9586
rect 31484 9522 31536 9528
rect 31668 9172 31720 9178
rect 31668 9114 31720 9120
rect 31680 8974 31708 9114
rect 31300 8968 31352 8974
rect 31300 8910 31352 8916
rect 31668 8968 31720 8974
rect 31668 8910 31720 8916
rect 31772 8906 31800 13194
rect 31864 9178 31892 13262
rect 31956 12442 31984 13262
rect 31944 12436 31996 12442
rect 31944 12378 31996 12384
rect 32036 9920 32088 9926
rect 32036 9862 32088 9868
rect 32048 9450 32076 9862
rect 32036 9444 32088 9450
rect 32036 9386 32088 9392
rect 31852 9172 31904 9178
rect 31852 9114 31904 9120
rect 32048 8974 32076 9386
rect 32140 8974 32168 13874
rect 32220 13456 32272 13462
rect 32220 13398 32272 13404
rect 32232 13326 32260 13398
rect 32220 13320 32272 13326
rect 32220 13262 32272 13268
rect 32416 12434 32444 13874
rect 32232 12406 32444 12434
rect 32036 8968 32088 8974
rect 32128 8968 32180 8974
rect 32036 8910 32088 8916
rect 32126 8936 32128 8945
rect 32180 8936 32182 8945
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31760 8900 31812 8906
rect 32126 8871 32182 8880
rect 31760 8842 31812 8848
rect 31208 8832 31260 8838
rect 31208 8774 31260 8780
rect 31220 7954 31248 8774
rect 31300 8492 31352 8498
rect 31300 8434 31352 8440
rect 31024 7948 31076 7954
rect 31024 7890 31076 7896
rect 31208 7948 31260 7954
rect 31208 7890 31260 7896
rect 31036 7834 31064 7890
rect 31312 7834 31340 8434
rect 31392 8288 31444 8294
rect 31392 8230 31444 8236
rect 31036 7806 31340 7834
rect 30932 7540 30984 7546
rect 30932 7482 30984 7488
rect 30840 7200 30892 7206
rect 30840 7142 30892 7148
rect 30944 6254 30972 7482
rect 31208 7200 31260 7206
rect 31208 7142 31260 7148
rect 31220 6798 31248 7142
rect 31208 6792 31260 6798
rect 31312 6764 31340 7806
rect 31404 6848 31432 8230
rect 31496 7954 31524 8842
rect 31944 8832 31996 8838
rect 31944 8774 31996 8780
rect 31576 8628 31628 8634
rect 31576 8570 31628 8576
rect 31588 8498 31616 8570
rect 31576 8492 31628 8498
rect 31576 8434 31628 8440
rect 31588 8401 31616 8434
rect 31668 8424 31720 8430
rect 31574 8392 31630 8401
rect 31668 8366 31720 8372
rect 31574 8327 31630 8336
rect 31484 7948 31536 7954
rect 31484 7890 31536 7896
rect 31588 7886 31616 8327
rect 31576 7880 31628 7886
rect 31576 7822 31628 7828
rect 31484 6860 31536 6866
rect 31404 6820 31484 6848
rect 31484 6802 31536 6808
rect 31208 6734 31260 6740
rect 31300 6758 31352 6764
rect 31588 6730 31616 7822
rect 31680 7750 31708 8366
rect 31760 7880 31812 7886
rect 31760 7822 31812 7828
rect 31668 7744 31720 7750
rect 31668 7686 31720 7692
rect 31668 6860 31720 6866
rect 31668 6802 31720 6808
rect 31300 6700 31352 6706
rect 31576 6724 31628 6730
rect 31208 6316 31260 6322
rect 31208 6258 31260 6264
rect 30932 6248 30984 6254
rect 30932 6190 30984 6196
rect 30944 4622 30972 6190
rect 31116 5908 31168 5914
rect 31116 5850 31168 5856
rect 31128 5166 31156 5850
rect 31116 5160 31168 5166
rect 31116 5102 31168 5108
rect 30932 4616 30984 4622
rect 30932 4558 30984 4564
rect 30944 3602 30972 4558
rect 31220 4010 31248 6258
rect 31312 6186 31340 6700
rect 31576 6666 31628 6672
rect 31300 6180 31352 6186
rect 31300 6122 31352 6128
rect 31680 5710 31708 6802
rect 31772 6662 31800 7822
rect 31760 6656 31812 6662
rect 31760 6598 31812 6604
rect 31850 6488 31906 6497
rect 31850 6423 31852 6432
rect 31904 6423 31906 6432
rect 31852 6394 31904 6400
rect 31956 6322 31984 8774
rect 32140 8566 32168 8871
rect 32128 8560 32180 8566
rect 32128 8502 32180 8508
rect 32036 8084 32088 8090
rect 32036 8026 32088 8032
rect 32128 8084 32180 8090
rect 32128 8026 32180 8032
rect 31944 6316 31996 6322
rect 31944 6258 31996 6264
rect 31668 5704 31720 5710
rect 31668 5646 31720 5652
rect 31944 5364 31996 5370
rect 31944 5306 31996 5312
rect 31760 4140 31812 4146
rect 31760 4082 31812 4088
rect 31208 4004 31260 4010
rect 31208 3946 31260 3952
rect 30932 3596 30984 3602
rect 30932 3538 30984 3544
rect 30748 3120 30800 3126
rect 30748 3062 30800 3068
rect 31220 3058 31248 3946
rect 31668 3936 31720 3942
rect 31668 3878 31720 3884
rect 31484 3392 31536 3398
rect 31484 3334 31536 3340
rect 31496 3058 31524 3334
rect 31208 3052 31260 3058
rect 31208 2994 31260 3000
rect 31484 3052 31536 3058
rect 31484 2994 31536 3000
rect 30748 2984 30800 2990
rect 30748 2926 30800 2932
rect 31576 2984 31628 2990
rect 31576 2926 31628 2932
rect 30472 2372 30524 2378
rect 30472 2314 30524 2320
rect 30484 800 30512 2314
rect 30760 800 30788 2926
rect 31208 2508 31260 2514
rect 31208 2450 31260 2456
rect 31024 2372 31076 2378
rect 31024 2314 31076 2320
rect 31036 800 31064 2314
rect 31220 1902 31248 2450
rect 31300 2304 31352 2310
rect 31300 2246 31352 2252
rect 31208 1896 31260 1902
rect 31208 1838 31260 1844
rect 31312 800 31340 2246
rect 31588 800 31616 2926
rect 31680 2038 31708 3878
rect 31772 2854 31800 4082
rect 31956 3534 31984 5306
rect 32048 4214 32076 8026
rect 32140 7954 32168 8026
rect 32128 7948 32180 7954
rect 32128 7890 32180 7896
rect 32128 5704 32180 5710
rect 32128 5646 32180 5652
rect 32140 4690 32168 5646
rect 32128 4684 32180 4690
rect 32128 4626 32180 4632
rect 32036 4208 32088 4214
rect 32036 4150 32088 4156
rect 31944 3528 31996 3534
rect 31944 3470 31996 3476
rect 32048 3466 32076 4150
rect 32036 3460 32088 3466
rect 32036 3402 32088 3408
rect 32232 3398 32260 12406
rect 32404 11076 32456 11082
rect 32404 11018 32456 11024
rect 32416 10538 32444 11018
rect 32404 10532 32456 10538
rect 32404 10474 32456 10480
rect 32312 10464 32364 10470
rect 32312 10406 32364 10412
rect 32324 8498 32352 10406
rect 32404 8900 32456 8906
rect 32404 8842 32456 8848
rect 32416 8566 32444 8842
rect 32404 8560 32456 8566
rect 32404 8502 32456 8508
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 32324 8294 32352 8434
rect 32312 8288 32364 8294
rect 32312 8230 32364 8236
rect 32324 7410 32352 8230
rect 32404 7948 32456 7954
rect 32404 7890 32456 7896
rect 32416 7546 32444 7890
rect 32404 7540 32456 7546
rect 32404 7482 32456 7488
rect 32312 7404 32364 7410
rect 32312 7346 32364 7352
rect 32404 7404 32456 7410
rect 32404 7346 32456 7352
rect 32416 5234 32444 7346
rect 32404 5228 32456 5234
rect 32404 5170 32456 5176
rect 32312 5024 32364 5030
rect 32312 4966 32364 4972
rect 32324 4622 32352 4966
rect 32312 4616 32364 4622
rect 32312 4558 32364 4564
rect 32416 4554 32444 5170
rect 32404 4548 32456 4554
rect 32404 4490 32456 4496
rect 32312 4480 32364 4486
rect 32312 4422 32364 4428
rect 32324 3534 32352 4422
rect 32312 3528 32364 3534
rect 32508 3516 32536 14232
rect 32588 12776 32640 12782
rect 32588 12718 32640 12724
rect 32600 11286 32628 12718
rect 32784 12646 32812 16050
rect 32772 12640 32824 12646
rect 32772 12582 32824 12588
rect 32680 12096 32732 12102
rect 32680 12038 32732 12044
rect 32588 11280 32640 11286
rect 32588 11222 32640 11228
rect 32692 11098 32720 12038
rect 32876 11898 32904 17614
rect 33060 17542 33088 17818
rect 33152 17678 33180 17847
rect 33140 17672 33192 17678
rect 33140 17614 33192 17620
rect 33244 17610 33272 22066
rect 33416 21616 33468 21622
rect 33416 21558 33468 21564
rect 33324 20528 33376 20534
rect 33324 20470 33376 20476
rect 33336 18086 33364 20470
rect 33428 18766 33456 21558
rect 33600 19168 33652 19174
rect 33600 19110 33652 19116
rect 33612 18902 33640 19110
rect 33600 18896 33652 18902
rect 33600 18838 33652 18844
rect 33612 18766 33640 18838
rect 33416 18760 33468 18766
rect 33416 18702 33468 18708
rect 33600 18760 33652 18766
rect 33600 18702 33652 18708
rect 33324 18080 33376 18086
rect 33324 18022 33376 18028
rect 33232 17604 33284 17610
rect 33232 17546 33284 17552
rect 33048 17536 33100 17542
rect 33048 17478 33100 17484
rect 33230 17504 33286 17513
rect 33230 17439 33286 17448
rect 33244 17270 33272 17439
rect 33232 17264 33284 17270
rect 33232 17206 33284 17212
rect 33140 15904 33192 15910
rect 33140 15846 33192 15852
rect 33152 15026 33180 15846
rect 33140 15020 33192 15026
rect 33140 14962 33192 14968
rect 33232 14340 33284 14346
rect 33232 14282 33284 14288
rect 32864 11892 32916 11898
rect 32864 11834 32916 11840
rect 33244 11354 33272 14282
rect 33232 11348 33284 11354
rect 33232 11290 33284 11296
rect 32600 11082 32720 11098
rect 33232 11144 33284 11150
rect 33232 11086 33284 11092
rect 32588 11076 32720 11082
rect 32640 11070 32720 11076
rect 32588 11018 32640 11024
rect 32772 11008 32824 11014
rect 32772 10950 32824 10956
rect 32588 9444 32640 9450
rect 32588 9386 32640 9392
rect 32600 7206 32628 9386
rect 32784 8498 32812 10950
rect 33244 10470 33272 11086
rect 33232 10464 33284 10470
rect 33232 10406 33284 10412
rect 32956 9920 33008 9926
rect 32956 9862 33008 9868
rect 32862 8936 32918 8945
rect 32862 8871 32864 8880
rect 32916 8871 32918 8880
rect 32864 8842 32916 8848
rect 32772 8492 32824 8498
rect 32772 8434 32824 8440
rect 32588 7200 32640 7206
rect 32588 7142 32640 7148
rect 32680 6316 32732 6322
rect 32680 6258 32732 6264
rect 32692 5574 32720 6258
rect 32680 5568 32732 5574
rect 32680 5510 32732 5516
rect 32784 5370 32812 8434
rect 32864 6792 32916 6798
rect 32864 6734 32916 6740
rect 32876 5914 32904 6734
rect 32864 5908 32916 5914
rect 32864 5850 32916 5856
rect 32772 5364 32824 5370
rect 32772 5306 32824 5312
rect 32680 5160 32732 5166
rect 32864 5160 32916 5166
rect 32732 5120 32864 5148
rect 32680 5102 32732 5108
rect 32864 5102 32916 5108
rect 32968 4146 32996 9862
rect 33244 9330 33272 10406
rect 33152 9302 33272 9330
rect 33048 6656 33100 6662
rect 33048 6598 33100 6604
rect 33060 6390 33088 6598
rect 33048 6384 33100 6390
rect 33048 6326 33100 6332
rect 33152 6118 33180 9302
rect 33336 8514 33364 18022
rect 33428 12918 33456 18702
rect 33508 18284 33560 18290
rect 33612 18272 33640 18702
rect 33704 18630 33732 59366
rect 33784 56432 33836 56438
rect 33784 56374 33836 56380
rect 33796 55214 33824 56374
rect 33968 56364 34020 56370
rect 33968 56306 34020 56312
rect 33980 56234 34008 56306
rect 33968 56228 34020 56234
rect 33968 56170 34020 56176
rect 33796 55186 34100 55214
rect 34072 33522 34100 55186
rect 34060 33516 34112 33522
rect 34060 33458 34112 33464
rect 34072 33114 34100 33458
rect 34060 33108 34112 33114
rect 34060 33050 34112 33056
rect 33968 32836 34020 32842
rect 33968 32778 34020 32784
rect 33784 32768 33836 32774
rect 33784 32710 33836 32716
rect 33796 31346 33824 32710
rect 33876 32428 33928 32434
rect 33876 32370 33928 32376
rect 33888 31890 33916 32370
rect 33876 31884 33928 31890
rect 33876 31826 33928 31832
rect 33980 31822 34008 32778
rect 34152 32360 34204 32366
rect 34152 32302 34204 32308
rect 33968 31816 34020 31822
rect 33968 31758 34020 31764
rect 34060 31680 34112 31686
rect 34060 31622 34112 31628
rect 34072 31346 34100 31622
rect 33784 31340 33836 31346
rect 33784 31282 33836 31288
rect 34060 31340 34112 31346
rect 34060 31282 34112 31288
rect 33784 30388 33836 30394
rect 33784 30330 33836 30336
rect 33796 19718 33824 30330
rect 34164 28966 34192 32302
rect 34256 29578 34284 60454
rect 34934 60412 35242 60421
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60347 35242 60356
rect 34934 59324 35242 59333
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59259 35242 59268
rect 34934 58236 35242 58245
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58171 35242 58180
rect 34520 57588 34572 57594
rect 34520 57530 34572 57536
rect 34532 57050 34560 57530
rect 35348 57248 35400 57254
rect 35348 57190 35400 57196
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 34520 57044 34572 57050
rect 34520 56986 34572 56992
rect 34980 57044 35032 57050
rect 34980 56986 35032 56992
rect 34992 56302 35020 56986
rect 35360 56681 35388 57190
rect 35346 56672 35402 56681
rect 35346 56607 35402 56616
rect 34980 56296 35032 56302
rect 34980 56238 35032 56244
rect 35532 56160 35584 56166
rect 35532 56102 35584 56108
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34428 40996 34480 41002
rect 34428 40938 34480 40944
rect 34336 40928 34388 40934
rect 34336 40870 34388 40876
rect 34244 29572 34296 29578
rect 34244 29514 34296 29520
rect 34152 28960 34204 28966
rect 34152 28902 34204 28908
rect 34348 26874 34376 40870
rect 34440 32450 34468 40938
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35440 35828 35492 35834
rect 35440 35770 35492 35776
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35452 34678 35480 35770
rect 35440 34672 35492 34678
rect 35440 34614 35492 34620
rect 34612 34400 34664 34406
rect 34612 34342 34664 34348
rect 34440 32422 34560 32450
rect 34532 31770 34560 32422
rect 34256 26846 34376 26874
rect 34440 31742 34560 31770
rect 33966 23624 34022 23633
rect 33966 23559 34022 23568
rect 33874 23080 33930 23089
rect 33874 23015 33876 23024
rect 33928 23015 33930 23024
rect 33876 22986 33928 22992
rect 33888 21894 33916 22986
rect 33980 22030 34008 23559
rect 34152 22976 34204 22982
rect 34152 22918 34204 22924
rect 34164 22681 34192 22918
rect 34150 22672 34206 22681
rect 34060 22636 34112 22642
rect 34150 22607 34206 22616
rect 34060 22578 34112 22584
rect 33968 22024 34020 22030
rect 33968 21966 34020 21972
rect 33876 21888 33928 21894
rect 33876 21830 33928 21836
rect 33968 21480 34020 21486
rect 33968 21422 34020 21428
rect 33980 20874 34008 21422
rect 33968 20868 34020 20874
rect 33968 20810 34020 20816
rect 33980 20398 34008 20810
rect 33968 20392 34020 20398
rect 33968 20334 34020 20340
rect 33784 19712 33836 19718
rect 33784 19654 33836 19660
rect 33796 19174 33824 19654
rect 33784 19168 33836 19174
rect 33784 19110 33836 19116
rect 33876 18760 33928 18766
rect 33928 18720 34008 18748
rect 33876 18702 33928 18708
rect 33784 18692 33836 18698
rect 33784 18634 33836 18640
rect 33692 18624 33744 18630
rect 33692 18566 33744 18572
rect 33796 18426 33824 18634
rect 33784 18420 33836 18426
rect 33784 18362 33836 18368
rect 33560 18244 33640 18272
rect 33876 18284 33928 18290
rect 33508 18226 33560 18232
rect 33876 18226 33928 18232
rect 33520 17746 33548 18226
rect 33508 17740 33560 17746
rect 33560 17700 33732 17728
rect 33508 17682 33560 17688
rect 33508 17332 33560 17338
rect 33704 17320 33732 17700
rect 33704 17292 33824 17320
rect 33508 17274 33560 17280
rect 33416 12912 33468 12918
rect 33416 12854 33468 12860
rect 33520 12434 33548 17274
rect 33598 17232 33654 17241
rect 33796 17202 33824 17292
rect 33598 17167 33654 17176
rect 33784 17196 33836 17202
rect 33612 17066 33640 17167
rect 33784 17138 33836 17144
rect 33600 17060 33652 17066
rect 33600 17002 33652 17008
rect 33888 14929 33916 18226
rect 33980 18222 34008 18720
rect 33968 18216 34020 18222
rect 33968 18158 34020 18164
rect 33980 17610 34008 18158
rect 33968 17604 34020 17610
rect 33968 17546 34020 17552
rect 33968 17196 34020 17202
rect 33968 17138 34020 17144
rect 33980 17066 34008 17138
rect 33968 17060 34020 17066
rect 33968 17002 34020 17008
rect 34072 16250 34100 22578
rect 34150 22536 34206 22545
rect 34150 22471 34206 22480
rect 34164 22166 34192 22471
rect 34152 22160 34204 22166
rect 34152 22102 34204 22108
rect 34152 21956 34204 21962
rect 34152 21898 34204 21904
rect 34164 20058 34192 21898
rect 34152 20052 34204 20058
rect 34152 19994 34204 20000
rect 33968 16244 34020 16250
rect 33968 16186 34020 16192
rect 34060 16244 34112 16250
rect 34060 16186 34112 16192
rect 33874 14920 33930 14929
rect 33874 14855 33930 14864
rect 33784 14816 33836 14822
rect 33784 14758 33836 14764
rect 33692 13252 33744 13258
rect 33692 13194 33744 13200
rect 33704 12986 33732 13194
rect 33692 12980 33744 12986
rect 33692 12922 33744 12928
rect 33520 12406 33640 12434
rect 33414 11656 33470 11665
rect 33470 11614 33548 11642
rect 33414 11591 33470 11600
rect 33244 8486 33364 8514
rect 33244 7562 33272 8486
rect 33324 8424 33376 8430
rect 33324 8366 33376 8372
rect 33336 7954 33364 8366
rect 33416 8356 33468 8362
rect 33416 8298 33468 8304
rect 33324 7948 33376 7954
rect 33324 7890 33376 7896
rect 33244 7534 33364 7562
rect 33232 7404 33284 7410
rect 33232 7346 33284 7352
rect 33244 6361 33272 7346
rect 33230 6352 33286 6361
rect 33230 6287 33286 6296
rect 33140 6112 33192 6118
rect 33140 6054 33192 6060
rect 33244 6066 33272 6287
rect 33336 6202 33364 7534
rect 33428 7410 33456 8298
rect 33416 7404 33468 7410
rect 33416 7346 33468 7352
rect 33520 6916 33548 11614
rect 33612 7818 33640 12406
rect 33690 11792 33746 11801
rect 33690 11727 33692 11736
rect 33744 11727 33746 11736
rect 33692 11698 33744 11704
rect 33692 11348 33744 11354
rect 33692 11290 33744 11296
rect 33704 9761 33732 11290
rect 33796 11082 33824 14758
rect 33876 12232 33928 12238
rect 33876 12174 33928 12180
rect 33888 11762 33916 12174
rect 33980 11801 34008 16186
rect 34164 14346 34192 19994
rect 34256 18358 34284 26846
rect 34336 23044 34388 23050
rect 34336 22986 34388 22992
rect 34348 21894 34376 22986
rect 34336 21888 34388 21894
rect 34336 21830 34388 21836
rect 34348 21554 34376 21830
rect 34336 21548 34388 21554
rect 34336 21490 34388 21496
rect 34336 19712 34388 19718
rect 34336 19654 34388 19660
rect 34244 18352 34296 18358
rect 34348 18329 34376 19654
rect 34244 18294 34296 18300
rect 34334 18320 34390 18329
rect 34440 18290 34468 31742
rect 34624 26874 34652 34342
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35348 33652 35400 33658
rect 35348 33594 35400 33600
rect 34704 33380 34756 33386
rect 34704 33322 34756 33328
rect 34716 31822 34744 33322
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35360 32842 35388 33594
rect 35348 32836 35400 32842
rect 35348 32778 35400 32784
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 35360 31754 35388 32778
rect 35268 31726 35388 31754
rect 35268 31414 35296 31726
rect 34796 31408 34848 31414
rect 34796 31350 34848 31356
rect 35256 31408 35308 31414
rect 35256 31350 35308 31356
rect 34808 29850 34836 31350
rect 35164 31340 35216 31346
rect 35164 31282 35216 31288
rect 35348 31340 35400 31346
rect 35348 31282 35400 31288
rect 35176 31249 35204 31282
rect 35162 31240 35218 31249
rect 35162 31175 35218 31184
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35360 30938 35388 31282
rect 35348 30932 35400 30938
rect 35348 30874 35400 30880
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34796 29844 34848 29850
rect 34796 29786 34848 29792
rect 34808 29714 35020 29730
rect 34796 29708 35032 29714
rect 34848 29702 34980 29708
rect 34796 29650 34848 29656
rect 34980 29650 35032 29656
rect 34888 29640 34940 29646
rect 34888 29582 34940 29588
rect 34900 29238 34928 29582
rect 35072 29572 35124 29578
rect 35072 29514 35124 29520
rect 35084 29306 35112 29514
rect 35072 29300 35124 29306
rect 35072 29242 35124 29248
rect 34888 29232 34940 29238
rect 34888 29174 34940 29180
rect 35452 28994 35480 34614
rect 35360 28966 35480 28994
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34532 26846 34652 26874
rect 34532 18358 34560 26846
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34796 24200 34848 24206
rect 34796 24142 34848 24148
rect 34704 23724 34756 23730
rect 34704 23666 34756 23672
rect 34612 23044 34664 23050
rect 34612 22986 34664 22992
rect 34624 22522 34652 22986
rect 34716 22778 34744 23666
rect 34808 23526 34836 24142
rect 35070 23624 35126 23633
rect 35070 23559 35072 23568
rect 35124 23559 35126 23568
rect 35072 23530 35124 23536
rect 34796 23520 34848 23526
rect 34796 23462 34848 23468
rect 34704 22772 34756 22778
rect 34704 22714 34756 22720
rect 34624 22494 34744 22522
rect 34612 22432 34664 22438
rect 34612 22374 34664 22380
rect 34624 21690 34652 22374
rect 34612 21684 34664 21690
rect 34612 21626 34664 21632
rect 34716 19514 34744 22494
rect 34704 19508 34756 19514
rect 34704 19450 34756 19456
rect 34716 19378 34744 19450
rect 34808 19378 34836 23462
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35360 22114 35388 28966
rect 35440 23588 35492 23594
rect 35440 23530 35492 23536
rect 35452 23118 35480 23530
rect 35440 23112 35492 23118
rect 35440 23054 35492 23060
rect 35351 22086 35388 22114
rect 35351 22012 35379 22086
rect 35440 22024 35492 22030
rect 35351 21984 35388 22012
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35360 20942 35388 21984
rect 35440 21966 35492 21972
rect 35452 21690 35480 21966
rect 35440 21684 35492 21690
rect 35440 21626 35492 21632
rect 35440 21548 35492 21554
rect 35440 21490 35492 21496
rect 35452 21010 35480 21490
rect 35440 21004 35492 21010
rect 35440 20946 35492 20952
rect 35348 20936 35400 20942
rect 35348 20878 35400 20884
rect 35440 20868 35492 20874
rect 35440 20810 35492 20816
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34888 19848 34940 19854
rect 34888 19790 34940 19796
rect 34704 19372 34756 19378
rect 34704 19314 34756 19320
rect 34796 19372 34848 19378
rect 34796 19314 34848 19320
rect 34702 19272 34758 19281
rect 34702 19207 34758 19216
rect 34716 18970 34744 19207
rect 34704 18964 34756 18970
rect 34704 18906 34756 18912
rect 34520 18352 34572 18358
rect 34520 18294 34572 18300
rect 34334 18255 34390 18264
rect 34428 18284 34480 18290
rect 34704 18284 34756 18290
rect 34428 18226 34480 18232
rect 34624 18244 34704 18272
rect 34518 16960 34574 16969
rect 34518 16895 34574 16904
rect 34428 16720 34480 16726
rect 34428 16662 34480 16668
rect 34244 16040 34296 16046
rect 34244 15982 34296 15988
rect 34256 14822 34284 15982
rect 34334 15600 34390 15609
rect 34334 15535 34390 15544
rect 34244 14816 34296 14822
rect 34244 14758 34296 14764
rect 34152 14340 34204 14346
rect 34152 14282 34204 14288
rect 34164 14006 34192 14282
rect 34152 14000 34204 14006
rect 34152 13942 34204 13948
rect 34244 13864 34296 13870
rect 34244 13806 34296 13812
rect 34152 13728 34204 13734
rect 34152 13670 34204 13676
rect 34164 12850 34192 13670
rect 34256 13530 34284 13806
rect 34244 13524 34296 13530
rect 34244 13466 34296 13472
rect 34152 12844 34204 12850
rect 34152 12786 34204 12792
rect 34152 11892 34204 11898
rect 34152 11834 34204 11840
rect 33966 11792 34022 11801
rect 33876 11756 33928 11762
rect 34164 11762 34192 11834
rect 34348 11830 34376 15535
rect 34440 14550 34468 16662
rect 34532 16250 34560 16895
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 34428 14544 34480 14550
rect 34428 14486 34480 14492
rect 34428 13932 34480 13938
rect 34428 13874 34480 13880
rect 34440 11914 34468 13874
rect 34440 11886 34560 11914
rect 34336 11824 34388 11830
rect 34336 11766 34388 11772
rect 33966 11727 33968 11736
rect 33876 11698 33928 11704
rect 34020 11727 34022 11736
rect 34152 11756 34204 11762
rect 33968 11698 34020 11704
rect 34152 11698 34204 11704
rect 34060 11688 34112 11694
rect 34060 11630 34112 11636
rect 33968 11620 34020 11626
rect 33968 11562 34020 11568
rect 33980 11098 34008 11562
rect 34072 11354 34100 11630
rect 34336 11552 34388 11558
rect 34336 11494 34388 11500
rect 34060 11348 34112 11354
rect 34060 11290 34112 11296
rect 34072 11218 34100 11290
rect 34060 11212 34112 11218
rect 34060 11154 34112 11160
rect 33980 11082 34192 11098
rect 33784 11076 33836 11082
rect 33980 11076 34204 11082
rect 33980 11070 34152 11076
rect 33784 11018 33836 11024
rect 34152 11018 34204 11024
rect 33876 11008 33928 11014
rect 33876 10950 33928 10956
rect 33784 10736 33836 10742
rect 33784 10678 33836 10684
rect 33796 10554 33824 10678
rect 33888 10656 33916 10950
rect 33968 10668 34020 10674
rect 33888 10628 33968 10656
rect 33968 10610 34020 10616
rect 33796 10526 34100 10554
rect 33690 9752 33746 9761
rect 33690 9687 33746 9696
rect 33704 8430 33732 9687
rect 33876 9648 33928 9654
rect 33876 9590 33928 9596
rect 33692 8424 33744 8430
rect 33692 8366 33744 8372
rect 33600 7812 33652 7818
rect 33600 7754 33652 7760
rect 33782 7440 33838 7449
rect 33782 7375 33838 7384
rect 33796 7342 33824 7375
rect 33784 7336 33836 7342
rect 33784 7278 33836 7284
rect 33888 7206 33916 9590
rect 33968 8424 34020 8430
rect 33968 8366 34020 8372
rect 33876 7200 33928 7206
rect 33876 7142 33928 7148
rect 33520 6888 33640 6916
rect 33336 6174 33548 6202
rect 33416 6112 33468 6118
rect 33244 6060 33416 6066
rect 33244 6054 33468 6060
rect 33244 6038 33456 6054
rect 33244 5710 33272 6038
rect 33232 5704 33284 5710
rect 33232 5646 33284 5652
rect 33416 5636 33468 5642
rect 33416 5578 33468 5584
rect 33048 5228 33100 5234
rect 33048 5170 33100 5176
rect 33060 4282 33088 5170
rect 33048 4276 33100 4282
rect 33048 4218 33100 4224
rect 33428 4214 33456 5578
rect 33416 4208 33468 4214
rect 33416 4150 33468 4156
rect 32956 4140 33008 4146
rect 32956 4082 33008 4088
rect 33232 3936 33284 3942
rect 33232 3878 33284 3884
rect 32588 3528 32640 3534
rect 32508 3488 32588 3516
rect 32312 3470 32364 3476
rect 32588 3470 32640 3476
rect 32220 3392 32272 3398
rect 32220 3334 32272 3340
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 32128 2916 32180 2922
rect 32128 2858 32180 2864
rect 31760 2848 31812 2854
rect 31760 2790 31812 2796
rect 31852 2848 31904 2854
rect 31852 2790 31904 2796
rect 31668 2032 31720 2038
rect 31668 1974 31720 1980
rect 31864 800 31892 2790
rect 32140 800 32168 2858
rect 32416 800 32444 3062
rect 32956 2984 33008 2990
rect 32956 2926 33008 2932
rect 32680 2372 32732 2378
rect 32680 2314 32732 2320
rect 32692 800 32720 2314
rect 32968 800 32996 2926
rect 33060 2446 33088 3334
rect 33244 3058 33272 3878
rect 33520 3738 33548 6174
rect 33612 5642 33640 6888
rect 33980 6730 34008 8366
rect 33968 6724 34020 6730
rect 33968 6666 34020 6672
rect 33784 6180 33836 6186
rect 33784 6122 33836 6128
rect 33796 5778 33824 6122
rect 33784 5772 33836 5778
rect 33784 5714 33836 5720
rect 33600 5636 33652 5642
rect 33600 5578 33652 5584
rect 33692 5228 33744 5234
rect 33692 5170 33744 5176
rect 33600 4820 33652 4826
rect 33600 4762 33652 4768
rect 33612 4146 33640 4762
rect 33600 4140 33652 4146
rect 33600 4082 33652 4088
rect 33508 3732 33560 3738
rect 33508 3674 33560 3680
rect 33508 3596 33560 3602
rect 33508 3538 33560 3544
rect 33416 3392 33468 3398
rect 33416 3334 33468 3340
rect 33428 3194 33456 3334
rect 33416 3188 33468 3194
rect 33416 3130 33468 3136
rect 33232 3052 33284 3058
rect 33232 2994 33284 3000
rect 33416 2848 33468 2854
rect 33416 2790 33468 2796
rect 33428 2514 33456 2790
rect 33416 2508 33468 2514
rect 33416 2450 33468 2456
rect 33048 2440 33100 2446
rect 33048 2382 33100 2388
rect 33232 1488 33284 1494
rect 33232 1430 33284 1436
rect 33244 800 33272 1430
rect 33520 800 33548 3538
rect 33704 3398 33732 5170
rect 33796 5166 33824 5714
rect 34072 5370 34100 10526
rect 34348 9586 34376 11494
rect 34532 10826 34560 11886
rect 34624 11830 34652 18244
rect 34704 18226 34756 18232
rect 34704 18080 34756 18086
rect 34704 18022 34756 18028
rect 34716 17202 34744 18022
rect 34704 17196 34756 17202
rect 34704 17138 34756 17144
rect 34704 15972 34756 15978
rect 34704 15914 34756 15920
rect 34716 15638 34744 15914
rect 34704 15632 34756 15638
rect 34704 15574 34756 15580
rect 34808 15570 34836 19314
rect 34900 19242 34928 19790
rect 35348 19372 35400 19378
rect 35348 19314 35400 19320
rect 34888 19236 34940 19242
rect 34888 19178 34940 19184
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18970 35388 19314
rect 35348 18964 35400 18970
rect 35348 18906 35400 18912
rect 34888 18896 34940 18902
rect 34888 18838 34940 18844
rect 34900 18465 34928 18838
rect 35256 18760 35308 18766
rect 35256 18702 35308 18708
rect 35348 18760 35400 18766
rect 35348 18702 35400 18708
rect 34886 18456 34942 18465
rect 34886 18391 34942 18400
rect 34900 18290 34928 18391
rect 34888 18284 34940 18290
rect 34888 18226 34940 18232
rect 35268 18154 35296 18702
rect 35360 18426 35388 18702
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 35348 18284 35400 18290
rect 35348 18226 35400 18232
rect 35256 18148 35308 18154
rect 35256 18090 35308 18096
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17814 35388 18226
rect 35348 17808 35400 17814
rect 35348 17750 35400 17756
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34796 15564 34848 15570
rect 34796 15506 34848 15512
rect 34808 15026 34836 15506
rect 34980 15360 35032 15366
rect 34980 15302 35032 15308
rect 35348 15360 35400 15366
rect 35348 15302 35400 15308
rect 34992 15026 35020 15302
rect 34796 15020 34848 15026
rect 34796 14962 34848 14968
rect 34980 15020 35032 15026
rect 34980 14962 35032 14968
rect 35360 14822 35388 15302
rect 35348 14816 35400 14822
rect 35348 14758 35400 14764
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34612 11824 34664 11830
rect 34612 11766 34664 11772
rect 34702 11792 34758 11801
rect 34702 11727 34758 11736
rect 34612 11620 34664 11626
rect 34612 11562 34664 11568
rect 34624 11286 34652 11562
rect 34612 11280 34664 11286
rect 34612 11222 34664 11228
rect 34612 11076 34664 11082
rect 34612 11018 34664 11024
rect 34440 10798 34560 10826
rect 34336 9580 34388 9586
rect 34336 9522 34388 9528
rect 34440 8922 34468 10798
rect 34520 9512 34572 9518
rect 34520 9454 34572 9460
rect 34348 8894 34468 8922
rect 34150 7984 34206 7993
rect 34150 7919 34152 7928
rect 34204 7919 34206 7928
rect 34152 7890 34204 7896
rect 34164 7410 34192 7890
rect 34152 7404 34204 7410
rect 34152 7346 34204 7352
rect 34060 5364 34112 5370
rect 34060 5306 34112 5312
rect 33784 5160 33836 5166
rect 33784 5102 33836 5108
rect 34348 3942 34376 8894
rect 34428 8832 34480 8838
rect 34428 8774 34480 8780
rect 34440 8498 34468 8774
rect 34428 8492 34480 8498
rect 34428 8434 34480 8440
rect 34532 7342 34560 9454
rect 34624 9194 34652 11018
rect 34716 9674 34744 11727
rect 35360 11665 35388 14758
rect 35452 12102 35480 20810
rect 35440 12096 35492 12102
rect 35440 12038 35492 12044
rect 35346 11656 35402 11665
rect 35346 11591 35402 11600
rect 34796 11552 34848 11558
rect 34796 11494 34848 11500
rect 34808 11218 34836 11494
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34796 11212 34848 11218
rect 34796 11154 34848 11160
rect 34888 11144 34940 11150
rect 34888 11086 34940 11092
rect 34900 10742 34928 11086
rect 34888 10736 34940 10742
rect 34940 10684 35112 10690
rect 34888 10678 35112 10684
rect 34900 10662 35112 10678
rect 34900 10613 34928 10662
rect 35084 10606 35112 10662
rect 35072 10600 35124 10606
rect 35072 10542 35124 10548
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34888 9988 34940 9994
rect 34888 9930 34940 9936
rect 34716 9646 34836 9674
rect 34900 9654 34928 9930
rect 34624 9166 34744 9194
rect 34612 9104 34664 9110
rect 34612 9046 34664 9052
rect 34624 8566 34652 9046
rect 34716 8566 34744 9166
rect 34808 8974 34836 9646
rect 34888 9648 34940 9654
rect 34888 9590 34940 9596
rect 35070 9616 35126 9625
rect 35070 9551 35072 9560
rect 35124 9551 35126 9560
rect 35072 9522 35124 9528
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 34612 8560 34664 8566
rect 34612 8502 34664 8508
rect 34704 8560 34756 8566
rect 34704 8502 34756 8508
rect 34612 7404 34664 7410
rect 34612 7346 34664 7352
rect 34520 7336 34572 7342
rect 34520 7278 34572 7284
rect 34624 7206 34652 7346
rect 34716 7274 34744 8502
rect 34704 7268 34756 7274
rect 34704 7210 34756 7216
rect 34612 7200 34664 7206
rect 34612 7142 34664 7148
rect 34612 6724 34664 6730
rect 34612 6666 34664 6672
rect 34624 5846 34652 6666
rect 34716 6662 34744 7210
rect 34704 6656 34756 6662
rect 34704 6598 34756 6604
rect 34808 6322 34836 8910
rect 34888 8900 34940 8906
rect 34888 8842 34940 8848
rect 34900 8537 34928 8842
rect 34886 8528 34942 8537
rect 34886 8463 34888 8472
rect 34940 8463 34942 8472
rect 34888 8434 34940 8440
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35452 8106 35480 12038
rect 35544 8974 35572 56102
rect 35714 31240 35770 31249
rect 35714 31175 35770 31184
rect 35624 30728 35676 30734
rect 35624 30670 35676 30676
rect 35636 30326 35664 30670
rect 35624 30320 35676 30326
rect 35624 30262 35676 30268
rect 35728 28694 35756 31175
rect 35808 30932 35860 30938
rect 35808 30874 35860 30880
rect 35716 28688 35768 28694
rect 35716 28630 35768 28636
rect 35716 27056 35768 27062
rect 35716 26998 35768 27004
rect 35624 24336 35676 24342
rect 35624 24278 35676 24284
rect 35636 22778 35664 24278
rect 35728 23066 35756 26998
rect 35820 23594 35848 30874
rect 35900 30728 35952 30734
rect 35900 30670 35952 30676
rect 35912 27538 35940 30670
rect 35900 27532 35952 27538
rect 35900 27474 35952 27480
rect 35900 23656 35952 23662
rect 35900 23598 35952 23604
rect 35808 23588 35860 23594
rect 35808 23530 35860 23536
rect 35728 23038 35848 23066
rect 35714 22944 35770 22953
rect 35714 22879 35770 22888
rect 35728 22778 35756 22879
rect 35624 22772 35676 22778
rect 35624 22714 35676 22720
rect 35716 22772 35768 22778
rect 35716 22714 35768 22720
rect 35714 22672 35770 22681
rect 35624 22636 35676 22642
rect 35714 22607 35770 22616
rect 35624 22578 35676 22584
rect 35636 22545 35664 22578
rect 35622 22536 35678 22545
rect 35622 22471 35678 22480
rect 35624 22024 35676 22030
rect 35624 21966 35676 21972
rect 35636 20874 35664 21966
rect 35728 21690 35756 22607
rect 35716 21684 35768 21690
rect 35716 21626 35768 21632
rect 35716 21548 35768 21554
rect 35820 21536 35848 23038
rect 35912 22778 35940 23598
rect 35900 22772 35952 22778
rect 35900 22714 35952 22720
rect 35900 22432 35952 22438
rect 35900 22374 35952 22380
rect 35768 21508 35848 21536
rect 35716 21490 35768 21496
rect 35624 20868 35676 20874
rect 35624 20810 35676 20816
rect 35624 18352 35676 18358
rect 35624 18294 35676 18300
rect 35532 8968 35584 8974
rect 35532 8910 35584 8916
rect 35532 8424 35584 8430
rect 35532 8366 35584 8372
rect 35268 8078 35480 8106
rect 34980 7812 35032 7818
rect 34980 7754 35032 7760
rect 34992 7546 35020 7754
rect 34980 7540 35032 7546
rect 34980 7482 35032 7488
rect 35164 7540 35216 7546
rect 35164 7482 35216 7488
rect 35176 7274 35204 7482
rect 35164 7268 35216 7274
rect 35164 7210 35216 7216
rect 35268 7206 35296 8078
rect 35348 7948 35400 7954
rect 35348 7890 35400 7896
rect 35256 7200 35308 7206
rect 35256 7142 35308 7148
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34796 6316 34848 6322
rect 34796 6258 34848 6264
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34612 5840 34664 5846
rect 34612 5782 34664 5788
rect 34520 5772 34572 5778
rect 34520 5714 34572 5720
rect 34532 5574 34560 5714
rect 34520 5568 34572 5574
rect 34520 5510 34572 5516
rect 34624 5234 34652 5782
rect 35360 5778 35388 7890
rect 35440 7404 35492 7410
rect 35440 7346 35492 7352
rect 35452 6866 35480 7346
rect 35544 7342 35572 8366
rect 35532 7336 35584 7342
rect 35532 7278 35584 7284
rect 35532 7200 35584 7206
rect 35532 7142 35584 7148
rect 35440 6860 35492 6866
rect 35440 6802 35492 6808
rect 35544 6746 35572 7142
rect 35636 6798 35664 18294
rect 35728 11898 35756 21490
rect 35912 21434 35940 22374
rect 35820 21406 35940 21434
rect 35820 21078 35848 21406
rect 35808 21072 35860 21078
rect 35808 21014 35860 21020
rect 35900 20256 35952 20262
rect 35900 20198 35952 20204
rect 35912 18970 35940 20198
rect 35900 18964 35952 18970
rect 35900 18906 35952 18912
rect 35808 18420 35860 18426
rect 35808 18362 35860 18368
rect 35820 15434 35848 18362
rect 35900 17264 35952 17270
rect 35900 17206 35952 17212
rect 35808 15428 35860 15434
rect 35808 15370 35860 15376
rect 35912 15314 35940 17206
rect 35820 15286 35940 15314
rect 35716 11892 35768 11898
rect 35716 11834 35768 11840
rect 35716 9580 35768 9586
rect 35716 9522 35768 9528
rect 35452 6718 35572 6746
rect 35624 6792 35676 6798
rect 35624 6734 35676 6740
rect 35348 5772 35400 5778
rect 35348 5714 35400 5720
rect 34796 5568 34848 5574
rect 34796 5510 34848 5516
rect 34704 5364 34756 5370
rect 34704 5306 34756 5312
rect 34612 5228 34664 5234
rect 34612 5170 34664 5176
rect 34428 4616 34480 4622
rect 34428 4558 34480 4564
rect 34336 3936 34388 3942
rect 34336 3878 34388 3884
rect 34440 3738 34468 4558
rect 34612 4548 34664 4554
rect 34612 4490 34664 4496
rect 34428 3732 34480 3738
rect 34428 3674 34480 3680
rect 34520 3528 34572 3534
rect 34520 3470 34572 3476
rect 33968 3460 34020 3466
rect 33968 3402 34020 3408
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 33600 2848 33652 2854
rect 33600 2790 33652 2796
rect 33612 1494 33640 2790
rect 33600 1488 33652 1494
rect 33600 1430 33652 1436
rect 33796 800 33824 3130
rect 33980 3058 34008 3402
rect 34532 3058 34560 3470
rect 33968 3052 34020 3058
rect 33968 2994 34020 3000
rect 34520 3052 34572 3058
rect 34520 2994 34572 3000
rect 34336 2304 34388 2310
rect 34336 2246 34388 2252
rect 34060 1420 34112 1426
rect 34060 1362 34112 1368
rect 34072 800 34100 1362
rect 34348 800 34376 2246
rect 34624 800 34652 4490
rect 34716 3534 34744 5306
rect 34808 4622 34836 5510
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34796 4616 34848 4622
rect 34796 4558 34848 4564
rect 35452 4026 35480 6718
rect 35624 6384 35676 6390
rect 35624 6326 35676 6332
rect 35532 5636 35584 5642
rect 35532 5578 35584 5584
rect 35544 5302 35572 5578
rect 35532 5296 35584 5302
rect 35532 5238 35584 5244
rect 35636 4146 35664 6326
rect 35728 4146 35756 9522
rect 35820 6390 35848 15286
rect 35900 11076 35952 11082
rect 35900 11018 35952 11024
rect 35912 10674 35940 11018
rect 36004 10742 36032 60998
rect 36372 60790 36400 63294
rect 36910 63294 37228 63322
rect 36910 63200 36966 63294
rect 37200 61180 37228 63294
rect 37646 63200 37702 64000
rect 38382 63200 38438 64000
rect 39118 63322 39174 64000
rect 39118 63294 39528 63322
rect 39118 63200 39174 63294
rect 37660 61198 37688 63200
rect 38396 61198 38424 63200
rect 37280 61192 37332 61198
rect 37200 61152 37280 61180
rect 37280 61134 37332 61140
rect 37648 61192 37700 61198
rect 37648 61134 37700 61140
rect 38384 61192 38436 61198
rect 38384 61134 38436 61140
rect 39500 61130 39528 63294
rect 39854 63200 39910 64000
rect 40590 63322 40646 64000
rect 40590 63294 41000 63322
rect 40590 63200 40646 63294
rect 39868 61180 39896 63200
rect 40972 61198 41000 63294
rect 41326 63200 41382 64000
rect 42062 63200 42118 64000
rect 42798 63200 42854 64000
rect 43534 63322 43590 64000
rect 44270 63322 44326 64000
rect 45006 63322 45062 64000
rect 45742 63322 45798 64000
rect 46478 63322 46534 64000
rect 43534 63294 44128 63322
rect 43534 63200 43590 63294
rect 40040 61192 40092 61198
rect 39868 61152 40040 61180
rect 40040 61134 40092 61140
rect 40960 61192 41012 61198
rect 40960 61134 41012 61140
rect 37740 61124 37792 61130
rect 37740 61066 37792 61072
rect 39488 61124 39540 61130
rect 39488 61066 39540 61072
rect 37280 61056 37332 61062
rect 37280 60998 37332 61004
rect 36360 60784 36412 60790
rect 36360 60726 36412 60732
rect 36452 60512 36504 60518
rect 36452 60454 36504 60460
rect 36084 57452 36136 57458
rect 36084 57394 36136 57400
rect 36360 57452 36412 57458
rect 36360 57394 36412 57400
rect 36096 57050 36124 57394
rect 36372 57254 36400 57394
rect 36360 57248 36412 57254
rect 36360 57190 36412 57196
rect 36084 57044 36136 57050
rect 36084 56986 36136 56992
rect 36372 35766 36400 57190
rect 36464 37262 36492 60454
rect 37292 57934 37320 60998
rect 37280 57928 37332 57934
rect 37280 57870 37332 57876
rect 37752 57526 37780 61066
rect 39764 61056 39816 61062
rect 39764 60998 39816 61004
rect 40224 61056 40276 61062
rect 40224 60998 40276 61004
rect 40960 61056 41012 61062
rect 40960 60998 41012 61004
rect 41052 61056 41104 61062
rect 41052 60998 41104 61004
rect 39776 58546 39804 60998
rect 40132 59016 40184 59022
rect 40132 58958 40184 58964
rect 39672 58540 39724 58546
rect 39672 58482 39724 58488
rect 39764 58540 39816 58546
rect 39764 58482 39816 58488
rect 38660 57928 38712 57934
rect 38660 57870 38712 57876
rect 38476 57860 38528 57866
rect 38476 57802 38528 57808
rect 37740 57520 37792 57526
rect 37740 57462 37792 57468
rect 36636 57452 36688 57458
rect 36636 57394 36688 57400
rect 38108 57452 38160 57458
rect 38108 57394 38160 57400
rect 38200 57452 38252 57458
rect 38200 57394 38252 57400
rect 36648 57050 36676 57394
rect 38120 57361 38148 57394
rect 38106 57352 38162 57361
rect 38016 57316 38068 57322
rect 38106 57287 38162 57296
rect 38016 57258 38068 57264
rect 38028 57202 38056 57258
rect 38212 57202 38240 57394
rect 38028 57174 38240 57202
rect 36636 57044 36688 57050
rect 36636 56986 36688 56992
rect 37924 39296 37976 39302
rect 37924 39238 37976 39244
rect 36452 37256 36504 37262
rect 36452 37198 36504 37204
rect 36544 36712 36596 36718
rect 36544 36654 36596 36660
rect 36360 35760 36412 35766
rect 36360 35702 36412 35708
rect 36556 35222 36584 36654
rect 36544 35216 36596 35222
rect 36544 35158 36596 35164
rect 36084 33516 36136 33522
rect 36084 33458 36136 33464
rect 36096 30734 36124 33458
rect 36544 32768 36596 32774
rect 36544 32710 36596 32716
rect 36556 32570 36584 32710
rect 36544 32564 36596 32570
rect 36544 32506 36596 32512
rect 37004 32292 37056 32298
rect 37004 32234 37056 32240
rect 36176 31952 36228 31958
rect 36176 31894 36228 31900
rect 36084 30728 36136 30734
rect 36084 30670 36136 30676
rect 36188 29646 36216 31894
rect 37016 31754 37044 32234
rect 37016 31726 37136 31754
rect 36268 31272 36320 31278
rect 36268 31214 36320 31220
rect 36280 30734 36308 31214
rect 36268 30728 36320 30734
rect 36268 30670 36320 30676
rect 36912 30728 36964 30734
rect 36912 30670 36964 30676
rect 37004 30728 37056 30734
rect 37004 30670 37056 30676
rect 36280 30394 36308 30670
rect 36924 30394 36952 30670
rect 36268 30388 36320 30394
rect 36268 30330 36320 30336
rect 36912 30388 36964 30394
rect 36912 30330 36964 30336
rect 36820 29844 36872 29850
rect 36820 29786 36872 29792
rect 36176 29640 36228 29646
rect 36176 29582 36228 29588
rect 36636 25424 36688 25430
rect 36636 25366 36688 25372
rect 36084 24812 36136 24818
rect 36084 24754 36136 24760
rect 36096 22642 36124 24754
rect 36176 23860 36228 23866
rect 36176 23802 36228 23808
rect 36188 23186 36216 23802
rect 36452 23724 36504 23730
rect 36452 23666 36504 23672
rect 36176 23180 36228 23186
rect 36176 23122 36228 23128
rect 36464 23089 36492 23666
rect 36544 23112 36596 23118
rect 36450 23080 36506 23089
rect 36268 23044 36320 23050
rect 36544 23054 36596 23060
rect 36450 23015 36506 23024
rect 36268 22986 36320 22992
rect 36176 22976 36228 22982
rect 36176 22918 36228 22924
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 36096 21554 36124 22578
rect 36188 22438 36216 22918
rect 36280 22778 36308 22986
rect 36450 22808 36506 22817
rect 36268 22772 36320 22778
rect 36450 22743 36506 22752
rect 36268 22714 36320 22720
rect 36268 22636 36320 22642
rect 36268 22578 36320 22584
rect 36176 22432 36228 22438
rect 36176 22374 36228 22380
rect 36280 21672 36308 22578
rect 36464 22438 36492 22743
rect 36452 22432 36504 22438
rect 36452 22374 36504 22380
rect 36556 22098 36584 23054
rect 36648 22778 36676 25366
rect 36728 23520 36780 23526
rect 36728 23462 36780 23468
rect 36740 22778 36768 23462
rect 36636 22772 36688 22778
rect 36636 22714 36688 22720
rect 36728 22772 36780 22778
rect 36728 22714 36780 22720
rect 36544 22092 36596 22098
rect 36544 22034 36596 22040
rect 36544 21956 36596 21962
rect 36544 21898 36596 21904
rect 36188 21644 36308 21672
rect 36452 21684 36504 21690
rect 36084 21548 36136 21554
rect 36084 21490 36136 21496
rect 36084 21004 36136 21010
rect 36084 20946 36136 20952
rect 36096 19310 36124 20946
rect 36084 19304 36136 19310
rect 36084 19246 36136 19252
rect 36096 18902 36124 19246
rect 36084 18896 36136 18902
rect 36084 18838 36136 18844
rect 36084 18760 36136 18766
rect 36084 18702 36136 18708
rect 36096 18222 36124 18702
rect 36084 18216 36136 18222
rect 36084 18158 36136 18164
rect 36188 16590 36216 21644
rect 36452 21626 36504 21632
rect 36268 21548 36320 21554
rect 36268 21490 36320 21496
rect 36280 21146 36308 21490
rect 36268 21140 36320 21146
rect 36268 21082 36320 21088
rect 36360 21140 36412 21146
rect 36360 21082 36412 21088
rect 36280 20942 36308 21082
rect 36268 20936 36320 20942
rect 36268 20878 36320 20884
rect 36268 20800 36320 20806
rect 36268 20742 36320 20748
rect 36280 18698 36308 20742
rect 36268 18692 36320 18698
rect 36268 18634 36320 18640
rect 36372 18601 36400 21082
rect 36464 20942 36492 21626
rect 36452 20936 36504 20942
rect 36452 20878 36504 20884
rect 36358 18592 36414 18601
rect 36358 18527 36414 18536
rect 36360 18080 36412 18086
rect 36360 18022 36412 18028
rect 36176 16584 36228 16590
rect 36372 16561 36400 18022
rect 36176 16526 36228 16532
rect 36358 16552 36414 16561
rect 36358 16487 36414 16496
rect 36268 16448 36320 16454
rect 36268 16390 36320 16396
rect 36280 16114 36308 16390
rect 36268 16108 36320 16114
rect 36268 16050 36320 16056
rect 36372 15688 36400 16487
rect 36188 15660 36400 15688
rect 36084 11756 36136 11762
rect 36084 11698 36136 11704
rect 35992 10736 36044 10742
rect 35992 10678 36044 10684
rect 36096 10674 36124 11698
rect 35900 10668 35952 10674
rect 35900 10610 35952 10616
rect 36084 10668 36136 10674
rect 36084 10610 36136 10616
rect 35912 10062 35940 10610
rect 35900 10056 35952 10062
rect 35900 9998 35952 10004
rect 36084 7948 36136 7954
rect 36084 7890 36136 7896
rect 36096 7546 36124 7890
rect 36084 7540 36136 7546
rect 36084 7482 36136 7488
rect 35900 7404 35952 7410
rect 35900 7346 35952 7352
rect 35912 6934 35940 7346
rect 35900 6928 35952 6934
rect 35900 6870 35952 6876
rect 35808 6384 35860 6390
rect 35808 6326 35860 6332
rect 35912 5794 35940 6870
rect 36188 6866 36216 15660
rect 36464 11014 36492 20878
rect 36556 20398 36584 21898
rect 36544 20392 36596 20398
rect 36544 20334 36596 20340
rect 36636 20256 36688 20262
rect 36636 20198 36688 20204
rect 36542 19272 36598 19281
rect 36542 19207 36598 19216
rect 36556 19174 36584 19207
rect 36544 19168 36596 19174
rect 36544 19110 36596 19116
rect 36544 18760 36596 18766
rect 36544 18702 36596 18708
rect 36556 17678 36584 18702
rect 36544 17672 36596 17678
rect 36544 17614 36596 17620
rect 36544 12912 36596 12918
rect 36544 12854 36596 12860
rect 36556 11218 36584 12854
rect 36544 11212 36596 11218
rect 36544 11154 36596 11160
rect 36648 11150 36676 20198
rect 36832 17134 36860 29786
rect 37016 28626 37044 30670
rect 37004 28620 37056 28626
rect 37004 28562 37056 28568
rect 37004 24812 37056 24818
rect 37004 24754 37056 24760
rect 37016 23050 37044 24754
rect 37004 23044 37056 23050
rect 37004 22986 37056 22992
rect 36912 22636 36964 22642
rect 36912 22578 36964 22584
rect 36924 21486 36952 22578
rect 37016 21622 37044 22986
rect 37108 22166 37136 31726
rect 37464 31272 37516 31278
rect 37464 31214 37516 31220
rect 37280 31136 37332 31142
rect 37280 31078 37332 31084
rect 37292 30734 37320 31078
rect 37476 30734 37504 31214
rect 37280 30728 37332 30734
rect 37280 30670 37332 30676
rect 37464 30728 37516 30734
rect 37464 30670 37516 30676
rect 37556 30592 37608 30598
rect 37556 30534 37608 30540
rect 37568 30326 37596 30534
rect 37556 30320 37608 30326
rect 37556 30262 37608 30268
rect 37648 30048 37700 30054
rect 37648 29990 37700 29996
rect 37280 29232 37332 29238
rect 37280 29174 37332 29180
rect 37292 27130 37320 29174
rect 37280 27124 37332 27130
rect 37280 27066 37332 27072
rect 37554 23624 37610 23633
rect 37554 23559 37610 23568
rect 37280 23044 37332 23050
rect 37280 22986 37332 22992
rect 37188 22568 37240 22574
rect 37188 22510 37240 22516
rect 37096 22160 37148 22166
rect 37096 22102 37148 22108
rect 37004 21616 37056 21622
rect 37004 21558 37056 21564
rect 36912 21480 36964 21486
rect 36912 21422 36964 21428
rect 36924 20942 36952 21422
rect 37004 21344 37056 21350
rect 37004 21286 37056 21292
rect 36912 20936 36964 20942
rect 36912 20878 36964 20884
rect 36924 20534 36952 20878
rect 37016 20874 37044 21286
rect 37004 20868 37056 20874
rect 37004 20810 37056 20816
rect 36912 20528 36964 20534
rect 36912 20470 36964 20476
rect 37002 18728 37058 18737
rect 37002 18663 37058 18672
rect 37016 17134 37044 18663
rect 36820 17128 36872 17134
rect 36820 17070 36872 17076
rect 37004 17128 37056 17134
rect 37004 17070 37056 17076
rect 36728 16652 36780 16658
rect 36728 16594 36780 16600
rect 36740 15638 36768 16594
rect 36820 16448 36872 16454
rect 36820 16390 36872 16396
rect 36832 15910 36860 16390
rect 36820 15904 36872 15910
rect 36820 15846 36872 15852
rect 36728 15632 36780 15638
rect 36728 15574 36780 15580
rect 36728 14612 36780 14618
rect 36728 14554 36780 14560
rect 36636 11144 36688 11150
rect 36636 11086 36688 11092
rect 36452 11008 36504 11014
rect 36452 10950 36504 10956
rect 36268 10464 36320 10470
rect 36268 10406 36320 10412
rect 36280 9042 36308 10406
rect 36360 10056 36412 10062
rect 36360 9998 36412 10004
rect 36268 9036 36320 9042
rect 36268 8978 36320 8984
rect 36372 8922 36400 9998
rect 36636 9444 36688 9450
rect 36636 9386 36688 9392
rect 36452 9104 36504 9110
rect 36452 9046 36504 9052
rect 36280 8894 36400 8922
rect 36176 6860 36228 6866
rect 36176 6802 36228 6808
rect 35912 5766 36032 5794
rect 35900 5636 35952 5642
rect 35900 5578 35952 5584
rect 35808 4480 35860 4486
rect 35808 4422 35860 4428
rect 35624 4140 35676 4146
rect 35624 4082 35676 4088
rect 35716 4140 35768 4146
rect 35716 4082 35768 4088
rect 35452 3998 35756 4026
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34796 3460 34848 3466
rect 34796 3402 34848 3408
rect 34704 3392 34756 3398
rect 34704 3334 34756 3340
rect 34716 1714 34744 3334
rect 34808 2446 34836 3402
rect 35624 2984 35676 2990
rect 35624 2926 35676 2932
rect 35348 2916 35400 2922
rect 35348 2858 35400 2864
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 34716 1686 34928 1714
rect 34900 800 34928 1686
rect 35360 1578 35388 2858
rect 35440 2372 35492 2378
rect 35440 2314 35492 2320
rect 35176 1550 35388 1578
rect 35176 800 35204 1550
rect 35452 800 35480 2314
rect 35636 1714 35664 2926
rect 35728 2446 35756 3998
rect 35820 3058 35848 4422
rect 35912 3534 35940 5578
rect 36004 5234 36032 5766
rect 35992 5228 36044 5234
rect 35992 5170 36044 5176
rect 36188 4622 36216 6802
rect 36176 4616 36228 4622
rect 36176 4558 36228 4564
rect 36084 4480 36136 4486
rect 36084 4422 36136 4428
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 35808 3052 35860 3058
rect 35808 2994 35860 3000
rect 36004 2938 36032 3538
rect 35912 2910 36032 2938
rect 35716 2440 35768 2446
rect 35716 2382 35768 2388
rect 35636 1686 35756 1714
rect 35728 800 35756 1686
rect 35912 1426 35940 2910
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 2514 36032 2790
rect 35992 2508 36044 2514
rect 35992 2450 36044 2456
rect 36096 2258 36124 4422
rect 36280 4146 36308 8894
rect 36464 7449 36492 9046
rect 36648 8090 36676 9386
rect 36636 8084 36688 8090
rect 36636 8026 36688 8032
rect 36450 7440 36506 7449
rect 36450 7375 36506 7384
rect 36544 6656 36596 6662
rect 36544 6598 36596 6604
rect 36556 5234 36584 6598
rect 36740 5794 36768 14554
rect 36832 10538 36860 15846
rect 37108 13938 37136 22102
rect 37200 22098 37228 22510
rect 37188 22092 37240 22098
rect 37188 22034 37240 22040
rect 37200 20618 37228 22034
rect 37292 21962 37320 22986
rect 37568 22710 37596 23559
rect 37556 22704 37608 22710
rect 37556 22646 37608 22652
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37476 22030 37504 22578
rect 37464 22024 37516 22030
rect 37464 21966 37516 21972
rect 37280 21956 37332 21962
rect 37280 21898 37332 21904
rect 37372 21548 37424 21554
rect 37372 21490 37424 21496
rect 37200 20590 37320 20618
rect 37188 20392 37240 20398
rect 37188 20334 37240 20340
rect 37200 19334 37228 20334
rect 37292 19854 37320 20590
rect 37280 19848 37332 19854
rect 37280 19790 37332 19796
rect 37384 19446 37412 21490
rect 37660 21486 37688 29990
rect 37832 23656 37884 23662
rect 37832 23598 37884 23604
rect 37844 23254 37872 23598
rect 37832 23248 37884 23254
rect 37832 23190 37884 23196
rect 37832 23112 37884 23118
rect 37832 23054 37884 23060
rect 37844 22778 37872 23054
rect 37832 22772 37884 22778
rect 37832 22714 37884 22720
rect 37936 22094 37964 39238
rect 38488 31754 38516 57802
rect 38672 57594 38700 57870
rect 39684 57866 39712 58482
rect 40040 58336 40092 58342
rect 40040 58278 40092 58284
rect 38936 57860 38988 57866
rect 38936 57802 38988 57808
rect 39672 57860 39724 57866
rect 39672 57802 39724 57808
rect 38844 57792 38896 57798
rect 38844 57734 38896 57740
rect 38856 57594 38884 57734
rect 38660 57588 38712 57594
rect 38660 57530 38712 57536
rect 38844 57588 38896 57594
rect 38844 57530 38896 57536
rect 38568 57452 38620 57458
rect 38568 57394 38620 57400
rect 38580 56846 38608 57394
rect 38568 56840 38620 56846
rect 38568 56782 38620 56788
rect 38948 36922 38976 57802
rect 39396 55888 39448 55894
rect 39396 55830 39448 55836
rect 39304 48680 39356 48686
rect 39304 48622 39356 48628
rect 38936 36916 38988 36922
rect 38936 36858 38988 36864
rect 38948 35834 38976 36858
rect 38936 35828 38988 35834
rect 38936 35770 38988 35776
rect 38660 32020 38712 32026
rect 38660 31962 38712 31968
rect 38476 31748 38528 31754
rect 38476 31690 38528 31696
rect 38672 30734 38700 31962
rect 38660 30728 38712 30734
rect 38660 30670 38712 30676
rect 38384 23724 38436 23730
rect 38384 23666 38436 23672
rect 39120 23724 39172 23730
rect 39120 23666 39172 23672
rect 38396 23322 38424 23666
rect 38752 23656 38804 23662
rect 38752 23598 38804 23604
rect 38936 23656 38988 23662
rect 38936 23598 38988 23604
rect 38384 23316 38436 23322
rect 38384 23258 38436 23264
rect 38108 23248 38160 23254
rect 38108 23190 38160 23196
rect 37844 22066 37964 22094
rect 37648 21480 37700 21486
rect 37648 21422 37700 21428
rect 37464 21344 37516 21350
rect 37464 21286 37516 21292
rect 37476 21078 37504 21286
rect 37464 21072 37516 21078
rect 37464 21014 37516 21020
rect 37556 20868 37608 20874
rect 37556 20810 37608 20816
rect 37648 20868 37700 20874
rect 37648 20810 37700 20816
rect 37464 20460 37516 20466
rect 37464 20402 37516 20408
rect 37372 19440 37424 19446
rect 37372 19382 37424 19388
rect 37200 19306 37320 19334
rect 37292 19258 37320 19306
rect 37292 19230 37412 19258
rect 37096 13932 37148 13938
rect 37096 13874 37148 13880
rect 37188 12912 37240 12918
rect 37188 12854 37240 12860
rect 37200 12102 37228 12854
rect 37188 12096 37240 12102
rect 37188 12038 37240 12044
rect 37004 11212 37056 11218
rect 37004 11154 37056 11160
rect 36820 10532 36872 10538
rect 36820 10474 36872 10480
rect 36912 7744 36964 7750
rect 36912 7686 36964 7692
rect 36924 7546 36952 7686
rect 36912 7540 36964 7546
rect 36912 7482 36964 7488
rect 37016 6662 37044 11154
rect 37280 9376 37332 9382
rect 37280 9318 37332 9324
rect 37292 9178 37320 9318
rect 37280 9172 37332 9178
rect 37280 9114 37332 9120
rect 37280 8968 37332 8974
rect 37280 8910 37332 8916
rect 37096 8900 37148 8906
rect 37096 8842 37148 8848
rect 36820 6656 36872 6662
rect 36820 6598 36872 6604
rect 37004 6656 37056 6662
rect 37004 6598 37056 6604
rect 36832 5914 36860 6598
rect 36820 5908 36872 5914
rect 36820 5850 36872 5856
rect 36740 5766 36860 5794
rect 36728 5636 36780 5642
rect 36728 5578 36780 5584
rect 36740 5370 36768 5578
rect 36832 5370 36860 5766
rect 36728 5364 36780 5370
rect 36728 5306 36780 5312
rect 36820 5364 36872 5370
rect 36820 5306 36872 5312
rect 36544 5228 36596 5234
rect 36544 5170 36596 5176
rect 37016 5166 37044 6598
rect 37108 5166 37136 8842
rect 37292 8401 37320 8910
rect 37278 8392 37334 8401
rect 37278 8327 37334 8336
rect 37292 8022 37320 8327
rect 37280 8016 37332 8022
rect 37280 7958 37332 7964
rect 37384 7886 37412 19230
rect 37476 18970 37504 20402
rect 37568 19922 37596 20810
rect 37660 20602 37688 20810
rect 37648 20596 37700 20602
rect 37648 20538 37700 20544
rect 37556 19916 37608 19922
rect 37556 19858 37608 19864
rect 37648 19848 37700 19854
rect 37648 19790 37700 19796
rect 37740 19848 37792 19854
rect 37740 19790 37792 19796
rect 37660 19446 37688 19790
rect 37752 19514 37780 19790
rect 37740 19508 37792 19514
rect 37740 19450 37792 19456
rect 37556 19440 37608 19446
rect 37556 19382 37608 19388
rect 37648 19440 37700 19446
rect 37844 19394 37872 22066
rect 38120 22030 38148 23190
rect 38108 22024 38160 22030
rect 38764 22012 38792 23598
rect 38842 23080 38898 23089
rect 38842 23015 38844 23024
rect 38896 23015 38898 23024
rect 38844 22986 38896 22992
rect 38948 22710 38976 23598
rect 39028 23520 39080 23526
rect 39028 23462 39080 23468
rect 38936 22704 38988 22710
rect 38936 22646 38988 22652
rect 38948 22574 38976 22646
rect 39040 22642 39068 23462
rect 39028 22636 39080 22642
rect 39028 22578 39080 22584
rect 38936 22568 38988 22574
rect 38936 22510 38988 22516
rect 39132 22098 39160 23666
rect 39120 22092 39172 22098
rect 39120 22034 39172 22040
rect 38844 22024 38896 22030
rect 38764 21984 38844 22012
rect 38108 21966 38160 21972
rect 38844 21966 38896 21972
rect 38856 21622 38884 21966
rect 38844 21616 38896 21622
rect 38672 21576 38844 21604
rect 38292 21412 38344 21418
rect 38292 21354 38344 21360
rect 38200 20936 38252 20942
rect 38200 20878 38252 20884
rect 37924 20800 37976 20806
rect 37924 20742 37976 20748
rect 37648 19382 37700 19388
rect 37568 18970 37596 19382
rect 37464 18964 37516 18970
rect 37464 18906 37516 18912
rect 37556 18964 37608 18970
rect 37556 18906 37608 18912
rect 37660 18766 37688 19382
rect 37752 19378 37872 19394
rect 37936 19378 37964 20742
rect 38016 20256 38068 20262
rect 38016 20198 38068 20204
rect 38108 20256 38160 20262
rect 38108 20198 38160 20204
rect 38028 19854 38056 20198
rect 38016 19848 38068 19854
rect 38016 19790 38068 19796
rect 38120 19666 38148 20198
rect 38028 19638 38148 19666
rect 37740 19372 37872 19378
rect 37792 19366 37872 19372
rect 37740 19314 37792 19320
rect 37740 18896 37792 18902
rect 37740 18838 37792 18844
rect 37648 18760 37700 18766
rect 37648 18702 37700 18708
rect 37752 18426 37780 18838
rect 37740 18420 37792 18426
rect 37740 18362 37792 18368
rect 37844 17678 37872 19366
rect 37924 19372 37976 19378
rect 37924 19314 37976 19320
rect 38028 19310 38056 19638
rect 38016 19304 38068 19310
rect 38016 19246 38068 19252
rect 38028 18834 38056 19246
rect 38016 18828 38068 18834
rect 38016 18770 38068 18776
rect 38108 18284 38160 18290
rect 38108 18226 38160 18232
rect 38120 18193 38148 18226
rect 38106 18184 38162 18193
rect 38106 18119 38162 18128
rect 38212 17785 38240 20878
rect 38198 17776 38254 17785
rect 37924 17740 37976 17746
rect 38198 17711 38254 17720
rect 37924 17682 37976 17688
rect 37832 17672 37884 17678
rect 37832 17614 37884 17620
rect 37740 17604 37792 17610
rect 37740 17546 37792 17552
rect 37752 16794 37780 17546
rect 37740 16788 37792 16794
rect 37740 16730 37792 16736
rect 37936 16658 37964 17682
rect 38108 17672 38160 17678
rect 38108 17614 38160 17620
rect 38120 17270 38148 17614
rect 38108 17264 38160 17270
rect 38108 17206 38160 17212
rect 37924 16652 37976 16658
rect 37924 16594 37976 16600
rect 37464 12640 37516 12646
rect 37464 12582 37516 12588
rect 37476 9178 37504 12582
rect 37936 11762 37964 16594
rect 37924 11756 37976 11762
rect 37924 11698 37976 11704
rect 37936 11218 37964 11698
rect 37924 11212 37976 11218
rect 37924 11154 37976 11160
rect 37740 10668 37792 10674
rect 37740 10610 37792 10616
rect 37752 10266 37780 10610
rect 37740 10260 37792 10266
rect 37740 10202 37792 10208
rect 38212 9674 38240 17711
rect 38304 12170 38332 21354
rect 38384 20800 38436 20806
rect 38384 20742 38436 20748
rect 38396 20466 38424 20742
rect 38384 20460 38436 20466
rect 38384 20402 38436 20408
rect 38672 19378 38700 21576
rect 38844 21558 38896 21564
rect 38844 20596 38896 20602
rect 38844 20538 38896 20544
rect 38856 20330 38884 20538
rect 38936 20460 38988 20466
rect 38936 20402 38988 20408
rect 38844 20324 38896 20330
rect 38844 20266 38896 20272
rect 38660 19372 38712 19378
rect 38712 19332 38792 19360
rect 38660 19314 38712 19320
rect 38384 19304 38436 19310
rect 38384 19246 38436 19252
rect 38396 18970 38424 19246
rect 38384 18964 38436 18970
rect 38384 18906 38436 18912
rect 38764 18902 38792 19332
rect 38752 18896 38804 18902
rect 38752 18838 38804 18844
rect 38568 18760 38620 18766
rect 38620 18720 38700 18748
rect 38568 18702 38620 18708
rect 38384 18624 38436 18630
rect 38384 18566 38436 18572
rect 38396 18290 38424 18566
rect 38384 18284 38436 18290
rect 38384 18226 38436 18232
rect 38568 18216 38620 18222
rect 38568 18158 38620 18164
rect 38292 12164 38344 12170
rect 38292 12106 38344 12112
rect 38384 11688 38436 11694
rect 38384 11630 38436 11636
rect 38396 10130 38424 11630
rect 38384 10124 38436 10130
rect 38384 10066 38436 10072
rect 38212 9646 38332 9674
rect 38304 9586 38332 9646
rect 37556 9580 37608 9586
rect 37556 9522 37608 9528
rect 38292 9580 38344 9586
rect 38292 9522 38344 9528
rect 37464 9172 37516 9178
rect 37464 9114 37516 9120
rect 37476 8430 37504 9114
rect 37464 8424 37516 8430
rect 37464 8366 37516 8372
rect 37372 7880 37424 7886
rect 37372 7822 37424 7828
rect 37568 7410 37596 9522
rect 37648 9512 37700 9518
rect 37648 9454 37700 9460
rect 37660 8294 37688 9454
rect 37832 9376 37884 9382
rect 37832 9318 37884 9324
rect 38016 9376 38068 9382
rect 38016 9318 38068 9324
rect 37844 9178 37872 9318
rect 37832 9172 37884 9178
rect 37832 9114 37884 9120
rect 37832 8832 37884 8838
rect 37832 8774 37884 8780
rect 37740 8492 37792 8498
rect 37740 8434 37792 8440
rect 37648 8288 37700 8294
rect 37648 8230 37700 8236
rect 37556 7404 37608 7410
rect 37556 7346 37608 7352
rect 37188 7200 37240 7206
rect 37188 7142 37240 7148
rect 37200 6866 37228 7142
rect 37568 6934 37596 7346
rect 37372 6928 37424 6934
rect 37372 6870 37424 6876
rect 37556 6928 37608 6934
rect 37556 6870 37608 6876
rect 37188 6860 37240 6866
rect 37188 6802 37240 6808
rect 37200 6186 37228 6802
rect 37384 6390 37412 6870
rect 37660 6730 37688 8230
rect 37752 7886 37780 8434
rect 37740 7880 37792 7886
rect 37740 7822 37792 7828
rect 37752 7342 37780 7822
rect 37740 7336 37792 7342
rect 37740 7278 37792 7284
rect 37844 6866 37872 8774
rect 38028 8090 38056 9318
rect 38108 9172 38160 9178
rect 38108 9114 38160 9120
rect 38292 9172 38344 9178
rect 38292 9114 38344 9120
rect 38120 8906 38148 9114
rect 38108 8900 38160 8906
rect 38108 8842 38160 8848
rect 38200 8900 38252 8906
rect 38200 8842 38252 8848
rect 38120 8498 38148 8842
rect 38108 8492 38160 8498
rect 38108 8434 38160 8440
rect 38108 8288 38160 8294
rect 38108 8230 38160 8236
rect 38016 8084 38068 8090
rect 38016 8026 38068 8032
rect 38120 7993 38148 8230
rect 38106 7984 38162 7993
rect 38212 7954 38240 8842
rect 38106 7919 38162 7928
rect 38200 7948 38252 7954
rect 38200 7890 38252 7896
rect 38108 7880 38160 7886
rect 38028 7828 38108 7834
rect 38028 7822 38160 7828
rect 38028 7806 38148 7822
rect 38028 7750 38056 7806
rect 38016 7744 38068 7750
rect 38016 7686 38068 7692
rect 38028 6866 38056 7686
rect 38304 7410 38332 9114
rect 38580 8974 38608 18158
rect 38672 16697 38700 18720
rect 38844 18284 38896 18290
rect 38844 18226 38896 18232
rect 38856 18086 38884 18226
rect 38844 18080 38896 18086
rect 38844 18022 38896 18028
rect 38658 16688 38714 16697
rect 38658 16623 38714 16632
rect 38672 10062 38700 16623
rect 38844 10464 38896 10470
rect 38844 10406 38896 10412
rect 38856 10198 38884 10406
rect 38844 10192 38896 10198
rect 38844 10134 38896 10140
rect 38660 10056 38712 10062
rect 38660 9998 38712 10004
rect 38660 9580 38712 9586
rect 38660 9522 38712 9528
rect 38568 8968 38620 8974
rect 38568 8910 38620 8916
rect 38672 8820 38700 9522
rect 38752 8968 38804 8974
rect 38752 8910 38804 8916
rect 38764 8838 38792 8910
rect 38580 8792 38700 8820
rect 38752 8832 38804 8838
rect 38384 7948 38436 7954
rect 38436 7908 38516 7936
rect 38384 7890 38436 7896
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 37832 6860 37884 6866
rect 37832 6802 37884 6808
rect 38016 6860 38068 6866
rect 38016 6802 38068 6808
rect 38304 6798 38332 7346
rect 38384 7200 38436 7206
rect 38384 7142 38436 7148
rect 38396 7002 38424 7142
rect 38384 6996 38436 7002
rect 38384 6938 38436 6944
rect 38292 6792 38344 6798
rect 38292 6734 38344 6740
rect 37648 6724 37700 6730
rect 37648 6666 37700 6672
rect 38488 6662 38516 7908
rect 38476 6656 38528 6662
rect 38476 6598 38528 6604
rect 37372 6384 37424 6390
rect 37372 6326 37424 6332
rect 38580 6254 38608 8792
rect 38752 8774 38804 8780
rect 38658 8528 38714 8537
rect 38658 8463 38660 8472
rect 38712 8463 38714 8472
rect 38660 8434 38712 8440
rect 38948 8362 38976 20402
rect 39028 18760 39080 18766
rect 39028 18702 39080 18708
rect 39040 17202 39068 18702
rect 39212 18692 39264 18698
rect 39212 18634 39264 18640
rect 39224 18358 39252 18634
rect 39212 18352 39264 18358
rect 39212 18294 39264 18300
rect 39316 17218 39344 48622
rect 39408 17338 39436 55830
rect 40052 33998 40080 58278
rect 40144 57458 40172 58958
rect 40236 57934 40264 60998
rect 40972 60858 41000 60998
rect 40960 60852 41012 60858
rect 40960 60794 41012 60800
rect 40224 57928 40276 57934
rect 40224 57870 40276 57876
rect 40132 57452 40184 57458
rect 40132 57394 40184 57400
rect 40592 57316 40644 57322
rect 40592 57258 40644 57264
rect 40604 56982 40632 57258
rect 40592 56976 40644 56982
rect 40592 56918 40644 56924
rect 41064 56846 41092 60998
rect 41340 60722 41368 63200
rect 42076 61198 42104 63200
rect 42812 61198 42840 63200
rect 42064 61192 42116 61198
rect 42064 61134 42116 61140
rect 42800 61192 42852 61198
rect 44100 61180 44128 63294
rect 44270 63294 44588 63322
rect 44270 63200 44326 63294
rect 44456 61260 44508 61266
rect 44456 61202 44508 61208
rect 44180 61192 44232 61198
rect 44100 61152 44180 61180
rect 42800 61134 42852 61140
rect 44180 61134 44232 61140
rect 42064 61056 42116 61062
rect 42064 60998 42116 61004
rect 42800 61056 42852 61062
rect 42800 60998 42852 61004
rect 43720 61056 43772 61062
rect 43720 60998 43772 61004
rect 44272 61056 44324 61062
rect 44272 60998 44324 61004
rect 41328 60716 41380 60722
rect 41328 60658 41380 60664
rect 41604 60512 41656 60518
rect 41604 60454 41656 60460
rect 41616 60314 41644 60454
rect 41604 60308 41656 60314
rect 41604 60250 41656 60256
rect 41052 56840 41104 56846
rect 41052 56782 41104 56788
rect 42076 53145 42104 60998
rect 42708 54120 42760 54126
rect 42708 54062 42760 54068
rect 42062 53136 42118 53145
rect 42062 53071 42118 53080
rect 41604 47660 41656 47666
rect 41604 47602 41656 47608
rect 41512 37936 41564 37942
rect 41512 37878 41564 37884
rect 40868 36100 40920 36106
rect 40868 36042 40920 36048
rect 40040 33992 40092 33998
rect 40040 33934 40092 33940
rect 40592 33992 40644 33998
rect 40592 33934 40644 33940
rect 40500 33924 40552 33930
rect 40500 33866 40552 33872
rect 40512 31754 40540 33866
rect 40604 33522 40632 33934
rect 40592 33516 40644 33522
rect 40592 33458 40644 33464
rect 40144 31726 40540 31754
rect 39856 29028 39908 29034
rect 39856 28970 39908 28976
rect 39580 27124 39632 27130
rect 39580 27066 39632 27072
rect 39488 23112 39540 23118
rect 39488 23054 39540 23060
rect 39500 21962 39528 23054
rect 39488 21956 39540 21962
rect 39488 21898 39540 21904
rect 39396 17332 39448 17338
rect 39396 17274 39448 17280
rect 39028 17196 39080 17202
rect 39316 17190 39436 17218
rect 39028 17138 39080 17144
rect 39040 16640 39068 17138
rect 39120 16652 39172 16658
rect 39040 16612 39120 16640
rect 39120 16594 39172 16600
rect 39304 13456 39356 13462
rect 39304 13398 39356 13404
rect 39120 11144 39172 11150
rect 39120 11086 39172 11092
rect 39028 8832 39080 8838
rect 39028 8774 39080 8780
rect 38936 8356 38988 8362
rect 38936 8298 38988 8304
rect 38948 8090 38976 8298
rect 38752 8084 38804 8090
rect 38752 8026 38804 8032
rect 38936 8084 38988 8090
rect 38936 8026 38988 8032
rect 38660 7472 38712 7478
rect 38658 7440 38660 7449
rect 38712 7440 38714 7449
rect 38764 7410 38792 8026
rect 38844 7948 38896 7954
rect 38844 7890 38896 7896
rect 38658 7375 38714 7384
rect 38752 7404 38804 7410
rect 38752 7346 38804 7352
rect 38660 7200 38712 7206
rect 38660 7142 38712 7148
rect 38672 7002 38700 7142
rect 38660 6996 38712 7002
rect 38660 6938 38712 6944
rect 38764 6798 38792 7346
rect 38856 7342 38884 7890
rect 38844 7336 38896 7342
rect 38844 7278 38896 7284
rect 38856 7206 38884 7278
rect 38844 7200 38896 7206
rect 38844 7142 38896 7148
rect 39040 6866 39068 8774
rect 39132 7256 39160 11086
rect 39212 8832 39264 8838
rect 39212 8774 39264 8780
rect 39224 8566 39252 8774
rect 39212 8560 39264 8566
rect 39212 8502 39264 8508
rect 39212 8424 39264 8430
rect 39212 8366 39264 8372
rect 39224 7410 39252 8366
rect 39316 8106 39344 13398
rect 39408 12434 39436 17190
rect 39408 12406 39528 12434
rect 39396 9104 39448 9110
rect 39396 9046 39448 9052
rect 39408 8566 39436 9046
rect 39396 8560 39448 8566
rect 39396 8502 39448 8508
rect 39316 8078 39436 8106
rect 39212 7404 39264 7410
rect 39212 7346 39264 7352
rect 39212 7268 39264 7274
rect 39132 7228 39212 7256
rect 39212 7210 39264 7216
rect 39028 6860 39080 6866
rect 39028 6802 39080 6808
rect 38752 6792 38804 6798
rect 38752 6734 38804 6740
rect 38568 6248 38620 6254
rect 38568 6190 38620 6196
rect 37188 6180 37240 6186
rect 37188 6122 37240 6128
rect 37372 5296 37424 5302
rect 37372 5238 37424 5244
rect 37004 5160 37056 5166
rect 37004 5102 37056 5108
rect 37096 5160 37148 5166
rect 37096 5102 37148 5108
rect 37280 5092 37332 5098
rect 37280 5034 37332 5040
rect 37188 4616 37240 4622
rect 37188 4558 37240 4564
rect 37096 4548 37148 4554
rect 37096 4490 37148 4496
rect 36912 4208 36964 4214
rect 36912 4150 36964 4156
rect 36268 4140 36320 4146
rect 36268 4082 36320 4088
rect 36280 3942 36308 4082
rect 36360 4072 36412 4078
rect 36360 4014 36412 4020
rect 36268 3936 36320 3942
rect 36268 3878 36320 3884
rect 36372 2774 36400 4014
rect 36924 3534 36952 4150
rect 36912 3528 36964 3534
rect 36912 3470 36964 3476
rect 36544 2848 36596 2854
rect 36544 2790 36596 2796
rect 36004 2230 36124 2258
rect 36280 2746 36400 2774
rect 35900 1420 35952 1426
rect 35900 1362 35952 1368
rect 36004 800 36032 2230
rect 36280 800 36308 2746
rect 36556 800 36584 2790
rect 36820 2576 36872 2582
rect 36820 2518 36872 2524
rect 36832 800 36860 2518
rect 37108 800 37136 4490
rect 37200 4214 37228 4558
rect 37188 4208 37240 4214
rect 37188 4150 37240 4156
rect 37188 3936 37240 3942
rect 37188 3878 37240 3884
rect 37200 3398 37228 3878
rect 37188 3392 37240 3398
rect 37188 3334 37240 3340
rect 37292 2378 37320 5034
rect 37280 2372 37332 2378
rect 37280 2314 37332 2320
rect 37384 800 37412 5238
rect 38568 5228 38620 5234
rect 38568 5170 38620 5176
rect 38660 5228 38712 5234
rect 38660 5170 38712 5176
rect 39120 5228 39172 5234
rect 39120 5170 39172 5176
rect 38580 4622 38608 5170
rect 38568 4616 38620 4622
rect 38568 4558 38620 4564
rect 38476 4480 38528 4486
rect 38476 4422 38528 4428
rect 37556 4140 37608 4146
rect 37556 4082 37608 4088
rect 37464 3936 37516 3942
rect 37464 3878 37516 3884
rect 37476 3058 37504 3878
rect 37568 3738 37596 4082
rect 38200 4072 38252 4078
rect 38200 4014 38252 4020
rect 37556 3732 37608 3738
rect 37556 3674 37608 3680
rect 37648 3596 37700 3602
rect 37648 3538 37700 3544
rect 37464 3052 37516 3058
rect 37464 2994 37516 3000
rect 37660 800 37688 3538
rect 38108 3528 38160 3534
rect 38108 3470 38160 3476
rect 37924 3188 37976 3194
rect 37924 3130 37976 3136
rect 37936 800 37964 3130
rect 38120 2038 38148 3470
rect 38108 2032 38160 2038
rect 38108 1974 38160 1980
rect 38212 800 38240 4014
rect 38488 800 38516 4422
rect 38580 4214 38608 4558
rect 38568 4208 38620 4214
rect 38568 4150 38620 4156
rect 38672 4078 38700 5170
rect 39132 4570 39160 5170
rect 39304 5092 39356 5098
rect 39304 5034 39356 5040
rect 38936 4548 38988 4554
rect 38936 4490 38988 4496
rect 39040 4542 39160 4570
rect 39212 4616 39264 4622
rect 39212 4558 39264 4564
rect 38752 4208 38804 4214
rect 38752 4150 38804 4156
rect 38660 4072 38712 4078
rect 38660 4014 38712 4020
rect 38660 3936 38712 3942
rect 38660 3878 38712 3884
rect 38672 3058 38700 3878
rect 38660 3052 38712 3058
rect 38660 2994 38712 3000
rect 38764 800 38792 4150
rect 38844 4072 38896 4078
rect 38844 4014 38896 4020
rect 38856 3466 38884 4014
rect 38948 3602 38976 4490
rect 38936 3596 38988 3602
rect 38936 3538 38988 3544
rect 38844 3460 38896 3466
rect 38844 3402 38896 3408
rect 39040 800 39068 4542
rect 39120 4480 39172 4486
rect 39120 4422 39172 4428
rect 39132 4078 39160 4422
rect 39120 4072 39172 4078
rect 39120 4014 39172 4020
rect 39120 3392 39172 3398
rect 39118 3360 39120 3369
rect 39172 3360 39174 3369
rect 39118 3295 39174 3304
rect 39224 1986 39252 4558
rect 39316 3058 39344 5034
rect 39408 3670 39436 8078
rect 39500 5681 39528 12406
rect 39486 5672 39542 5681
rect 39486 5607 39542 5616
rect 39592 4758 39620 27066
rect 39672 22976 39724 22982
rect 39670 22944 39672 22953
rect 39764 22976 39816 22982
rect 39724 22944 39726 22953
rect 39764 22918 39816 22924
rect 39670 22879 39726 22888
rect 39776 22250 39804 22918
rect 39684 22222 39804 22250
rect 39684 22030 39712 22222
rect 39672 22024 39724 22030
rect 39672 21966 39724 21972
rect 39672 20052 39724 20058
rect 39672 19994 39724 20000
rect 39684 19854 39712 19994
rect 39672 19848 39724 19854
rect 39672 19790 39724 19796
rect 39764 19168 39816 19174
rect 39764 19110 39816 19116
rect 39672 18284 39724 18290
rect 39776 18272 39804 19110
rect 39724 18244 39804 18272
rect 39672 18226 39724 18232
rect 39764 16992 39816 16998
rect 39764 16934 39816 16940
rect 39672 16584 39724 16590
rect 39672 16526 39724 16532
rect 39684 9518 39712 16526
rect 39776 16114 39804 16934
rect 39764 16108 39816 16114
rect 39764 16050 39816 16056
rect 39672 9512 39724 9518
rect 39672 9454 39724 9460
rect 39764 9172 39816 9178
rect 39764 9114 39816 9120
rect 39776 7954 39804 9114
rect 39764 7948 39816 7954
rect 39764 7890 39816 7896
rect 39764 7812 39816 7818
rect 39764 7754 39816 7760
rect 39776 7478 39804 7754
rect 39764 7472 39816 7478
rect 39764 7414 39816 7420
rect 39672 7404 39724 7410
rect 39672 7346 39724 7352
rect 39684 6934 39712 7346
rect 39672 6928 39724 6934
rect 39672 6870 39724 6876
rect 39868 5370 39896 28970
rect 40040 24404 40092 24410
rect 40040 24346 40092 24352
rect 40052 23594 40080 24346
rect 40040 23588 40092 23594
rect 40040 23530 40092 23536
rect 40040 22160 40092 22166
rect 39960 22108 40040 22114
rect 39960 22102 40092 22108
rect 39960 22086 40080 22102
rect 39960 20641 39988 22086
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 39946 20632 40002 20641
rect 39946 20567 40002 20576
rect 39948 20528 40000 20534
rect 39948 20470 40000 20476
rect 39960 19174 39988 20470
rect 40052 19514 40080 21966
rect 40040 19508 40092 19514
rect 40040 19450 40092 19456
rect 39948 19168 40000 19174
rect 39948 19110 40000 19116
rect 40052 18222 40080 19450
rect 40040 18216 40092 18222
rect 40040 18158 40092 18164
rect 40040 17264 40092 17270
rect 40040 17206 40092 17212
rect 40052 16794 40080 17206
rect 40040 16788 40092 16794
rect 40040 16730 40092 16736
rect 39948 15496 40000 15502
rect 39948 15438 40000 15444
rect 39960 14074 39988 15438
rect 39948 14068 40000 14074
rect 39948 14010 40000 14016
rect 40040 12232 40092 12238
rect 40040 12174 40092 12180
rect 39948 9988 40000 9994
rect 39948 9930 40000 9936
rect 39960 9586 39988 9930
rect 39948 9580 40000 9586
rect 39948 9522 40000 9528
rect 39948 9444 40000 9450
rect 39948 9386 40000 9392
rect 39960 9178 39988 9386
rect 39948 9172 40000 9178
rect 39948 9114 40000 9120
rect 40052 7698 40080 12174
rect 40144 11014 40172 31726
rect 40408 26376 40460 26382
rect 40408 26318 40460 26324
rect 40420 23866 40448 26318
rect 40408 23860 40460 23866
rect 40408 23802 40460 23808
rect 40420 23746 40448 23802
rect 40420 23718 40540 23746
rect 40408 23656 40460 23662
rect 40408 23598 40460 23604
rect 40316 23248 40368 23254
rect 40316 23190 40368 23196
rect 40224 22976 40276 22982
rect 40222 22944 40224 22953
rect 40276 22944 40278 22953
rect 40222 22879 40278 22888
rect 40328 22778 40356 23190
rect 40316 22772 40368 22778
rect 40316 22714 40368 22720
rect 40420 22710 40448 23598
rect 40512 23186 40540 23718
rect 40592 23316 40644 23322
rect 40592 23258 40644 23264
rect 40500 23180 40552 23186
rect 40500 23122 40552 23128
rect 40500 23044 40552 23050
rect 40500 22986 40552 22992
rect 40408 22704 40460 22710
rect 40408 22646 40460 22652
rect 40316 22024 40368 22030
rect 40316 21966 40368 21972
rect 40328 21729 40356 21966
rect 40314 21720 40370 21729
rect 40314 21655 40370 21664
rect 40420 21554 40448 22646
rect 40512 21672 40540 22986
rect 40604 22710 40632 23258
rect 40682 23080 40738 23089
rect 40682 23015 40738 23024
rect 40696 22982 40724 23015
rect 40684 22976 40736 22982
rect 40684 22918 40736 22924
rect 40592 22704 40644 22710
rect 40592 22646 40644 22652
rect 40696 22556 40724 22918
rect 40604 22528 40724 22556
rect 40604 22030 40632 22528
rect 40682 22128 40738 22137
rect 40880 22094 40908 36042
rect 41144 28756 41196 28762
rect 41144 28698 41196 28704
rect 40682 22063 40738 22072
rect 40788 22066 40908 22094
rect 40592 22024 40644 22030
rect 40592 21966 40644 21972
rect 40512 21644 40632 21672
rect 40604 21593 40632 21644
rect 40590 21584 40646 21593
rect 40408 21548 40460 21554
rect 40408 21490 40460 21496
rect 40500 21548 40552 21554
rect 40590 21519 40646 21528
rect 40500 21490 40552 21496
rect 40224 21004 40276 21010
rect 40224 20946 40276 20952
rect 40236 20058 40264 20946
rect 40316 20800 40368 20806
rect 40316 20742 40368 20748
rect 40328 20466 40356 20742
rect 40512 20602 40540 21490
rect 40604 20806 40632 21519
rect 40696 20874 40724 22063
rect 40684 20868 40736 20874
rect 40684 20810 40736 20816
rect 40592 20800 40644 20806
rect 40592 20742 40644 20748
rect 40500 20596 40552 20602
rect 40500 20538 40552 20544
rect 40316 20460 40368 20466
rect 40316 20402 40368 20408
rect 40224 20052 40276 20058
rect 40224 19994 40276 20000
rect 40236 18086 40264 19994
rect 40604 19854 40632 20742
rect 40592 19848 40644 19854
rect 40592 19790 40644 19796
rect 40224 18080 40276 18086
rect 40224 18022 40276 18028
rect 40592 17264 40644 17270
rect 40592 17206 40644 17212
rect 40408 17196 40460 17202
rect 40408 17138 40460 17144
rect 40420 12434 40448 17138
rect 40604 16658 40632 17206
rect 40684 17060 40736 17066
rect 40684 17002 40736 17008
rect 40592 16652 40644 16658
rect 40592 16594 40644 16600
rect 40500 16176 40552 16182
rect 40500 16118 40552 16124
rect 40328 12406 40448 12434
rect 40132 11008 40184 11014
rect 40132 10950 40184 10956
rect 40328 9518 40356 12406
rect 40408 11076 40460 11082
rect 40408 11018 40460 11024
rect 40132 9512 40184 9518
rect 40132 9454 40184 9460
rect 40316 9512 40368 9518
rect 40316 9454 40368 9460
rect 40144 9110 40172 9454
rect 40316 9376 40368 9382
rect 40316 9318 40368 9324
rect 40132 9104 40184 9110
rect 40132 9046 40184 9052
rect 40328 8974 40356 9318
rect 40316 8968 40368 8974
rect 40316 8910 40368 8916
rect 40224 8900 40276 8906
rect 40224 8842 40276 8848
rect 40236 8634 40264 8842
rect 40316 8832 40368 8838
rect 40316 8774 40368 8780
rect 40224 8628 40276 8634
rect 40224 8570 40276 8576
rect 40328 8498 40356 8774
rect 40132 8492 40184 8498
rect 40132 8434 40184 8440
rect 40316 8492 40368 8498
rect 40316 8434 40368 8440
rect 40144 8090 40172 8434
rect 40132 8084 40184 8090
rect 40132 8026 40184 8032
rect 40144 7818 40172 8026
rect 40132 7812 40184 7818
rect 40132 7754 40184 7760
rect 40052 7670 40264 7698
rect 39946 7440 40002 7449
rect 39946 7375 40002 7384
rect 39960 7342 39988 7375
rect 39948 7336 40000 7342
rect 39948 7278 40000 7284
rect 39856 5364 39908 5370
rect 39856 5306 39908 5312
rect 40040 5228 40092 5234
rect 40040 5170 40092 5176
rect 39580 4752 39632 4758
rect 39580 4694 39632 4700
rect 39488 4684 39540 4690
rect 39488 4626 39540 4632
rect 39396 3664 39448 3670
rect 39396 3606 39448 3612
rect 39500 3534 39528 4626
rect 39948 4140 40000 4146
rect 39948 4082 40000 4088
rect 39672 3664 39724 3670
rect 39672 3606 39724 3612
rect 39488 3528 39540 3534
rect 39488 3470 39540 3476
rect 39396 3120 39448 3126
rect 39396 3062 39448 3068
rect 39304 3052 39356 3058
rect 39304 2994 39356 3000
rect 39408 2446 39436 3062
rect 39500 2446 39528 3470
rect 39684 3126 39712 3606
rect 39960 3194 39988 4082
rect 39948 3188 40000 3194
rect 39948 3130 40000 3136
rect 39672 3120 39724 3126
rect 39672 3062 39724 3068
rect 39580 3052 39632 3058
rect 39580 2994 39632 3000
rect 39396 2440 39448 2446
rect 39396 2382 39448 2388
rect 39488 2440 39540 2446
rect 39488 2382 39540 2388
rect 39224 1958 39344 1986
rect 39316 800 39344 1958
rect 39592 800 39620 2994
rect 40052 2774 40080 5170
rect 40132 4072 40184 4078
rect 40132 4014 40184 4020
rect 40144 3534 40172 4014
rect 40236 3942 40264 7670
rect 40224 3936 40276 3942
rect 40224 3878 40276 3884
rect 40420 3670 40448 11018
rect 40512 9586 40540 16118
rect 40500 9580 40552 9586
rect 40500 9522 40552 9528
rect 40500 9444 40552 9450
rect 40500 9386 40552 9392
rect 40512 8974 40540 9386
rect 40500 8968 40552 8974
rect 40500 8910 40552 8916
rect 40512 8430 40540 8910
rect 40500 8424 40552 8430
rect 40500 8366 40552 8372
rect 40696 3942 40724 17002
rect 40788 12646 40816 22066
rect 41052 19848 41104 19854
rect 41052 19790 41104 19796
rect 41064 18834 41092 19790
rect 41052 18828 41104 18834
rect 41052 18770 41104 18776
rect 41064 18290 41092 18770
rect 41052 18284 41104 18290
rect 41052 18226 41104 18232
rect 41064 17542 41092 18226
rect 41052 17536 41104 17542
rect 41052 17478 41104 17484
rect 41064 17338 41092 17478
rect 40960 17332 41012 17338
rect 40960 17274 41012 17280
rect 41052 17332 41104 17338
rect 41052 17274 41104 17280
rect 40868 16516 40920 16522
rect 40868 16458 40920 16464
rect 40880 15978 40908 16458
rect 40868 15972 40920 15978
rect 40868 15914 40920 15920
rect 40776 12640 40828 12646
rect 40776 12582 40828 12588
rect 40972 12434 41000 17274
rect 41156 17218 41184 28698
rect 41420 22976 41472 22982
rect 41420 22918 41472 22924
rect 41328 20936 41380 20942
rect 41328 20878 41380 20884
rect 41236 20052 41288 20058
rect 41236 19994 41288 20000
rect 41248 19854 41276 19994
rect 41340 19922 41368 20878
rect 41328 19916 41380 19922
rect 41328 19858 41380 19864
rect 41236 19848 41288 19854
rect 41236 19790 41288 19796
rect 41248 18358 41276 19790
rect 41236 18352 41288 18358
rect 41236 18294 41288 18300
rect 41236 17672 41288 17678
rect 41236 17614 41288 17620
rect 41248 17338 41276 17614
rect 41236 17332 41288 17338
rect 41236 17274 41288 17280
rect 40880 12406 41000 12434
rect 41064 17190 41184 17218
rect 41432 17202 41460 22918
rect 41420 17196 41472 17202
rect 40684 3936 40736 3942
rect 40684 3878 40736 3884
rect 40408 3664 40460 3670
rect 40408 3606 40460 3612
rect 40132 3528 40184 3534
rect 40132 3470 40184 3476
rect 40880 3126 40908 12406
rect 41064 9704 41092 17190
rect 41420 17138 41472 17144
rect 41142 13696 41198 13705
rect 41142 13631 41198 13640
rect 40972 9676 41092 9704
rect 40972 5370 41000 9676
rect 41052 9580 41104 9586
rect 41052 9522 41104 9528
rect 41064 9178 41092 9522
rect 41052 9172 41104 9178
rect 41052 9114 41104 9120
rect 41052 9036 41104 9042
rect 41052 8978 41104 8984
rect 41064 8838 41092 8978
rect 41052 8832 41104 8838
rect 41052 8774 41104 8780
rect 40960 5364 41012 5370
rect 40960 5306 41012 5312
rect 41050 3632 41106 3641
rect 41050 3567 41052 3576
rect 41104 3567 41106 3576
rect 41052 3538 41104 3544
rect 40868 3120 40920 3126
rect 40868 3062 40920 3068
rect 40408 3052 40460 3058
rect 40408 2994 40460 3000
rect 39868 2746 40080 2774
rect 39868 800 39896 2746
rect 40132 2440 40184 2446
rect 40132 2382 40184 2388
rect 40144 800 40172 2382
rect 40420 800 40448 2994
rect 40684 2848 40736 2854
rect 40684 2790 40736 2796
rect 40500 2372 40552 2378
rect 40500 2314 40552 2320
rect 40512 1970 40540 2314
rect 40500 1964 40552 1970
rect 40500 1906 40552 1912
rect 40696 800 40724 2790
rect 41156 2650 41184 13631
rect 41524 6914 41552 37878
rect 41616 11744 41644 47602
rect 42524 39364 42576 39370
rect 42524 39306 42576 39312
rect 41696 37460 41748 37466
rect 41696 37402 41748 37408
rect 41708 35894 41736 37402
rect 41708 35866 41828 35894
rect 41696 28960 41748 28966
rect 41696 28902 41748 28908
rect 41708 12434 41736 28902
rect 41800 21350 41828 35866
rect 42340 31952 42392 31958
rect 42340 31894 42392 31900
rect 42352 30258 42380 31894
rect 42432 31816 42484 31822
rect 42432 31758 42484 31764
rect 42444 31142 42472 31758
rect 42432 31136 42484 31142
rect 42432 31078 42484 31084
rect 42340 30252 42392 30258
rect 42340 30194 42392 30200
rect 42064 27532 42116 27538
rect 42064 27474 42116 27480
rect 41880 23724 41932 23730
rect 41880 23666 41932 23672
rect 41892 23322 41920 23666
rect 41880 23316 41932 23322
rect 41880 23258 41932 23264
rect 41788 21344 41840 21350
rect 41788 21286 41840 21292
rect 41800 21010 41828 21286
rect 41788 21004 41840 21010
rect 41788 20946 41840 20952
rect 41880 19916 41932 19922
rect 41880 19858 41932 19864
rect 41892 18630 41920 19858
rect 41880 18624 41932 18630
rect 41880 18566 41932 18572
rect 41788 18284 41840 18290
rect 41788 18226 41840 18232
rect 41800 17882 41828 18226
rect 41788 17876 41840 17882
rect 41788 17818 41840 17824
rect 41708 12406 41920 12434
rect 41616 11716 41828 11744
rect 41696 11008 41748 11014
rect 41696 10950 41748 10956
rect 41604 9444 41656 9450
rect 41604 9386 41656 9392
rect 41616 8566 41644 9386
rect 41604 8560 41656 8566
rect 41604 8502 41656 8508
rect 41524 6886 41644 6914
rect 41420 4548 41472 4554
rect 41420 4490 41472 4496
rect 41328 3052 41380 3058
rect 41328 2994 41380 3000
rect 41340 2774 41368 2994
rect 41432 2854 41460 4490
rect 41512 4140 41564 4146
rect 41512 4082 41564 4088
rect 41420 2848 41472 2854
rect 41420 2790 41472 2796
rect 41248 2746 41368 2774
rect 41144 2644 41196 2650
rect 41144 2586 41196 2592
rect 41144 2440 41196 2446
rect 40972 2400 41144 2428
rect 40972 800 41000 2400
rect 41144 2382 41196 2388
rect 41248 800 41276 2746
rect 41524 800 41552 4082
rect 41616 3126 41644 6886
rect 41708 4826 41736 10950
rect 41696 4820 41748 4826
rect 41696 4762 41748 4768
rect 41800 4078 41828 11716
rect 41788 4072 41840 4078
rect 41788 4014 41840 4020
rect 41892 3602 41920 12406
rect 42076 5098 42104 27474
rect 42536 24970 42564 39306
rect 42616 32292 42668 32298
rect 42616 32234 42668 32240
rect 42628 31822 42656 32234
rect 42616 31816 42668 31822
rect 42616 31758 42668 31764
rect 42536 24942 42656 24970
rect 42524 23316 42576 23322
rect 42524 23258 42576 23264
rect 42536 23225 42564 23258
rect 42522 23216 42578 23225
rect 42522 23151 42578 23160
rect 42628 22094 42656 24942
rect 42536 22066 42656 22094
rect 42432 18624 42484 18630
rect 42432 18566 42484 18572
rect 42248 17808 42300 17814
rect 42248 17750 42300 17756
rect 42156 10056 42208 10062
rect 42156 9998 42208 10004
rect 42168 5370 42196 9998
rect 42156 5364 42208 5370
rect 42156 5306 42208 5312
rect 42064 5092 42116 5098
rect 42064 5034 42116 5040
rect 42064 4548 42116 4554
rect 42064 4490 42116 4496
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 41788 3528 41840 3534
rect 41788 3470 41840 3476
rect 41604 3120 41656 3126
rect 41604 3062 41656 3068
rect 41800 800 41828 3470
rect 42076 800 42104 4490
rect 42260 3942 42288 17750
rect 42444 17678 42472 18566
rect 42432 17672 42484 17678
rect 42432 17614 42484 17620
rect 42444 16590 42472 17614
rect 42432 16584 42484 16590
rect 42432 16526 42484 16532
rect 42536 4146 42564 22066
rect 42616 19372 42668 19378
rect 42616 19314 42668 19320
rect 42628 18290 42656 19314
rect 42616 18284 42668 18290
rect 42616 18226 42668 18232
rect 42720 11762 42748 54062
rect 42812 32570 42840 60998
rect 43444 55616 43496 55622
rect 43444 55558 43496 55564
rect 43456 55282 43484 55558
rect 43536 55412 43588 55418
rect 43536 55354 43588 55360
rect 43444 55276 43496 55282
rect 43444 55218 43496 55224
rect 43260 54188 43312 54194
rect 43260 54130 43312 54136
rect 43168 36780 43220 36786
rect 43168 36722 43220 36728
rect 43180 33538 43208 36722
rect 43272 34406 43300 54130
rect 43260 34400 43312 34406
rect 43260 34342 43312 34348
rect 43180 33510 43392 33538
rect 43364 32910 43392 33510
rect 42892 32904 42944 32910
rect 42892 32846 42944 32852
rect 43076 32904 43128 32910
rect 43076 32846 43128 32852
rect 43352 32904 43404 32910
rect 43352 32846 43404 32852
rect 42800 32564 42852 32570
rect 42800 32506 42852 32512
rect 42904 30394 42932 32846
rect 43088 31278 43116 32846
rect 43364 32366 43392 32846
rect 43352 32360 43404 32366
rect 43352 32302 43404 32308
rect 43444 31816 43496 31822
rect 43444 31758 43496 31764
rect 43076 31272 43128 31278
rect 43076 31214 43128 31220
rect 42892 30388 42944 30394
rect 42892 30330 42944 30336
rect 43168 30388 43220 30394
rect 43168 30330 43220 30336
rect 43076 29708 43128 29714
rect 43076 29650 43128 29656
rect 43088 29306 43116 29650
rect 43180 29646 43208 30330
rect 43456 29646 43484 31758
rect 43168 29640 43220 29646
rect 43168 29582 43220 29588
rect 43444 29640 43496 29646
rect 43444 29582 43496 29588
rect 43076 29300 43128 29306
rect 43076 29242 43128 29248
rect 42892 28552 42944 28558
rect 42892 28494 42944 28500
rect 42800 23112 42852 23118
rect 42798 23080 42800 23089
rect 42852 23080 42854 23089
rect 42798 23015 42854 23024
rect 42812 20942 42840 23015
rect 42800 20936 42852 20942
rect 42800 20878 42852 20884
rect 42708 11756 42760 11762
rect 42708 11698 42760 11704
rect 42904 6914 42932 28494
rect 43352 24064 43404 24070
rect 43352 24006 43404 24012
rect 43364 23118 43392 24006
rect 43352 23112 43404 23118
rect 43352 23054 43404 23060
rect 43260 22772 43312 22778
rect 43260 22714 43312 22720
rect 43168 22568 43220 22574
rect 43168 22510 43220 22516
rect 43180 18766 43208 22510
rect 43272 21962 43300 22714
rect 43352 22024 43404 22030
rect 43404 21984 43484 22012
rect 43352 21966 43404 21972
rect 43260 21956 43312 21962
rect 43260 21898 43312 21904
rect 43352 21480 43404 21486
rect 43352 21422 43404 21428
rect 43364 21010 43392 21422
rect 43456 21010 43484 21984
rect 43352 21004 43404 21010
rect 43352 20946 43404 20952
rect 43444 21004 43496 21010
rect 43444 20946 43496 20952
rect 43364 19378 43392 20946
rect 43456 20466 43484 20946
rect 43444 20460 43496 20466
rect 43444 20402 43496 20408
rect 43352 19372 43404 19378
rect 43352 19314 43404 19320
rect 43444 19236 43496 19242
rect 43444 19178 43496 19184
rect 43168 18760 43220 18766
rect 43168 18702 43220 18708
rect 43180 18290 43208 18702
rect 43456 18630 43484 19178
rect 43444 18624 43496 18630
rect 43444 18566 43496 18572
rect 43168 18284 43220 18290
rect 43168 18226 43220 18232
rect 42812 6886 42932 6914
rect 42524 4140 42576 4146
rect 42524 4082 42576 4088
rect 42248 3936 42300 3942
rect 42248 3878 42300 3884
rect 42614 3768 42670 3777
rect 42614 3703 42670 3712
rect 42628 3602 42656 3703
rect 42616 3596 42668 3602
rect 42616 3538 42668 3544
rect 42812 3194 42840 6886
rect 43180 5302 43208 18226
rect 43260 12640 43312 12646
rect 43260 12582 43312 12588
rect 43168 5296 43220 5302
rect 43168 5238 43220 5244
rect 43272 4758 43300 12582
rect 43444 11756 43496 11762
rect 43444 11698 43496 11704
rect 43352 9036 43404 9042
rect 43352 8978 43404 8984
rect 43364 8838 43392 8978
rect 43352 8832 43404 8838
rect 43352 8774 43404 8780
rect 43260 4752 43312 4758
rect 43260 4694 43312 4700
rect 42892 4548 42944 4554
rect 42892 4490 42944 4496
rect 42984 4548 43036 4554
rect 42984 4490 43036 4496
rect 43168 4548 43220 4554
rect 43168 4490 43220 4496
rect 42904 3534 42932 4490
rect 42892 3528 42944 3534
rect 42892 3470 42944 3476
rect 42800 3188 42852 3194
rect 42800 3130 42852 3136
rect 42340 2984 42392 2990
rect 42340 2926 42392 2932
rect 42352 800 42380 2926
rect 42616 2304 42668 2310
rect 42996 2258 43024 4490
rect 43076 4004 43128 4010
rect 43076 3946 43128 3952
rect 43088 3233 43116 3946
rect 43074 3224 43130 3233
rect 43074 3159 43130 3168
rect 42616 2246 42668 2252
rect 42628 800 42656 2246
rect 42904 2230 43024 2258
rect 42904 800 42932 2230
rect 43180 800 43208 4490
rect 43260 4140 43312 4146
rect 43312 4100 43392 4128
rect 43260 4082 43312 4088
rect 43364 3466 43392 4100
rect 43456 3534 43484 11698
rect 43444 3528 43496 3534
rect 43444 3470 43496 3476
rect 43352 3460 43404 3466
rect 43352 3402 43404 3408
rect 43364 3369 43392 3402
rect 43350 3360 43406 3369
rect 43350 3295 43406 3304
rect 43364 3097 43392 3295
rect 43350 3088 43406 3097
rect 43350 3023 43406 3032
rect 43364 2378 43392 3023
rect 43444 2848 43496 2854
rect 43444 2790 43496 2796
rect 43352 2372 43404 2378
rect 43352 2314 43404 2320
rect 43456 800 43484 2790
rect 43548 2446 43576 55354
rect 43732 51338 43760 60998
rect 44088 59016 44140 59022
rect 44088 58958 44140 58964
rect 43996 58540 44048 58546
rect 43996 58482 44048 58488
rect 43904 58404 43956 58410
rect 43904 58346 43956 58352
rect 43916 58002 43944 58346
rect 44008 58002 44036 58482
rect 43904 57996 43956 58002
rect 43904 57938 43956 57944
rect 43996 57996 44048 58002
rect 43996 57938 44048 57944
rect 43812 57928 43864 57934
rect 43812 57870 43864 57876
rect 43824 56982 43852 57870
rect 43812 56976 43864 56982
rect 43812 56918 43864 56924
rect 43824 55282 43852 56918
rect 44008 56846 44036 57938
rect 44100 57934 44128 58958
rect 44088 57928 44140 57934
rect 44088 57870 44140 57876
rect 44088 57792 44140 57798
rect 44088 57734 44140 57740
rect 43996 56840 44048 56846
rect 43916 56788 43996 56794
rect 43916 56782 44048 56788
rect 43916 56766 44036 56782
rect 43812 55276 43864 55282
rect 43812 55218 43864 55224
rect 43916 55214 43944 56766
rect 43996 56704 44048 56710
rect 43996 56646 44048 56652
rect 44008 55962 44036 56646
rect 43996 55956 44048 55962
rect 43996 55898 44048 55904
rect 43904 55208 43956 55214
rect 43904 55150 43956 55156
rect 43916 54126 43944 55150
rect 43904 54120 43956 54126
rect 43904 54062 43956 54068
rect 43720 51332 43772 51338
rect 43720 51274 43772 51280
rect 43916 37126 43944 54062
rect 44100 52698 44128 57734
rect 44088 52692 44140 52698
rect 44088 52634 44140 52640
rect 44088 37188 44140 37194
rect 44088 37130 44140 37136
rect 43904 37120 43956 37126
rect 43904 37062 43956 37068
rect 44100 33862 44128 37130
rect 44088 33856 44140 33862
rect 44088 33798 44140 33804
rect 43996 33040 44048 33046
rect 43996 32982 44048 32988
rect 44008 31822 44036 32982
rect 44100 32502 44128 33798
rect 44284 32842 44312 60998
rect 44468 56846 44496 61202
rect 44560 61198 44588 63294
rect 45006 63294 45508 63322
rect 45006 63200 45062 63294
rect 45480 61282 45508 63294
rect 45742 63294 46152 63322
rect 45742 63200 45798 63294
rect 45480 61254 45600 61282
rect 45572 61198 45600 61254
rect 46124 61198 46152 63294
rect 46478 63294 46704 63322
rect 46478 63200 46534 63294
rect 44548 61192 44600 61198
rect 44548 61134 44600 61140
rect 45560 61192 45612 61198
rect 45560 61134 45612 61140
rect 46112 61192 46164 61198
rect 46112 61134 46164 61140
rect 45376 61056 45428 61062
rect 45376 60998 45428 61004
rect 46112 61056 46164 61062
rect 46112 60998 46164 61004
rect 44824 58880 44876 58886
rect 44824 58822 44876 58828
rect 44456 56840 44508 56846
rect 44456 56782 44508 56788
rect 44272 32836 44324 32842
rect 44272 32778 44324 32784
rect 44088 32496 44140 32502
rect 44088 32438 44140 32444
rect 44100 31906 44128 32438
rect 44732 32428 44784 32434
rect 44732 32370 44784 32376
rect 44456 32360 44508 32366
rect 44456 32302 44508 32308
rect 44468 31958 44496 32302
rect 44744 31958 44772 32370
rect 44456 31952 44508 31958
rect 44100 31878 44220 31906
rect 44456 31894 44508 31900
rect 44732 31952 44784 31958
rect 44732 31894 44784 31900
rect 43996 31816 44048 31822
rect 43996 31758 44048 31764
rect 44088 31816 44140 31822
rect 44088 31758 44140 31764
rect 44100 31210 44128 31758
rect 44192 31754 44220 31878
rect 44180 31748 44232 31754
rect 44180 31690 44232 31696
rect 44088 31204 44140 31210
rect 44088 31146 44140 31152
rect 43812 30864 43864 30870
rect 43812 30806 43864 30812
rect 43824 29850 43852 30806
rect 43812 29844 43864 29850
rect 43812 29786 43864 29792
rect 44640 29572 44692 29578
rect 44640 29514 44692 29520
rect 43628 29504 43680 29510
rect 43628 29446 43680 29452
rect 43640 4826 43668 29446
rect 43996 28552 44048 28558
rect 43996 28494 44048 28500
rect 44008 23526 44036 28494
rect 44180 28212 44232 28218
rect 44180 28154 44232 28160
rect 43996 23520 44048 23526
rect 43996 23462 44048 23468
rect 44008 23186 44036 23462
rect 43996 23180 44048 23186
rect 43996 23122 44048 23128
rect 43720 23112 43772 23118
rect 43904 23112 43956 23118
rect 43720 23054 43772 23060
rect 43902 23080 43904 23089
rect 43956 23080 43958 23089
rect 43732 22506 43760 23054
rect 43902 23015 43958 23024
rect 43812 22636 43864 22642
rect 43812 22578 43864 22584
rect 43720 22500 43772 22506
rect 43720 22442 43772 22448
rect 43824 21894 43852 22578
rect 43996 22024 44048 22030
rect 43996 21966 44048 21972
rect 43812 21888 43864 21894
rect 43812 21830 43864 21836
rect 43904 21888 43956 21894
rect 44008 21865 44036 21966
rect 43904 21830 43956 21836
rect 43994 21856 44050 21865
rect 43916 21593 43944 21830
rect 43994 21791 44050 21800
rect 43902 21584 43958 21593
rect 43902 21519 43958 21528
rect 43996 18896 44048 18902
rect 43996 18838 44048 18844
rect 43904 18692 43956 18698
rect 43904 18634 43956 18640
rect 43916 16697 43944 18634
rect 44008 18630 44036 18838
rect 43996 18624 44048 18630
rect 43996 18566 44048 18572
rect 43996 18080 44048 18086
rect 43996 18022 44048 18028
rect 44008 17678 44036 18022
rect 43996 17672 44048 17678
rect 43996 17614 44048 17620
rect 43902 16688 43958 16697
rect 43902 16623 43958 16632
rect 43812 5228 43864 5234
rect 43812 5170 43864 5176
rect 43996 5228 44048 5234
rect 43996 5170 44048 5176
rect 43628 4820 43680 4826
rect 43628 4762 43680 4768
rect 43718 3632 43774 3641
rect 43718 3567 43774 3576
rect 43732 3534 43760 3567
rect 43720 3528 43772 3534
rect 43720 3470 43772 3476
rect 43824 2666 43852 5170
rect 43904 4140 43956 4146
rect 43904 4082 43956 4088
rect 43916 3602 43944 4082
rect 43904 3596 43956 3602
rect 43904 3538 43956 3544
rect 43904 3460 43956 3466
rect 43904 3402 43956 3408
rect 43916 3194 43944 3402
rect 43904 3188 43956 3194
rect 43904 3130 43956 3136
rect 43732 2638 43852 2666
rect 43536 2440 43588 2446
rect 43536 2382 43588 2388
rect 43732 800 43760 2638
rect 44008 800 44036 5170
rect 44192 4758 44220 28154
rect 44652 24342 44680 29514
rect 44836 27674 44864 58822
rect 45388 57322 45416 60998
rect 45376 57316 45428 57322
rect 45376 57258 45428 57264
rect 44916 55956 44968 55962
rect 44916 55898 44968 55904
rect 44824 27668 44876 27674
rect 44824 27610 44876 27616
rect 44640 24336 44692 24342
rect 44640 24278 44692 24284
rect 44548 24200 44600 24206
rect 44548 24142 44600 24148
rect 44456 24132 44508 24138
rect 44456 24074 44508 24080
rect 44364 23724 44416 23730
rect 44364 23666 44416 23672
rect 44376 23322 44404 23666
rect 44468 23526 44496 24074
rect 44560 23662 44588 24142
rect 44652 24070 44680 24278
rect 44824 24268 44876 24274
rect 44824 24210 44876 24216
rect 44640 24064 44692 24070
rect 44640 24006 44692 24012
rect 44640 23724 44692 23730
rect 44640 23666 44692 23672
rect 44548 23656 44600 23662
rect 44548 23598 44600 23604
rect 44456 23520 44508 23526
rect 44456 23462 44508 23468
rect 44364 23316 44416 23322
rect 44364 23258 44416 23264
rect 44364 23112 44416 23118
rect 44364 23054 44416 23060
rect 44272 22432 44324 22438
rect 44272 22374 44324 22380
rect 44284 21554 44312 22374
rect 44376 22030 44404 23054
rect 44560 22642 44588 23598
rect 44548 22636 44600 22642
rect 44548 22578 44600 22584
rect 44560 22094 44588 22578
rect 44468 22066 44588 22094
rect 44364 22024 44416 22030
rect 44364 21966 44416 21972
rect 44272 21548 44324 21554
rect 44272 21490 44324 21496
rect 44272 19372 44324 19378
rect 44272 19314 44324 19320
rect 44376 19334 44404 21966
rect 44468 21146 44496 22066
rect 44456 21140 44508 21146
rect 44456 21082 44508 21088
rect 44652 21010 44680 23666
rect 44732 22772 44784 22778
rect 44732 22714 44784 22720
rect 44744 22642 44772 22714
rect 44732 22636 44784 22642
rect 44732 22578 44784 22584
rect 44640 21004 44692 21010
rect 44640 20946 44692 20952
rect 44284 18834 44312 19314
rect 44376 19306 44496 19334
rect 44364 19168 44416 19174
rect 44364 19110 44416 19116
rect 44376 18902 44404 19110
rect 44364 18896 44416 18902
rect 44364 18838 44416 18844
rect 44272 18828 44324 18834
rect 44272 18770 44324 18776
rect 44468 18766 44496 19306
rect 44456 18760 44508 18766
rect 44456 18702 44508 18708
rect 44272 18148 44324 18154
rect 44272 18090 44324 18096
rect 44180 4752 44232 4758
rect 44180 4694 44232 4700
rect 44284 3738 44312 18090
rect 44836 13802 44864 24210
rect 44824 13796 44876 13802
rect 44824 13738 44876 13744
rect 44824 9716 44876 9722
rect 44824 9658 44876 9664
rect 44732 5024 44784 5030
rect 44732 4966 44784 4972
rect 44364 4548 44416 4554
rect 44364 4490 44416 4496
rect 44272 3732 44324 3738
rect 44272 3674 44324 3680
rect 44272 3528 44324 3534
rect 44272 3470 44324 3476
rect 44284 3058 44312 3470
rect 44272 3052 44324 3058
rect 44272 2994 44324 3000
rect 44284 2446 44312 2994
rect 44272 2440 44324 2446
rect 44272 2382 44324 2388
rect 44376 2258 44404 4490
rect 44456 3732 44508 3738
rect 44456 3674 44508 3680
rect 44468 2990 44496 3674
rect 44640 3596 44692 3602
rect 44640 3538 44692 3544
rect 44548 3392 44600 3398
rect 44548 3334 44600 3340
rect 44456 2984 44508 2990
rect 44456 2926 44508 2932
rect 44284 2230 44404 2258
rect 44284 800 44312 2230
rect 44560 800 44588 3334
rect 44652 2650 44680 3538
rect 44640 2644 44692 2650
rect 44640 2586 44692 2592
rect 44744 2378 44772 4966
rect 44836 2922 44864 9658
rect 44928 3058 44956 55898
rect 46020 52692 46072 52698
rect 46020 52634 46072 52640
rect 45928 44940 45980 44946
rect 45928 44882 45980 44888
rect 45376 37324 45428 37330
rect 45376 37266 45428 37272
rect 45192 37256 45244 37262
rect 45192 37198 45244 37204
rect 45008 24608 45060 24614
rect 45008 24550 45060 24556
rect 45020 24274 45048 24550
rect 45008 24268 45060 24274
rect 45008 24210 45060 24216
rect 45100 19780 45152 19786
rect 45100 19722 45152 19728
rect 45112 19446 45140 19722
rect 45100 19440 45152 19446
rect 45100 19382 45152 19388
rect 45006 14920 45062 14929
rect 45006 14855 45062 14864
rect 45020 6914 45048 14855
rect 45112 9994 45140 19382
rect 45100 9988 45152 9994
rect 45100 9930 45152 9936
rect 45020 6886 45140 6914
rect 45008 4480 45060 4486
rect 45008 4422 45060 4428
rect 45020 3210 45048 4422
rect 45112 3602 45140 6886
rect 45204 4758 45232 37198
rect 45388 36922 45416 37266
rect 45652 37120 45704 37126
rect 45652 37062 45704 37068
rect 45376 36916 45428 36922
rect 45376 36858 45428 36864
rect 45664 36854 45692 37062
rect 45652 36848 45704 36854
rect 45652 36790 45704 36796
rect 45744 32360 45796 32366
rect 45744 32302 45796 32308
rect 45652 27668 45704 27674
rect 45652 27610 45704 27616
rect 45284 24812 45336 24818
rect 45284 24754 45336 24760
rect 45468 24812 45520 24818
rect 45468 24754 45520 24760
rect 45296 24614 45324 24754
rect 45284 24608 45336 24614
rect 45284 24550 45336 24556
rect 45376 22160 45428 22166
rect 45374 22128 45376 22137
rect 45428 22128 45430 22137
rect 45374 22063 45430 22072
rect 45374 21856 45430 21865
rect 45374 21791 45430 21800
rect 45388 21350 45416 21791
rect 45376 21344 45428 21350
rect 45376 21286 45428 21292
rect 45376 19780 45428 19786
rect 45376 19722 45428 19728
rect 45388 19514 45416 19722
rect 45376 19508 45428 19514
rect 45376 19450 45428 19456
rect 45388 18834 45416 19450
rect 45376 18828 45428 18834
rect 45376 18770 45428 18776
rect 45480 6914 45508 24754
rect 45560 22772 45612 22778
rect 45560 22714 45612 22720
rect 45572 22030 45600 22714
rect 45560 22024 45612 22030
rect 45560 21966 45612 21972
rect 45560 20800 45612 20806
rect 45560 20742 45612 20748
rect 45572 20466 45600 20742
rect 45560 20460 45612 20466
rect 45560 20402 45612 20408
rect 45572 17338 45600 20402
rect 45560 17332 45612 17338
rect 45560 17274 45612 17280
rect 45388 6886 45508 6914
rect 45192 4752 45244 4758
rect 45192 4694 45244 4700
rect 45192 4072 45244 4078
rect 45192 4014 45244 4020
rect 45204 3618 45232 4014
rect 45100 3596 45152 3602
rect 45204 3590 45324 3618
rect 45100 3538 45152 3544
rect 45192 3528 45244 3534
rect 45190 3496 45192 3505
rect 45244 3496 45246 3505
rect 45190 3431 45246 3440
rect 45020 3182 45232 3210
rect 45008 3120 45060 3126
rect 45008 3062 45060 3068
rect 45098 3088 45154 3097
rect 44916 3052 44968 3058
rect 44916 2994 44968 3000
rect 44914 2952 44970 2961
rect 44824 2916 44876 2922
rect 44914 2887 44970 2896
rect 44824 2858 44876 2864
rect 44928 2854 44956 2887
rect 44916 2848 44968 2854
rect 44916 2790 44968 2796
rect 44732 2372 44784 2378
rect 44732 2314 44784 2320
rect 45020 1578 45048 3062
rect 45098 3023 45100 3032
rect 45152 3023 45154 3032
rect 45100 2994 45152 3000
rect 45112 2650 45140 2994
rect 45100 2644 45152 2650
rect 45100 2586 45152 2592
rect 45204 2530 45232 3182
rect 45296 2854 45324 3590
rect 45284 2848 45336 2854
rect 45284 2790 45336 2796
rect 45388 2650 45416 6886
rect 45468 4684 45520 4690
rect 45468 4626 45520 4632
rect 45284 2644 45336 2650
rect 45284 2586 45336 2592
rect 45376 2644 45428 2650
rect 45376 2586 45428 2592
rect 44836 1550 45048 1578
rect 45112 2502 45232 2530
rect 44836 800 44864 1550
rect 45112 800 45140 2502
rect 45296 2446 45324 2586
rect 45192 2440 45244 2446
rect 45192 2382 45244 2388
rect 45284 2440 45336 2446
rect 45284 2382 45336 2388
rect 45204 2106 45232 2382
rect 45480 2360 45508 4626
rect 45664 4146 45692 27610
rect 45756 24750 45784 32302
rect 45836 31816 45888 31822
rect 45836 31758 45888 31764
rect 45744 24744 45796 24750
rect 45744 24686 45796 24692
rect 45756 20466 45784 24686
rect 45848 22778 45876 31758
rect 45836 22772 45888 22778
rect 45836 22714 45888 22720
rect 45744 20460 45796 20466
rect 45744 20402 45796 20408
rect 45836 20256 45888 20262
rect 45836 20198 45888 20204
rect 45848 19854 45876 20198
rect 45940 19922 45968 44882
rect 45928 19916 45980 19922
rect 45928 19858 45980 19864
rect 45836 19848 45888 19854
rect 45836 19790 45888 19796
rect 45928 4616 45980 4622
rect 45928 4558 45980 4564
rect 45744 4480 45796 4486
rect 45744 4422 45796 4428
rect 45652 4140 45704 4146
rect 45652 4082 45704 4088
rect 45560 3596 45612 3602
rect 45560 3538 45612 3544
rect 45572 2446 45600 3538
rect 45756 3534 45784 4422
rect 45836 3596 45888 3602
rect 45836 3538 45888 3544
rect 45744 3528 45796 3534
rect 45744 3470 45796 3476
rect 45742 3088 45798 3097
rect 45742 3023 45744 3032
rect 45796 3023 45798 3032
rect 45744 2994 45796 3000
rect 45652 2984 45704 2990
rect 45650 2952 45652 2961
rect 45704 2952 45706 2961
rect 45650 2887 45706 2896
rect 45560 2440 45612 2446
rect 45560 2382 45612 2388
rect 45388 2332 45508 2360
rect 45192 2100 45244 2106
rect 45192 2042 45244 2048
rect 45388 800 45416 2332
rect 45848 1714 45876 3538
rect 45664 1686 45876 1714
rect 45664 800 45692 1686
rect 45940 800 45968 4558
rect 46032 3534 46060 52634
rect 46124 32502 46152 60998
rect 46676 60790 46704 63294
rect 47214 63200 47270 64000
rect 47950 63322 48006 64000
rect 47950 63294 48268 63322
rect 47950 63200 48006 63294
rect 47228 61198 47256 63200
rect 48240 61282 48268 63294
rect 48686 63200 48742 64000
rect 49422 63322 49478 64000
rect 49422 63294 49556 63322
rect 49422 63200 49478 63294
rect 48240 61254 48360 61282
rect 48332 61198 48360 61254
rect 48700 61198 48728 63200
rect 47216 61192 47268 61198
rect 47216 61134 47268 61140
rect 48320 61192 48372 61198
rect 48320 61134 48372 61140
rect 48688 61192 48740 61198
rect 48688 61134 48740 61140
rect 46940 61124 46992 61130
rect 46940 61066 46992 61072
rect 46664 60784 46716 60790
rect 46664 60726 46716 60732
rect 46756 60512 46808 60518
rect 46756 60454 46808 60460
rect 46296 37188 46348 37194
rect 46296 37130 46348 37136
rect 46308 36378 46336 37130
rect 46296 36372 46348 36378
rect 46296 36314 46348 36320
rect 46112 32496 46164 32502
rect 46112 32438 46164 32444
rect 46768 31890 46796 60454
rect 46952 54194 46980 61066
rect 47952 61056 48004 61062
rect 47952 60998 48004 61004
rect 48688 61056 48740 61062
rect 48688 60998 48740 61004
rect 47964 55282 47992 60998
rect 48700 56506 48728 60998
rect 49528 60722 49556 63294
rect 50158 63200 50214 64000
rect 50894 63322 50950 64000
rect 51630 63322 51686 64000
rect 50894 63294 51028 63322
rect 50894 63200 50950 63294
rect 50172 60790 50200 63200
rect 51000 62098 51028 63294
rect 51630 63294 52040 63322
rect 51630 63200 51686 63294
rect 51000 62070 51120 62098
rect 51092 61198 51120 62070
rect 52012 61198 52040 63294
rect 52366 63200 52422 64000
rect 53102 63322 53158 64000
rect 53838 63322 53894 64000
rect 54574 63322 54630 64000
rect 55310 63322 55366 64000
rect 56046 63322 56102 64000
rect 53102 63294 53236 63322
rect 53102 63200 53158 63294
rect 51080 61192 51132 61198
rect 51080 61134 51132 61140
rect 52000 61192 52052 61198
rect 52000 61134 52052 61140
rect 51172 61056 51224 61062
rect 51172 60998 51224 61004
rect 52092 61056 52144 61062
rect 52092 60998 52144 61004
rect 50294 60956 50602 60965
rect 50294 60954 50300 60956
rect 50356 60954 50380 60956
rect 50436 60954 50460 60956
rect 50516 60954 50540 60956
rect 50596 60954 50602 60956
rect 50356 60902 50358 60954
rect 50538 60902 50540 60954
rect 50294 60900 50300 60902
rect 50356 60900 50380 60902
rect 50436 60900 50460 60902
rect 50516 60900 50540 60902
rect 50596 60900 50602 60902
rect 50294 60891 50602 60900
rect 50160 60784 50212 60790
rect 50160 60726 50212 60732
rect 49516 60716 49568 60722
rect 49516 60658 49568 60664
rect 49700 60512 49752 60518
rect 49700 60454 49752 60460
rect 49792 60512 49844 60518
rect 49792 60454 49844 60460
rect 49608 60308 49660 60314
rect 49608 60250 49660 60256
rect 49620 57594 49648 60250
rect 49608 57588 49660 57594
rect 49608 57530 49660 57536
rect 48688 56500 48740 56506
rect 48688 56442 48740 56448
rect 47952 55276 48004 55282
rect 47952 55218 48004 55224
rect 46940 54188 46992 54194
rect 46940 54130 46992 54136
rect 47584 43784 47636 43790
rect 47584 43726 47636 43732
rect 46940 37392 46992 37398
rect 46940 37334 46992 37340
rect 46952 33318 46980 37334
rect 46940 33312 46992 33318
rect 46940 33254 46992 33260
rect 46756 31884 46808 31890
rect 46756 31826 46808 31832
rect 47596 31822 47624 43726
rect 49148 41608 49200 41614
rect 49148 41550 49200 41556
rect 48228 40520 48280 40526
rect 48228 40462 48280 40468
rect 48240 37466 48268 40462
rect 48228 37460 48280 37466
rect 48228 37402 48280 37408
rect 48688 36780 48740 36786
rect 48688 36722 48740 36728
rect 47676 35080 47728 35086
rect 47676 35022 47728 35028
rect 47584 31816 47636 31822
rect 47584 31758 47636 31764
rect 47216 29708 47268 29714
rect 47216 29650 47268 29656
rect 46112 29640 46164 29646
rect 46112 29582 46164 29588
rect 46124 20806 46152 29582
rect 47228 28966 47256 29650
rect 47216 28960 47268 28966
rect 47216 28902 47268 28908
rect 47584 28688 47636 28694
rect 47584 28630 47636 28636
rect 46480 26988 46532 26994
rect 46480 26930 46532 26936
rect 46216 24682 46428 24698
rect 46204 24676 46440 24682
rect 46256 24670 46388 24676
rect 46204 24618 46256 24624
rect 46388 24618 46440 24624
rect 46112 20800 46164 20806
rect 46112 20742 46164 20748
rect 46388 19984 46440 19990
rect 46388 19926 46440 19932
rect 46204 19848 46256 19854
rect 46204 19790 46256 19796
rect 46216 19514 46244 19790
rect 46400 19718 46428 19926
rect 46388 19712 46440 19718
rect 46388 19654 46440 19660
rect 46204 19508 46256 19514
rect 46204 19450 46256 19456
rect 46204 19236 46256 19242
rect 46204 19178 46256 19184
rect 46216 18970 46244 19178
rect 46204 18964 46256 18970
rect 46204 18906 46256 18912
rect 46204 17536 46256 17542
rect 46204 17478 46256 17484
rect 46216 17134 46244 17478
rect 46204 17128 46256 17134
rect 46204 17070 46256 17076
rect 46204 13252 46256 13258
rect 46204 13194 46256 13200
rect 46216 12986 46244 13194
rect 46204 12980 46256 12986
rect 46204 12922 46256 12928
rect 46204 4480 46256 4486
rect 46204 4422 46256 4428
rect 46216 4214 46244 4422
rect 46204 4208 46256 4214
rect 46204 4150 46256 4156
rect 46296 4208 46348 4214
rect 46296 4150 46348 4156
rect 46204 4072 46256 4078
rect 46204 4014 46256 4020
rect 46112 3732 46164 3738
rect 46112 3674 46164 3680
rect 46020 3528 46072 3534
rect 46020 3470 46072 3476
rect 46124 3058 46152 3674
rect 46216 3534 46244 4014
rect 46204 3528 46256 3534
rect 46204 3470 46256 3476
rect 46112 3052 46164 3058
rect 46112 2994 46164 3000
rect 46216 2582 46244 3470
rect 46204 2576 46256 2582
rect 46204 2518 46256 2524
rect 46308 2088 46336 4150
rect 46388 4004 46440 4010
rect 46388 3946 46440 3952
rect 46400 2854 46428 3946
rect 46388 2848 46440 2854
rect 46388 2790 46440 2796
rect 46492 2650 46520 26930
rect 47492 22024 47544 22030
rect 47492 21966 47544 21972
rect 47504 21078 47532 21966
rect 47492 21072 47544 21078
rect 47492 21014 47544 21020
rect 46848 20868 46900 20874
rect 46848 20810 46900 20816
rect 46860 15434 46888 20810
rect 47124 19780 47176 19786
rect 47124 19722 47176 19728
rect 47136 19446 47164 19722
rect 47124 19440 47176 19446
rect 47124 19382 47176 19388
rect 46848 15428 46900 15434
rect 46848 15370 46900 15376
rect 46860 12918 46888 15370
rect 46848 12912 46900 12918
rect 46848 12854 46900 12860
rect 47124 7200 47176 7206
rect 47124 7142 47176 7148
rect 47136 7002 47164 7142
rect 47124 6996 47176 7002
rect 47124 6938 47176 6944
rect 47596 4826 47624 28630
rect 47688 11762 47716 35022
rect 48044 32768 48096 32774
rect 48044 32710 48096 32716
rect 47952 28620 48004 28626
rect 47952 28562 48004 28568
rect 47860 23044 47912 23050
rect 47860 22986 47912 22992
rect 47872 22030 47900 22986
rect 47860 22024 47912 22030
rect 47860 21966 47912 21972
rect 47860 21888 47912 21894
rect 47860 21830 47912 21836
rect 47872 21729 47900 21830
rect 47858 21720 47914 21729
rect 47858 21655 47860 21664
rect 47912 21655 47914 21664
rect 47860 21626 47912 21632
rect 47872 21595 47900 21626
rect 47860 11824 47912 11830
rect 47860 11766 47912 11772
rect 47676 11756 47728 11762
rect 47676 11698 47728 11704
rect 47676 10804 47728 10810
rect 47676 10746 47728 10752
rect 47584 4820 47636 4826
rect 47584 4762 47636 4768
rect 46848 4684 46900 4690
rect 46848 4626 46900 4632
rect 46572 4616 46624 4622
rect 46572 4558 46624 4564
rect 46480 2644 46532 2650
rect 46480 2586 46532 2592
rect 46584 2360 46612 4558
rect 46860 4214 46888 4626
rect 47492 4616 47544 4622
rect 47492 4558 47544 4564
rect 46848 4208 46900 4214
rect 46848 4150 46900 4156
rect 47032 4208 47084 4214
rect 47032 4150 47084 4156
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 46676 2446 46704 3878
rect 46768 3602 46980 3618
rect 46768 3596 46992 3602
rect 46768 3590 46940 3596
rect 46664 2440 46716 2446
rect 46664 2382 46716 2388
rect 46216 2060 46336 2088
rect 46492 2332 46612 2360
rect 46216 800 46244 2060
rect 46492 800 46520 2332
rect 46768 800 46796 3590
rect 46940 3538 46992 3544
rect 46848 3528 46900 3534
rect 46848 3470 46900 3476
rect 46860 3233 46888 3470
rect 46846 3224 46902 3233
rect 46846 3159 46902 3168
rect 47044 800 47072 4150
rect 47122 3768 47178 3777
rect 47122 3703 47178 3712
rect 47136 3670 47164 3703
rect 47124 3664 47176 3670
rect 47124 3606 47176 3612
rect 47136 3466 47440 3482
rect 47124 3460 47452 3466
rect 47176 3454 47400 3460
rect 47124 3402 47176 3408
rect 47400 3402 47452 3408
rect 47308 3392 47360 3398
rect 47308 3334 47360 3340
rect 47320 2922 47348 3334
rect 47308 2916 47360 2922
rect 47308 2858 47360 2864
rect 47504 2394 47532 4558
rect 47688 4078 47716 10746
rect 47676 4072 47728 4078
rect 47676 4014 47728 4020
rect 47872 3942 47900 11766
rect 47860 3936 47912 3942
rect 47860 3878 47912 3884
rect 47584 3732 47636 3738
rect 47584 3674 47636 3680
rect 47596 3398 47624 3674
rect 47584 3392 47636 3398
rect 47584 3334 47636 3340
rect 47964 3194 47992 28562
rect 48056 27062 48084 32710
rect 48044 27056 48096 27062
rect 48044 26998 48096 27004
rect 48136 23112 48188 23118
rect 48136 23054 48188 23060
rect 48148 22710 48176 23054
rect 48136 22704 48188 22710
rect 48136 22646 48188 22652
rect 48136 22432 48188 22438
rect 48136 22374 48188 22380
rect 48148 20942 48176 22374
rect 48504 22024 48556 22030
rect 48504 21966 48556 21972
rect 48516 21554 48544 21966
rect 48504 21548 48556 21554
rect 48504 21490 48556 21496
rect 48228 21004 48280 21010
rect 48228 20946 48280 20952
rect 48136 20936 48188 20942
rect 48136 20878 48188 20884
rect 48044 20528 48096 20534
rect 48044 20470 48096 20476
rect 48056 3738 48084 20470
rect 48148 16182 48176 20878
rect 48240 20534 48268 20946
rect 48320 20800 48372 20806
rect 48320 20742 48372 20748
rect 48332 20602 48360 20742
rect 48320 20596 48372 20602
rect 48320 20538 48372 20544
rect 48228 20528 48280 20534
rect 48228 20470 48280 20476
rect 48136 16176 48188 16182
rect 48136 16118 48188 16124
rect 48148 15706 48176 16118
rect 48136 15700 48188 15706
rect 48136 15642 48188 15648
rect 48044 3732 48096 3738
rect 48044 3674 48096 3680
rect 48700 3194 48728 36722
rect 48964 33312 49016 33318
rect 48964 33254 49016 33260
rect 48872 22636 48924 22642
rect 48872 22578 48924 22584
rect 48884 22098 48912 22578
rect 48872 22092 48924 22098
rect 48872 22034 48924 22040
rect 48780 21888 48832 21894
rect 48780 21830 48832 21836
rect 48792 21350 48820 21830
rect 48780 21344 48832 21350
rect 48780 21286 48832 21292
rect 47952 3188 48004 3194
rect 47952 3130 48004 3136
rect 48688 3188 48740 3194
rect 48688 3130 48740 3136
rect 48412 3052 48464 3058
rect 48412 2994 48464 3000
rect 48688 3052 48740 3058
rect 48688 2994 48740 3000
rect 48136 2984 48188 2990
rect 48136 2926 48188 2932
rect 48044 2440 48096 2446
rect 47320 2366 47532 2394
rect 47950 2408 48006 2417
rect 47584 2372 47636 2378
rect 47320 800 47348 2366
rect 48044 2382 48096 2388
rect 47950 2343 48006 2352
rect 47584 2314 47636 2320
rect 47596 800 47624 2314
rect 47964 2310 47992 2343
rect 47952 2304 48004 2310
rect 47952 2246 48004 2252
rect 48056 1306 48084 2382
rect 47872 1278 48084 1306
rect 47872 800 47900 1278
rect 48148 800 48176 2926
rect 48424 800 48452 2994
rect 48700 800 48728 2994
rect 48976 2514 49004 33254
rect 49056 29300 49108 29306
rect 49056 29242 49108 29248
rect 49068 2650 49096 29242
rect 49160 22778 49188 41550
rect 49712 32298 49740 60454
rect 49804 57866 49832 60454
rect 50294 59868 50602 59877
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59803 50602 59812
rect 50294 58780 50602 58789
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58715 50602 58724
rect 50068 57928 50120 57934
rect 50068 57870 50120 57876
rect 49792 57860 49844 57866
rect 49792 57802 49844 57808
rect 50080 56166 50108 57870
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 51080 57520 51132 57526
rect 51080 57462 51132 57468
rect 51092 57322 51120 57462
rect 51080 57316 51132 57322
rect 51080 57258 51132 57264
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 50068 56160 50120 56166
rect 50068 56102 50120 56108
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 49884 35216 49936 35222
rect 49884 35158 49936 35164
rect 49700 32292 49752 32298
rect 49700 32234 49752 32240
rect 49240 31952 49292 31958
rect 49240 31894 49292 31900
rect 49148 22772 49200 22778
rect 49148 22714 49200 22720
rect 49160 22166 49188 22714
rect 49148 22160 49200 22166
rect 49148 22102 49200 22108
rect 49252 11014 49280 31894
rect 49792 26920 49844 26926
rect 49792 26862 49844 26868
rect 49700 20460 49752 20466
rect 49700 20402 49752 20408
rect 49712 19417 49740 20402
rect 49698 19408 49754 19417
rect 49698 19343 49754 19352
rect 49240 11008 49292 11014
rect 49240 10950 49292 10956
rect 49240 3460 49292 3466
rect 49240 3402 49292 3408
rect 49516 3460 49568 3466
rect 49516 3402 49568 3408
rect 49056 2644 49108 2650
rect 49056 2586 49108 2592
rect 48964 2508 49016 2514
rect 48964 2450 49016 2456
rect 48964 2372 49016 2378
rect 48964 2314 49016 2320
rect 48976 800 49004 2314
rect 49252 800 49280 3402
rect 49528 800 49556 3402
rect 49804 3194 49832 26862
rect 49896 3738 49924 35158
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50988 33924 51040 33930
rect 50988 33866 51040 33872
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50068 24608 50120 24614
rect 50068 24550 50120 24556
rect 50080 24206 50108 24550
rect 50068 24200 50120 24206
rect 50068 24142 50120 24148
rect 50896 24200 50948 24206
rect 50896 24142 50948 24148
rect 49976 23044 50028 23050
rect 49976 22986 50028 22992
rect 49988 20466 50016 22986
rect 49976 20460 50028 20466
rect 49976 20402 50028 20408
rect 49988 19854 50016 20402
rect 49976 19848 50028 19854
rect 49976 19790 50028 19796
rect 49988 19378 50016 19790
rect 49976 19372 50028 19378
rect 49976 19314 50028 19320
rect 50080 9518 50108 24142
rect 50804 24132 50856 24138
rect 50724 24092 50804 24120
rect 50620 24064 50672 24070
rect 50620 24006 50672 24012
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50632 23730 50660 24006
rect 50620 23724 50672 23730
rect 50620 23666 50672 23672
rect 50724 23118 50752 24092
rect 50804 24074 50856 24080
rect 50908 23322 50936 24142
rect 50896 23316 50948 23322
rect 50896 23258 50948 23264
rect 50712 23112 50764 23118
rect 50712 23054 50764 23060
rect 50724 22982 50752 23054
rect 50712 22976 50764 22982
rect 50712 22918 50764 22924
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50160 21548 50212 21554
rect 50160 21490 50212 21496
rect 50172 20602 50200 21490
rect 50436 21344 50488 21350
rect 50436 21286 50488 21292
rect 50448 20874 50476 21286
rect 50436 20868 50488 20874
rect 50436 20810 50488 20816
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50160 20596 50212 20602
rect 50160 20538 50212 20544
rect 50724 20466 50752 22918
rect 50712 20460 50764 20466
rect 50712 20402 50764 20408
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50712 13932 50764 13938
rect 50712 13874 50764 13880
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50068 9512 50120 9518
rect 50068 9454 50120 9460
rect 50080 8974 50108 9454
rect 50068 8968 50120 8974
rect 50068 8910 50120 8916
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50160 7812 50212 7818
rect 50160 7754 50212 7760
rect 50172 7478 50200 7754
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50160 7472 50212 7478
rect 50160 7414 50212 7420
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 49884 3732 49936 3738
rect 49884 3674 49936 3680
rect 50620 3528 50672 3534
rect 50620 3470 50672 3476
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 49792 3188 49844 3194
rect 49792 3130 49844 3136
rect 49792 2984 49844 2990
rect 49792 2926 49844 2932
rect 49804 800 49832 2926
rect 50068 2916 50120 2922
rect 50068 2858 50120 2864
rect 50080 800 50108 2858
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50344 1420 50396 1426
rect 50344 1362 50396 1368
rect 50356 800 50384 1362
rect 50632 800 50660 3470
rect 50724 1358 50752 13874
rect 50804 9512 50856 9518
rect 50804 9454 50856 9460
rect 50816 3602 50844 9454
rect 50896 3664 50948 3670
rect 50894 3632 50896 3641
rect 50948 3632 50950 3641
rect 50804 3596 50856 3602
rect 50894 3567 50950 3576
rect 50804 3538 50856 3544
rect 50896 3460 50948 3466
rect 50896 3402 50948 3408
rect 50712 1352 50764 1358
rect 50712 1294 50764 1300
rect 50908 800 50936 3402
rect 51000 3194 51028 33866
rect 51184 24818 51212 60998
rect 51724 35080 51776 35086
rect 51724 35022 51776 35028
rect 51172 24812 51224 24818
rect 51172 24754 51224 24760
rect 51540 24268 51592 24274
rect 51540 24210 51592 24216
rect 51356 24132 51408 24138
rect 51552 24120 51580 24210
rect 51632 24200 51684 24206
rect 51632 24142 51684 24148
rect 51408 24092 51580 24120
rect 51356 24074 51408 24080
rect 51644 22098 51672 24142
rect 51736 23594 51764 35022
rect 51816 24744 51868 24750
rect 51816 24686 51868 24692
rect 51828 24138 51856 24686
rect 51816 24132 51868 24138
rect 51816 24074 51868 24080
rect 51724 23588 51776 23594
rect 51724 23530 51776 23536
rect 51736 23050 51764 23530
rect 51724 23044 51776 23050
rect 51724 22986 51776 22992
rect 51632 22092 51684 22098
rect 51632 22034 51684 22040
rect 51644 21690 51672 22034
rect 51724 22024 51776 22030
rect 51724 21966 51776 21972
rect 51632 21684 51684 21690
rect 51632 21626 51684 21632
rect 51736 21146 51764 21966
rect 51724 21140 51776 21146
rect 51724 21082 51776 21088
rect 51736 20398 51764 21082
rect 51724 20392 51776 20398
rect 51724 20334 51776 20340
rect 51828 20262 51856 24074
rect 52000 23656 52052 23662
rect 52000 23598 52052 23604
rect 52012 21486 52040 23598
rect 52000 21480 52052 21486
rect 52000 21422 52052 21428
rect 51816 20256 51868 20262
rect 51816 20198 51868 20204
rect 52012 19310 52040 21422
rect 52104 20330 52132 60998
rect 52380 60772 52408 63200
rect 53208 61198 53236 63294
rect 53838 63294 54248 63322
rect 53838 63200 53894 63294
rect 54220 61198 54248 63294
rect 54574 63294 54800 63322
rect 54574 63200 54630 63294
rect 53196 61192 53248 61198
rect 53196 61134 53248 61140
rect 54208 61192 54260 61198
rect 54208 61134 54260 61140
rect 54392 61124 54444 61130
rect 54392 61066 54444 61072
rect 52460 60784 52512 60790
rect 52380 60744 52460 60772
rect 52460 60726 52512 60732
rect 53104 60512 53156 60518
rect 53104 60454 53156 60460
rect 53116 59090 53144 60454
rect 53104 59084 53156 59090
rect 53104 59026 53156 59032
rect 54024 57860 54076 57866
rect 54024 57802 54076 57808
rect 54036 57458 54064 57802
rect 54024 57452 54076 57458
rect 54024 57394 54076 57400
rect 53932 57384 53984 57390
rect 53932 57326 53984 57332
rect 53472 56704 53524 56710
rect 53472 56646 53524 56652
rect 52276 31272 52328 31278
rect 52276 31214 52328 31220
rect 52092 20324 52144 20330
rect 52092 20266 52144 20272
rect 52184 19712 52236 19718
rect 52184 19654 52236 19660
rect 52196 19378 52224 19654
rect 52184 19372 52236 19378
rect 52184 19314 52236 19320
rect 52000 19304 52052 19310
rect 52000 19246 52052 19252
rect 52012 16658 52040 19246
rect 52000 16652 52052 16658
rect 52000 16594 52052 16600
rect 51448 11756 51500 11762
rect 51448 11698 51500 11704
rect 51264 11008 51316 11014
rect 51264 10950 51316 10956
rect 51276 3738 51304 10950
rect 51264 3732 51316 3738
rect 51264 3674 51316 3680
rect 50988 3188 51040 3194
rect 50988 3130 51040 3136
rect 51356 2848 51408 2854
rect 51356 2790 51408 2796
rect 51368 2582 51396 2790
rect 51460 2650 51488 11698
rect 52288 6914 52316 31214
rect 53012 31204 53064 31210
rect 53012 31146 53064 31152
rect 52920 31136 52972 31142
rect 52920 31078 52972 31084
rect 52736 28960 52788 28966
rect 52736 28902 52788 28908
rect 52552 24200 52604 24206
rect 52552 24142 52604 24148
rect 52564 23798 52592 24142
rect 52552 23792 52604 23798
rect 52552 23734 52604 23740
rect 52368 20936 52420 20942
rect 52368 20878 52420 20884
rect 52380 20466 52408 20878
rect 52368 20460 52420 20466
rect 52368 20402 52420 20408
rect 52552 20392 52604 20398
rect 52552 20334 52604 20340
rect 52368 20256 52420 20262
rect 52368 20198 52420 20204
rect 52380 19786 52408 20198
rect 52564 19786 52592 20334
rect 52368 19780 52420 19786
rect 52368 19722 52420 19728
rect 52552 19780 52604 19786
rect 52552 19722 52604 19728
rect 52460 19440 52512 19446
rect 52460 19382 52512 19388
rect 52472 18426 52500 19382
rect 52460 18420 52512 18426
rect 52460 18362 52512 18368
rect 52196 6886 52316 6914
rect 51724 3528 51776 3534
rect 51724 3470 51776 3476
rect 51540 3120 51592 3126
rect 51540 3062 51592 3068
rect 51448 2644 51500 2650
rect 51448 2586 51500 2592
rect 51356 2576 51408 2582
rect 51356 2518 51408 2524
rect 51172 2440 51224 2446
rect 51172 2382 51224 2388
rect 51184 800 51212 2382
rect 51356 2372 51408 2378
rect 51356 2314 51408 2320
rect 51368 1426 51396 2314
rect 51552 1578 51580 3062
rect 51460 1550 51580 1578
rect 51356 1420 51408 1426
rect 51356 1362 51408 1368
rect 51460 800 51488 1550
rect 51736 800 51764 3470
rect 52196 3194 52224 6886
rect 52748 3738 52776 28902
rect 52932 3738 52960 31078
rect 53024 16574 53052 31146
rect 53484 29782 53512 56646
rect 53944 31686 53972 57326
rect 54036 57254 54064 57394
rect 54024 57248 54076 57254
rect 54024 57190 54076 57196
rect 54036 56846 54064 57190
rect 54404 56846 54432 61066
rect 54772 60790 54800 63294
rect 55310 63294 55536 63322
rect 55310 63200 55366 63294
rect 55508 60790 55536 63294
rect 56046 63294 56272 63322
rect 56046 63200 56102 63294
rect 56046 62656 56102 62665
rect 56046 62591 56102 62600
rect 54760 60784 54812 60790
rect 54760 60726 54812 60732
rect 55496 60784 55548 60790
rect 55496 60726 55548 60732
rect 54852 60512 54904 60518
rect 54852 60454 54904 60460
rect 55588 60512 55640 60518
rect 55588 60454 55640 60460
rect 54484 60240 54536 60246
rect 54484 60182 54536 60188
rect 54024 56840 54076 56846
rect 54024 56782 54076 56788
rect 54392 56840 54444 56846
rect 54392 56782 54444 56788
rect 54496 44878 54524 60182
rect 54760 59968 54812 59974
rect 54760 59910 54812 59916
rect 54576 57928 54628 57934
rect 54576 57870 54628 57876
rect 54588 57594 54616 57870
rect 54772 57866 54800 59910
rect 54760 57860 54812 57866
rect 54760 57802 54812 57808
rect 54576 57588 54628 57594
rect 54576 57530 54628 57536
rect 54588 56846 54616 57530
rect 54864 57458 54892 60454
rect 55220 58336 55272 58342
rect 55220 58278 55272 58284
rect 55232 57934 55260 58278
rect 55220 57928 55272 57934
rect 55220 57870 55272 57876
rect 54852 57452 54904 57458
rect 54852 57394 54904 57400
rect 55600 57254 55628 60454
rect 56060 60042 56088 62591
rect 56138 62112 56194 62121
rect 56138 62047 56194 62056
rect 56152 61198 56180 62047
rect 56140 61192 56192 61198
rect 56140 61134 56192 61140
rect 56138 61024 56194 61033
rect 56138 60959 56194 60968
rect 56152 60722 56180 60959
rect 56140 60716 56192 60722
rect 56140 60658 56192 60664
rect 56244 60110 56272 63294
rect 56782 63200 56838 64000
rect 57518 63200 57574 64000
rect 58254 63200 58310 64000
rect 58990 63322 59046 64000
rect 58728 63294 59046 63322
rect 56506 61568 56562 61577
rect 56506 61503 56562 61512
rect 56416 61124 56468 61130
rect 56416 61066 56468 61072
rect 56324 60648 56376 60654
rect 56324 60590 56376 60596
rect 56232 60104 56284 60110
rect 56232 60046 56284 60052
rect 56048 60036 56100 60042
rect 56048 59978 56100 59984
rect 55588 57248 55640 57254
rect 55588 57190 55640 57196
rect 54576 56840 54628 56846
rect 54576 56782 54628 56788
rect 54484 44872 54536 44878
rect 54484 44814 54536 44820
rect 55956 44872 56008 44878
rect 55956 44814 56008 44820
rect 55968 31754 55996 44814
rect 56048 39840 56100 39846
rect 56048 39782 56100 39788
rect 55876 31726 55996 31754
rect 53932 31680 53984 31686
rect 53932 31622 53984 31628
rect 53472 29776 53524 29782
rect 53472 29718 53524 29724
rect 54760 28416 54812 28422
rect 54760 28358 54812 28364
rect 53840 25220 53892 25226
rect 53840 25162 53892 25168
rect 53288 24132 53340 24138
rect 53288 24074 53340 24080
rect 53104 24064 53156 24070
rect 53104 24006 53156 24012
rect 53116 23730 53144 24006
rect 53300 23730 53328 24074
rect 53104 23724 53156 23730
rect 53104 23666 53156 23672
rect 53288 23724 53340 23730
rect 53288 23666 53340 23672
rect 53852 23254 53880 25162
rect 54116 24744 54168 24750
rect 54116 24686 54168 24692
rect 54024 24132 54076 24138
rect 54024 24074 54076 24080
rect 54036 23526 54064 24074
rect 54024 23520 54076 23526
rect 54024 23462 54076 23468
rect 53840 23248 53892 23254
rect 53840 23190 53892 23196
rect 54128 23118 54156 24686
rect 54484 24608 54536 24614
rect 54484 24550 54536 24556
rect 54496 24274 54524 24550
rect 54484 24268 54536 24274
rect 54484 24210 54536 24216
rect 54668 24200 54720 24206
rect 54668 24142 54720 24148
rect 54392 23520 54444 23526
rect 54392 23462 54444 23468
rect 54404 23186 54432 23462
rect 54680 23322 54708 24142
rect 54668 23316 54720 23322
rect 54668 23258 54720 23264
rect 54392 23180 54444 23186
rect 54392 23122 54444 23128
rect 53932 23112 53984 23118
rect 53932 23054 53984 23060
rect 54116 23112 54168 23118
rect 54116 23054 54168 23060
rect 53944 22982 53972 23054
rect 53380 22976 53432 22982
rect 53380 22918 53432 22924
rect 53932 22976 53984 22982
rect 53932 22918 53984 22924
rect 53392 22234 53420 22918
rect 53380 22228 53432 22234
rect 53380 22170 53432 22176
rect 53944 22098 53972 22918
rect 53932 22092 53984 22098
rect 53932 22034 53984 22040
rect 53944 20806 53972 22034
rect 53932 20800 53984 20806
rect 53932 20742 53984 20748
rect 54300 20596 54352 20602
rect 54300 20538 54352 20544
rect 53196 20460 53248 20466
rect 53196 20402 53248 20408
rect 53208 19514 53236 20402
rect 54312 20262 54340 20538
rect 54300 20256 54352 20262
rect 54300 20198 54352 20204
rect 54312 19922 54340 20198
rect 54300 19916 54352 19922
rect 54300 19858 54352 19864
rect 53196 19508 53248 19514
rect 53196 19450 53248 19456
rect 53196 19372 53248 19378
rect 53196 19314 53248 19320
rect 53024 16546 53144 16574
rect 52736 3732 52788 3738
rect 52736 3674 52788 3680
rect 52920 3732 52972 3738
rect 52920 3674 52972 3680
rect 52276 3460 52328 3466
rect 52276 3402 52328 3408
rect 52184 3188 52236 3194
rect 52184 3130 52236 3136
rect 52000 3052 52052 3058
rect 52000 2994 52052 3000
rect 52012 800 52040 2994
rect 52288 800 52316 3402
rect 52460 3188 52512 3194
rect 52460 3130 52512 3136
rect 52472 3097 52500 3130
rect 52458 3088 52514 3097
rect 52458 3023 52514 3032
rect 52552 2984 52604 2990
rect 52552 2926 52604 2932
rect 52564 800 52592 2926
rect 53116 2650 53144 16546
rect 53208 3670 53236 19314
rect 53840 10056 53892 10062
rect 53840 9998 53892 10004
rect 53852 9382 53880 9998
rect 53840 9376 53892 9382
rect 53840 9318 53892 9324
rect 53564 7404 53616 7410
rect 53564 7346 53616 7352
rect 53576 3738 53604 7346
rect 53932 4004 53984 4010
rect 53932 3946 53984 3952
rect 53564 3732 53616 3738
rect 53564 3674 53616 3680
rect 53196 3664 53248 3670
rect 53196 3606 53248 3612
rect 53196 3460 53248 3466
rect 53196 3402 53248 3408
rect 53104 2644 53156 2650
rect 53104 2586 53156 2592
rect 52828 2304 52880 2310
rect 52828 2246 52880 2252
rect 52840 800 52868 2246
rect 53208 898 53236 3402
rect 53944 3194 53972 3946
rect 54668 3392 54720 3398
rect 54668 3334 54720 3340
rect 53932 3188 53984 3194
rect 53932 3130 53984 3136
rect 53380 3120 53432 3126
rect 53380 3062 53432 3068
rect 53116 870 53236 898
rect 53116 800 53144 870
rect 53392 800 53420 3062
rect 54680 3058 54708 3334
rect 54668 3052 54720 3058
rect 54668 2994 54720 3000
rect 54772 2514 54800 28358
rect 55312 28212 55364 28218
rect 55312 28154 55364 28160
rect 55324 24818 55352 28154
rect 55496 25492 55548 25498
rect 55496 25434 55548 25440
rect 55588 25492 55640 25498
rect 55588 25434 55640 25440
rect 55508 24818 55536 25434
rect 55600 24886 55628 25434
rect 55772 25288 55824 25294
rect 55772 25230 55824 25236
rect 55588 24880 55640 24886
rect 55588 24822 55640 24828
rect 55312 24812 55364 24818
rect 55312 24754 55364 24760
rect 55496 24812 55548 24818
rect 55496 24754 55548 24760
rect 55128 24744 55180 24750
rect 55128 24686 55180 24692
rect 55036 24676 55088 24682
rect 55036 24618 55088 24624
rect 55048 24138 55076 24618
rect 55036 24132 55088 24138
rect 55036 24074 55088 24080
rect 54852 24064 54904 24070
rect 54852 24006 54904 24012
rect 54864 23730 54892 24006
rect 54852 23724 54904 23730
rect 54852 23666 54904 23672
rect 55140 22982 55168 24686
rect 55784 24614 55812 25230
rect 55772 24608 55824 24614
rect 55772 24550 55824 24556
rect 55876 24342 55904 31726
rect 56060 28218 56088 39782
rect 56336 38010 56364 60590
rect 56324 38004 56376 38010
rect 56324 37946 56376 37952
rect 56428 34542 56456 61066
rect 56520 58954 56548 61503
rect 56796 61266 56824 63200
rect 56784 61260 56836 61266
rect 56784 61202 56836 61208
rect 57532 61198 57560 63200
rect 57520 61192 57572 61198
rect 57520 61134 57572 61140
rect 56876 61056 56928 61062
rect 56876 60998 56928 61004
rect 58164 61056 58216 61062
rect 58164 60998 58216 61004
rect 56508 58948 56560 58954
rect 56508 58890 56560 58896
rect 56888 51074 56916 60998
rect 57796 60784 57848 60790
rect 57796 60726 57848 60732
rect 57060 60512 57112 60518
rect 57060 60454 57112 60460
rect 57334 60480 57390 60489
rect 56796 51046 56916 51074
rect 56796 45898 56824 51046
rect 56876 48136 56928 48142
rect 56876 48078 56928 48084
rect 56784 45892 56836 45898
rect 56784 45834 56836 45840
rect 56416 34536 56468 34542
rect 56416 34478 56468 34484
rect 56888 31754 56916 48078
rect 57072 47598 57100 60454
rect 57334 60415 57390 60424
rect 57244 59560 57296 59566
rect 57244 59502 57296 59508
rect 57060 47592 57112 47598
rect 57060 47534 57112 47540
rect 57256 45554 57284 59502
rect 57348 59022 57376 60415
rect 57808 59401 57836 60726
rect 57980 60036 58032 60042
rect 57980 59978 58032 59984
rect 57992 59945 58020 59978
rect 57978 59936 58034 59945
rect 57978 59871 58034 59880
rect 57888 59628 57940 59634
rect 57888 59570 57940 59576
rect 57794 59392 57850 59401
rect 57794 59327 57850 59336
rect 57336 59016 57388 59022
rect 57336 58958 57388 58964
rect 57336 58880 57388 58886
rect 57900 58857 57928 59570
rect 58072 58880 58124 58886
rect 57336 58822 57388 58828
rect 57886 58848 57942 58857
rect 57348 58478 57376 58822
rect 58072 58822 58124 58828
rect 57886 58783 57942 58792
rect 57336 58472 57388 58478
rect 57336 58414 57388 58420
rect 57796 50312 57848 50318
rect 57796 50254 57848 50260
rect 57336 48068 57388 48074
rect 57336 48010 57388 48016
rect 57348 47977 57376 48010
rect 57334 47968 57390 47977
rect 57334 47903 57390 47912
rect 57612 47048 57664 47054
rect 57612 46990 57664 46996
rect 57164 45526 57284 45554
rect 56968 42696 57020 42702
rect 56968 42638 57020 42644
rect 56980 42537 57008 42638
rect 56966 42528 57022 42537
rect 56966 42463 57022 42472
rect 57060 39364 57112 39370
rect 57060 39306 57112 39312
rect 57072 39273 57100 39306
rect 57058 39264 57114 39273
rect 57058 39199 57114 39208
rect 57164 34950 57192 45526
rect 57244 44804 57296 44810
rect 57244 44746 57296 44752
rect 57256 44713 57284 44746
rect 57242 44704 57298 44713
rect 57242 44639 57298 44648
rect 57244 41540 57296 41546
rect 57244 41482 57296 41488
rect 57256 41449 57284 41482
rect 57242 41440 57298 41449
rect 57242 41375 57298 41384
rect 57244 38276 57296 38282
rect 57244 38218 57296 38224
rect 57256 38185 57284 38218
rect 57242 38176 57298 38185
rect 57242 38111 57298 38120
rect 57152 34944 57204 34950
rect 57152 34886 57204 34892
rect 57520 32904 57572 32910
rect 57520 32846 57572 32852
rect 57060 32836 57112 32842
rect 57060 32778 57112 32784
rect 57072 32745 57100 32778
rect 57058 32736 57114 32745
rect 57058 32671 57114 32680
rect 57428 31816 57480 31822
rect 57428 31758 57480 31764
rect 56888 31726 57008 31754
rect 56048 28212 56100 28218
rect 56048 28154 56100 28160
rect 56048 25288 56100 25294
rect 56048 25230 56100 25236
rect 56876 25288 56928 25294
rect 56876 25230 56928 25236
rect 56060 24954 56088 25230
rect 56324 25152 56376 25158
rect 56324 25094 56376 25100
rect 56048 24948 56100 24954
rect 56048 24890 56100 24896
rect 56232 24812 56284 24818
rect 56232 24754 56284 24760
rect 56244 24682 56272 24754
rect 56232 24676 56284 24682
rect 56232 24618 56284 24624
rect 55864 24336 55916 24342
rect 55864 24278 55916 24284
rect 56048 24200 56100 24206
rect 56048 24142 56100 24148
rect 56060 23798 56088 24142
rect 56048 23792 56100 23798
rect 56048 23734 56100 23740
rect 56048 23112 56100 23118
rect 56048 23054 56100 23060
rect 56244 23100 56272 24618
rect 56336 24206 56364 25094
rect 56888 24954 56916 25230
rect 56876 24948 56928 24954
rect 56876 24890 56928 24896
rect 56508 24812 56560 24818
rect 56508 24754 56560 24760
rect 56692 24812 56744 24818
rect 56692 24754 56744 24760
rect 56876 24812 56928 24818
rect 56876 24754 56928 24760
rect 56324 24200 56376 24206
rect 56324 24142 56376 24148
rect 56520 23866 56548 24754
rect 56704 24614 56732 24754
rect 56888 24682 56916 24754
rect 56876 24676 56928 24682
rect 56876 24618 56928 24624
rect 56692 24608 56744 24614
rect 56692 24550 56744 24556
rect 56508 23860 56560 23866
rect 56508 23802 56560 23808
rect 56876 23792 56928 23798
rect 56876 23734 56928 23740
rect 56416 23724 56468 23730
rect 56416 23666 56468 23672
rect 56324 23112 56376 23118
rect 56244 23072 56324 23100
rect 55956 23044 56008 23050
rect 55956 22986 56008 22992
rect 55128 22976 55180 22982
rect 55128 22918 55180 22924
rect 55968 21418 55996 22986
rect 55956 21412 56008 21418
rect 55956 21354 56008 21360
rect 56060 20942 56088 23054
rect 56244 21842 56272 23072
rect 56324 23054 56376 23060
rect 56428 22506 56456 23666
rect 56888 23186 56916 23734
rect 56508 23180 56560 23186
rect 56508 23122 56560 23128
rect 56876 23180 56928 23186
rect 56876 23122 56928 23128
rect 56520 22642 56548 23122
rect 56508 22636 56560 22642
rect 56508 22578 56560 22584
rect 56784 22636 56836 22642
rect 56784 22578 56836 22584
rect 56416 22500 56468 22506
rect 56416 22442 56468 22448
rect 56324 22432 56376 22438
rect 56324 22374 56376 22380
rect 56336 22001 56364 22374
rect 56322 21992 56378 22001
rect 56322 21927 56378 21936
rect 56244 21814 56364 21842
rect 56232 21548 56284 21554
rect 56232 21490 56284 21496
rect 56244 21010 56272 21490
rect 56232 21004 56284 21010
rect 56232 20946 56284 20952
rect 56048 20936 56100 20942
rect 56048 20878 56100 20884
rect 56140 20868 56192 20874
rect 56140 20810 56192 20816
rect 56048 16516 56100 16522
rect 56048 16458 56100 16464
rect 56060 15502 56088 16458
rect 56152 16182 56180 20810
rect 56336 19786 56364 21814
rect 56796 21554 56824 22578
rect 56784 21548 56836 21554
rect 56784 21490 56836 21496
rect 56416 20868 56468 20874
rect 56416 20810 56468 20816
rect 56324 19780 56376 19786
rect 56324 19722 56376 19728
rect 56140 16176 56192 16182
rect 56140 16118 56192 16124
rect 56048 15496 56100 15502
rect 56048 15438 56100 15444
rect 56428 12782 56456 20810
rect 56796 20262 56824 21490
rect 56888 21010 56916 23122
rect 56980 22094 57008 31726
rect 57060 29572 57112 29578
rect 57060 29514 57112 29520
rect 57072 29481 57100 29514
rect 57152 29504 57204 29510
rect 57058 29472 57114 29481
rect 57152 29446 57204 29452
rect 57058 29407 57114 29416
rect 57164 29170 57192 29446
rect 57152 29164 57204 29170
rect 57152 29106 57204 29112
rect 57152 25152 57204 25158
rect 57152 25094 57204 25100
rect 57164 23118 57192 25094
rect 57440 24750 57468 31758
rect 57428 24744 57480 24750
rect 57428 24686 57480 24692
rect 57440 24342 57468 24686
rect 57428 24336 57480 24342
rect 57428 24278 57480 24284
rect 57532 23866 57560 32846
rect 57520 23860 57572 23866
rect 57520 23802 57572 23808
rect 57152 23112 57204 23118
rect 57152 23054 57204 23060
rect 57532 23050 57560 23802
rect 57520 23044 57572 23050
rect 57520 22986 57572 22992
rect 56980 22066 57100 22094
rect 56968 21344 57020 21350
rect 56968 21286 57020 21292
rect 56876 21004 56928 21010
rect 56876 20946 56928 20952
rect 56980 20942 57008 21286
rect 56968 20936 57020 20942
rect 56968 20878 57020 20884
rect 56784 20256 56836 20262
rect 56784 20198 56836 20204
rect 56508 19780 56560 19786
rect 56508 19722 56560 19728
rect 56520 18358 56548 19722
rect 56796 19378 56824 20198
rect 57072 19938 57100 22066
rect 57152 21548 57204 21554
rect 57152 21490 57204 21496
rect 57164 21321 57192 21490
rect 57244 21344 57296 21350
rect 57150 21312 57206 21321
rect 57244 21286 57296 21292
rect 57150 21247 57206 21256
rect 57072 19910 57192 19938
rect 57060 19780 57112 19786
rect 57060 19722 57112 19728
rect 57072 19689 57100 19722
rect 57058 19680 57114 19689
rect 57058 19615 57114 19624
rect 56784 19372 56836 19378
rect 56784 19314 56836 19320
rect 56796 18426 56824 19314
rect 56968 19168 57020 19174
rect 56968 19110 57020 19116
rect 56980 18766 57008 19110
rect 57164 18970 57192 19910
rect 57152 18964 57204 18970
rect 57152 18906 57204 18912
rect 57256 18873 57284 21286
rect 57624 20602 57652 46990
rect 57704 37256 57756 37262
rect 57704 37198 57756 37204
rect 57716 21162 57744 37198
rect 57808 23526 57836 50254
rect 57888 50176 57940 50182
rect 57888 50118 57940 50124
rect 57900 49609 57928 50118
rect 57886 49600 57942 49609
rect 57886 49535 57942 49544
rect 57980 49156 58032 49162
rect 57980 49098 58032 49104
rect 57992 49065 58020 49098
rect 57978 49056 58034 49065
rect 57978 48991 58034 49000
rect 57980 48068 58032 48074
rect 57980 48010 58032 48016
rect 57992 47433 58020 48010
rect 57978 47424 58034 47433
rect 57978 47359 58034 47368
rect 57888 46912 57940 46918
rect 57888 46854 57940 46860
rect 57900 46345 57928 46854
rect 57886 46336 57942 46345
rect 57886 46271 57942 46280
rect 57980 45892 58032 45898
rect 57980 45834 58032 45840
rect 57992 45801 58020 45834
rect 57978 45792 58034 45801
rect 57978 45727 58034 45736
rect 57888 44804 57940 44810
rect 57888 44746 57940 44752
rect 57900 44169 57928 44746
rect 57886 44160 57942 44169
rect 57886 44095 57942 44104
rect 57888 42696 57940 42702
rect 57888 42638 57940 42644
rect 57900 41993 57928 42638
rect 57886 41984 57942 41993
rect 57886 41919 57942 41928
rect 57888 41540 57940 41546
rect 57888 41482 57940 41488
rect 57900 40905 57928 41482
rect 57886 40896 57942 40905
rect 57886 40831 57942 40840
rect 57888 40384 57940 40390
rect 57888 40326 57940 40332
rect 57900 39817 57928 40326
rect 57886 39808 57942 39817
rect 57886 39743 57942 39752
rect 57980 39364 58032 39370
rect 57980 39306 58032 39312
rect 57992 38729 58020 39306
rect 57978 38720 58034 38729
rect 57978 38655 58034 38664
rect 57888 38344 57940 38350
rect 57888 38286 57940 38292
rect 57900 37641 57928 38286
rect 57886 37632 57942 37641
rect 57886 37567 57942 37576
rect 57980 36100 58032 36106
rect 57980 36042 58032 36048
rect 57992 36009 58020 36042
rect 57978 36000 58034 36009
rect 57978 35935 58034 35944
rect 58084 35086 58112 58822
rect 58176 58682 58204 60998
rect 58268 60858 58296 63200
rect 58256 60852 58308 60858
rect 58256 60794 58308 60800
rect 58256 60512 58308 60518
rect 58256 60454 58308 60460
rect 58268 60314 58296 60454
rect 58256 60308 58308 60314
rect 58256 60250 58308 60256
rect 58728 59702 58756 63294
rect 58990 63200 59046 63294
rect 58992 60036 59044 60042
rect 58992 59978 59044 59984
rect 58716 59696 58768 59702
rect 58716 59638 58768 59644
rect 58164 58676 58216 58682
rect 58164 58618 58216 58624
rect 58164 58540 58216 58546
rect 58164 58482 58216 58488
rect 58176 58313 58204 58482
rect 58162 58304 58218 58313
rect 58162 58239 58218 58248
rect 58164 57860 58216 57866
rect 58164 57802 58216 57808
rect 58176 57769 58204 57802
rect 58256 57792 58308 57798
rect 58162 57760 58218 57769
rect 58256 57734 58308 57740
rect 58162 57695 58218 57704
rect 58164 57452 58216 57458
rect 58164 57394 58216 57400
rect 58176 57225 58204 57394
rect 58162 57216 58218 57225
rect 58162 57151 58218 57160
rect 58268 57050 58296 57734
rect 58256 57044 58308 57050
rect 58256 56986 58308 56992
rect 58164 56772 58216 56778
rect 58164 56714 58216 56720
rect 58176 56681 58204 56714
rect 58162 56672 58218 56681
rect 58162 56607 58218 56616
rect 58348 56160 58400 56166
rect 58346 56128 58348 56137
rect 58400 56128 58402 56137
rect 58346 56063 58402 56072
rect 58348 54664 58400 54670
rect 58348 54606 58400 54612
rect 58360 54505 58388 54606
rect 58346 54496 58402 54505
rect 58346 54431 58402 54440
rect 58348 52896 58400 52902
rect 58346 52864 58348 52873
rect 58400 52864 58402 52873
rect 58346 52799 58402 52808
rect 58348 51400 58400 51406
rect 58348 51342 58400 51348
rect 58360 51241 58388 51342
rect 58346 51232 58402 51241
rect 58346 51167 58402 51176
rect 58900 49156 58952 49162
rect 58900 49098 58952 49104
rect 58348 48068 58400 48074
rect 58348 48010 58400 48016
rect 58164 43716 58216 43722
rect 58164 43658 58216 43664
rect 58176 43081 58204 43658
rect 58162 43072 58218 43081
rect 58162 43007 58218 43016
rect 58162 40352 58218 40361
rect 58162 40287 58218 40296
rect 58176 40118 58204 40287
rect 58164 40112 58216 40118
rect 58164 40054 58216 40060
rect 58256 38208 58308 38214
rect 58256 38150 58308 38156
rect 58164 37188 58216 37194
rect 58164 37130 58216 37136
rect 58176 36553 58204 37130
rect 58162 36544 58218 36553
rect 58162 36479 58218 36488
rect 58072 35080 58124 35086
rect 58072 35022 58124 35028
rect 58164 35012 58216 35018
rect 58164 34954 58216 34960
rect 58176 34921 58204 34954
rect 58162 34912 58218 34921
rect 58162 34847 58218 34856
rect 57978 34368 58034 34377
rect 57978 34303 58034 34312
rect 57992 33998 58020 34303
rect 57980 33992 58032 33998
rect 57980 33934 58032 33940
rect 58162 33280 58218 33289
rect 58162 33215 58218 33224
rect 58176 32978 58204 33215
rect 58164 32972 58216 32978
rect 58164 32914 58216 32920
rect 58164 31816 58216 31822
rect 58164 31758 58216 31764
rect 58176 31657 58204 31758
rect 58162 31648 58218 31657
rect 58162 31583 58218 31592
rect 57978 31104 58034 31113
rect 57978 31039 58034 31048
rect 57992 30734 58020 31039
rect 57980 30728 58032 30734
rect 57980 30670 58032 30676
rect 58072 30592 58124 30598
rect 58072 30534 58124 30540
rect 57978 27840 58034 27849
rect 57978 27775 58034 27784
rect 57992 27470 58020 27775
rect 57980 27464 58032 27470
rect 57980 27406 58032 27412
rect 58084 26330 58112 30534
rect 58162 30016 58218 30025
rect 58162 29951 58218 29960
rect 58176 29714 58204 29951
rect 58164 29708 58216 29714
rect 58164 29650 58216 29656
rect 58164 28484 58216 28490
rect 58164 28426 58216 28432
rect 58176 28393 58204 28426
rect 58162 28384 58218 28393
rect 58162 28319 58218 28328
rect 58162 26752 58218 26761
rect 58162 26687 58218 26696
rect 58176 26450 58204 26687
rect 58164 26444 58216 26450
rect 58164 26386 58216 26392
rect 57992 26302 58112 26330
rect 57888 24200 57940 24206
rect 57888 24142 57940 24148
rect 57796 23520 57848 23526
rect 57796 23462 57848 23468
rect 57900 21894 57928 24142
rect 57992 24070 58020 26302
rect 58070 26208 58126 26217
rect 58070 26143 58126 26152
rect 58084 25906 58112 26143
rect 58072 25900 58124 25906
rect 58072 25842 58124 25848
rect 58268 25786 58296 38150
rect 58360 26246 58388 48010
rect 58716 45892 58768 45898
rect 58716 45834 58768 45840
rect 58440 44804 58492 44810
rect 58440 44746 58492 44752
rect 58348 26240 58400 26246
rect 58348 26182 58400 26188
rect 58268 25758 58388 25786
rect 58452 25770 58480 44746
rect 58624 42628 58676 42634
rect 58624 42570 58676 42576
rect 58532 39364 58584 39370
rect 58532 39306 58584 39312
rect 58256 25696 58308 25702
rect 58256 25638 58308 25644
rect 58268 25430 58296 25638
rect 58256 25424 58308 25430
rect 58256 25366 58308 25372
rect 58164 25220 58216 25226
rect 58164 25162 58216 25168
rect 58176 25129 58204 25162
rect 58162 25120 58218 25129
rect 58162 25055 58218 25064
rect 58072 24812 58124 24818
rect 58072 24754 58124 24760
rect 58084 24585 58112 24754
rect 58360 24750 58388 25758
rect 58440 25764 58492 25770
rect 58440 25706 58492 25712
rect 58348 24744 58400 24750
rect 58348 24686 58400 24692
rect 58256 24608 58308 24614
rect 58070 24576 58126 24585
rect 58256 24550 58308 24556
rect 58070 24511 58126 24520
rect 58268 24410 58296 24550
rect 58256 24404 58308 24410
rect 58256 24346 58308 24352
rect 58164 24132 58216 24138
rect 58164 24074 58216 24080
rect 57980 24064 58032 24070
rect 57980 24006 58032 24012
rect 58176 23497 58204 24074
rect 58162 23488 58218 23497
rect 58162 23423 58218 23432
rect 58360 23322 58388 24686
rect 58348 23316 58400 23322
rect 58348 23258 58400 23264
rect 58070 22944 58126 22953
rect 58070 22879 58126 22888
rect 58084 22642 58112 22879
rect 58072 22636 58124 22642
rect 58072 22578 58124 22584
rect 58164 21956 58216 21962
rect 58164 21898 58216 21904
rect 57888 21888 57940 21894
rect 58176 21865 58204 21898
rect 57888 21830 57940 21836
rect 58162 21856 58218 21865
rect 58162 21791 58218 21800
rect 57716 21146 57836 21162
rect 57716 21140 57848 21146
rect 57716 21134 57796 21140
rect 57716 20806 57744 21134
rect 57796 21082 57848 21088
rect 57704 20800 57756 20806
rect 57704 20742 57756 20748
rect 57612 20596 57664 20602
rect 57612 20538 57664 20544
rect 58162 20224 58218 20233
rect 58162 20159 58218 20168
rect 58176 19922 58204 20159
rect 58164 19916 58216 19922
rect 58164 19858 58216 19864
rect 58072 19508 58124 19514
rect 58072 19450 58124 19456
rect 57888 18964 57940 18970
rect 57888 18906 57940 18912
rect 57242 18864 57298 18873
rect 57242 18799 57298 18808
rect 56876 18760 56928 18766
rect 56876 18702 56928 18708
rect 56968 18760 57020 18766
rect 56968 18702 57020 18708
rect 56784 18420 56836 18426
rect 56784 18362 56836 18368
rect 56508 18352 56560 18358
rect 56508 18294 56560 18300
rect 56692 18284 56744 18290
rect 56692 18226 56744 18232
rect 56600 16584 56652 16590
rect 56600 16526 56652 16532
rect 56612 16250 56640 16526
rect 56600 16244 56652 16250
rect 56600 16186 56652 16192
rect 56600 12844 56652 12850
rect 56600 12786 56652 12792
rect 56416 12776 56468 12782
rect 56416 12718 56468 12724
rect 56612 10742 56640 12786
rect 56600 10736 56652 10742
rect 56600 10678 56652 10684
rect 56600 10600 56652 10606
rect 56600 10542 56652 10548
rect 56324 9580 56376 9586
rect 56324 9522 56376 9528
rect 56336 8634 56364 9522
rect 56612 8838 56640 10542
rect 56600 8832 56652 8838
rect 56600 8774 56652 8780
rect 56704 8650 56732 18226
rect 56888 16658 56916 18702
rect 57900 18358 57928 18906
rect 58084 18426 58112 19450
rect 58162 18592 58218 18601
rect 58162 18527 58218 18536
rect 58072 18420 58124 18426
rect 58072 18362 58124 18368
rect 57888 18352 57940 18358
rect 57888 18294 57940 18300
rect 57980 18284 58032 18290
rect 57980 18226 58032 18232
rect 57058 18048 57114 18057
rect 57058 17983 57114 17992
rect 57072 17610 57100 17983
rect 57060 17604 57112 17610
rect 57060 17546 57112 17552
rect 57060 17196 57112 17202
rect 57060 17138 57112 17144
rect 56876 16652 56928 16658
rect 56876 16594 56928 16600
rect 56888 13394 56916 16594
rect 57072 16574 57100 17138
rect 57336 17128 57388 17134
rect 57336 17070 57388 17076
rect 57348 16969 57376 17070
rect 57334 16960 57390 16969
rect 57334 16895 57390 16904
rect 56980 16546 57100 16574
rect 57992 16574 58020 18226
rect 58176 17746 58204 18527
rect 58164 17740 58216 17746
rect 58164 17682 58216 17688
rect 57992 16546 58112 16574
rect 56980 16454 57008 16546
rect 56968 16448 57020 16454
rect 56968 16390 57020 16396
rect 57978 16416 58034 16425
rect 56980 16182 57008 16390
rect 57978 16351 58034 16360
rect 56968 16176 57020 16182
rect 56968 16118 57020 16124
rect 57992 15502 58020 16351
rect 58084 16114 58112 16546
rect 58072 16108 58124 16114
rect 58072 16050 58124 16056
rect 57980 15496 58032 15502
rect 57980 15438 58032 15444
rect 57244 15428 57296 15434
rect 57244 15370 57296 15376
rect 57256 15337 57284 15370
rect 57242 15328 57298 15337
rect 57242 15263 57298 15272
rect 57978 14784 58034 14793
rect 57978 14719 58034 14728
rect 57992 14414 58020 14719
rect 58072 14612 58124 14618
rect 58072 14554 58124 14560
rect 58084 14521 58112 14554
rect 58070 14512 58126 14521
rect 58070 14447 58126 14456
rect 57980 14408 58032 14414
rect 57980 14350 58032 14356
rect 58256 13932 58308 13938
rect 58256 13874 58308 13880
rect 57336 13864 57388 13870
rect 57336 13806 57388 13812
rect 57348 13705 57376 13806
rect 57334 13696 57390 13705
rect 57334 13631 57390 13640
rect 58268 13530 58296 13874
rect 58256 13524 58308 13530
rect 58256 13466 58308 13472
rect 56876 13388 56928 13394
rect 56876 13330 56928 13336
rect 56784 13252 56836 13258
rect 56784 13194 56836 13200
rect 56796 12714 56824 13194
rect 56784 12708 56836 12714
rect 56784 12650 56836 12656
rect 56888 12646 56916 13330
rect 57978 13152 58034 13161
rect 57978 13087 58034 13096
rect 57888 12776 57940 12782
rect 57888 12718 57940 12724
rect 56876 12640 56928 12646
rect 56876 12582 56928 12588
rect 56888 11218 56916 12582
rect 57244 12164 57296 12170
rect 57244 12106 57296 12112
rect 57256 12073 57284 12106
rect 57242 12064 57298 12073
rect 57242 11999 57298 12008
rect 57152 11756 57204 11762
rect 57152 11698 57204 11704
rect 57164 11529 57192 11698
rect 57244 11552 57296 11558
rect 57150 11520 57206 11529
rect 57244 11494 57296 11500
rect 57150 11455 57206 11464
rect 56876 11212 56928 11218
rect 56876 11154 56928 11160
rect 56784 11076 56836 11082
rect 56784 11018 56836 11024
rect 56796 10538 56824 11018
rect 56784 10532 56836 10538
rect 56784 10474 56836 10480
rect 56888 9042 56916 11154
rect 57152 10804 57204 10810
rect 57152 10746 57204 10752
rect 57060 9988 57112 9994
rect 57060 9930 57112 9936
rect 57072 9897 57100 9930
rect 57058 9888 57114 9897
rect 57058 9823 57114 9832
rect 56876 9036 56928 9042
rect 56876 8978 56928 8984
rect 56324 8628 56376 8634
rect 56324 8570 56376 8576
rect 56612 8622 56732 8650
rect 56232 8492 56284 8498
rect 56232 8434 56284 8440
rect 56140 8288 56192 8294
rect 56244 8265 56272 8434
rect 56140 8230 56192 8236
rect 56230 8256 56286 8265
rect 55312 7880 55364 7886
rect 55312 7822 55364 7828
rect 55324 2990 55352 7822
rect 56152 7818 56180 8230
rect 56230 8191 56286 8200
rect 56416 7880 56468 7886
rect 56416 7822 56468 7828
rect 56140 7812 56192 7818
rect 56140 7754 56192 7760
rect 55404 7268 55456 7274
rect 55404 7210 55456 7216
rect 55416 4826 55444 7210
rect 56152 5370 56180 7754
rect 56428 7698 56456 7822
rect 56244 7670 56456 7698
rect 56508 7744 56560 7750
rect 56508 7686 56560 7692
rect 56244 7342 56272 7670
rect 56520 7410 56548 7686
rect 56508 7404 56560 7410
rect 56508 7346 56560 7352
rect 56232 7336 56284 7342
rect 56232 7278 56284 7284
rect 56416 7336 56468 7342
rect 56416 7278 56468 7284
rect 56428 7177 56456 7278
rect 56612 7206 56640 8622
rect 56888 7954 56916 8978
rect 57164 8634 57192 10746
rect 57256 9654 57284 11494
rect 57900 10674 57928 12718
rect 57992 12238 58020 13087
rect 58268 12850 58296 13466
rect 58256 12844 58308 12850
rect 58256 12786 58308 12792
rect 57980 12232 58032 12238
rect 57980 12174 58032 12180
rect 58256 12164 58308 12170
rect 58256 12106 58308 12112
rect 58268 11354 58296 12106
rect 58256 11348 58308 11354
rect 58256 11290 58308 11296
rect 58268 10674 58296 11290
rect 57888 10668 57940 10674
rect 57888 10610 57940 10616
rect 58256 10668 58308 10674
rect 58256 10610 58308 10616
rect 57900 9654 57928 10610
rect 58162 10432 58218 10441
rect 58162 10367 58218 10376
rect 58176 10130 58204 10367
rect 58164 10124 58216 10130
rect 58164 10066 58216 10072
rect 57244 9648 57296 9654
rect 57244 9590 57296 9596
rect 57428 9648 57480 9654
rect 57428 9590 57480 9596
rect 57888 9648 57940 9654
rect 57888 9590 57940 9596
rect 57334 8800 57390 8809
rect 57334 8735 57390 8744
rect 57152 8628 57204 8634
rect 57152 8570 57204 8576
rect 57164 8294 57192 8570
rect 57348 8566 57376 8735
rect 57336 8560 57388 8566
rect 57336 8502 57388 8508
rect 57152 8288 57204 8294
rect 57152 8230 57204 8236
rect 56876 7948 56928 7954
rect 56876 7890 56928 7896
rect 56600 7200 56652 7206
rect 56414 7168 56470 7177
rect 56600 7142 56652 7148
rect 56414 7103 56470 7112
rect 55588 5364 55640 5370
rect 55588 5306 55640 5312
rect 56140 5364 56192 5370
rect 56140 5306 56192 5312
rect 55404 4820 55456 4826
rect 55404 4762 55456 4768
rect 55416 4146 55444 4762
rect 55600 4146 55628 5306
rect 56612 5234 56640 7142
rect 56888 6914 56916 7890
rect 57164 7410 57192 8230
rect 57440 8106 57468 9590
rect 57520 9580 57572 9586
rect 57520 9522 57572 9528
rect 57532 8838 57560 9522
rect 58256 9376 58308 9382
rect 58256 9318 58308 9324
rect 58072 8900 58124 8906
rect 58072 8842 58124 8848
rect 57520 8832 57572 8838
rect 57520 8774 57572 8780
rect 57532 8498 57560 8774
rect 57520 8492 57572 8498
rect 57520 8434 57572 8440
rect 58084 8362 58112 8842
rect 58268 8634 58296 9318
rect 58348 9172 58400 9178
rect 58348 9114 58400 9120
rect 58256 8628 58308 8634
rect 58256 8570 58308 8576
rect 58360 8498 58388 9114
rect 58348 8492 58400 8498
rect 58348 8434 58400 8440
rect 58544 8430 58572 39306
rect 58636 20058 58664 42570
rect 58728 26518 58756 45834
rect 58808 41540 58860 41546
rect 58808 41482 58860 41488
rect 58716 26512 58768 26518
rect 58716 26454 58768 26460
rect 58820 21622 58848 41482
rect 58912 25498 58940 49098
rect 59004 36650 59032 59978
rect 59176 59424 59228 59430
rect 59176 59366 59228 59372
rect 59084 38276 59136 38282
rect 59084 38218 59136 38224
rect 58992 36644 59044 36650
rect 58992 36586 59044 36592
rect 58992 33924 59044 33930
rect 58992 33866 59044 33872
rect 58900 25492 58952 25498
rect 58900 25434 58952 25440
rect 58808 21616 58860 21622
rect 58808 21558 58860 21564
rect 58624 20052 58676 20058
rect 58624 19994 58676 20000
rect 59004 19242 59032 33866
rect 59096 24206 59124 38218
rect 59188 37126 59216 59366
rect 59176 37120 59228 37126
rect 59176 37062 59228 37068
rect 59176 36100 59228 36106
rect 59176 36042 59228 36048
rect 59084 24200 59136 24206
rect 59084 24142 59136 24148
rect 58992 19236 59044 19242
rect 58992 19178 59044 19184
rect 59188 18630 59216 36042
rect 59176 18624 59228 18630
rect 59176 18566 59228 18572
rect 58532 8424 58584 8430
rect 58532 8366 58584 8372
rect 58072 8356 58124 8362
rect 58072 8298 58124 8304
rect 57256 8090 57468 8106
rect 57244 8084 57468 8090
rect 57296 8078 57468 8084
rect 57244 8026 57296 8032
rect 57440 7478 57468 8078
rect 57244 7472 57296 7478
rect 57244 7414 57296 7420
rect 57428 7472 57480 7478
rect 57428 7414 57480 7420
rect 57612 7472 57664 7478
rect 57612 7414 57664 7420
rect 57152 7404 57204 7410
rect 57152 7346 57204 7352
rect 56704 6886 56916 6914
rect 56704 6798 56732 6886
rect 56692 6792 56744 6798
rect 56692 6734 56744 6740
rect 56600 5228 56652 5234
rect 56600 5170 56652 5176
rect 56612 4690 56640 5170
rect 56600 4684 56652 4690
rect 56600 4626 56652 4632
rect 56600 4548 56652 4554
rect 56600 4490 56652 4496
rect 55404 4140 55456 4146
rect 55404 4082 55456 4088
rect 55588 4140 55640 4146
rect 55588 4082 55640 4088
rect 56612 3126 56640 4490
rect 56704 3942 56732 6734
rect 57256 6322 57284 7414
rect 57520 7200 57572 7206
rect 57520 7142 57572 7148
rect 57532 6798 57560 7142
rect 57520 6792 57572 6798
rect 57520 6734 57572 6740
rect 57520 6656 57572 6662
rect 57520 6598 57572 6604
rect 57532 6322 57560 6598
rect 57624 6458 57652 7414
rect 57978 6624 58034 6633
rect 57978 6559 58034 6568
rect 57612 6452 57664 6458
rect 57612 6394 57664 6400
rect 57244 6316 57296 6322
rect 57244 6258 57296 6264
rect 57520 6316 57572 6322
rect 57520 6258 57572 6264
rect 57532 5710 57560 6258
rect 57992 5710 58020 6559
rect 57520 5704 57572 5710
rect 57520 5646 57572 5652
rect 57980 5704 58032 5710
rect 57980 5646 58032 5652
rect 57244 5636 57296 5642
rect 57244 5578 57296 5584
rect 57256 5545 57284 5578
rect 57242 5536 57298 5545
rect 57242 5471 57298 5480
rect 58072 5228 58124 5234
rect 58072 5170 58124 5176
rect 58084 5001 58112 5170
rect 58256 5024 58308 5030
rect 58070 4992 58126 5001
rect 58256 4966 58308 4972
rect 58070 4927 58126 4936
rect 57980 4616 58032 4622
rect 57980 4558 58032 4564
rect 58164 4616 58216 4622
rect 58164 4558 58216 4564
rect 56692 3936 56744 3942
rect 56692 3878 56744 3884
rect 57428 3936 57480 3942
rect 57428 3878 57480 3884
rect 56704 3602 56732 3878
rect 56692 3596 56744 3602
rect 56692 3538 56744 3544
rect 57440 3534 57468 3878
rect 57428 3528 57480 3534
rect 57428 3470 57480 3476
rect 57244 3392 57296 3398
rect 57244 3334 57296 3340
rect 56600 3120 56652 3126
rect 56600 3062 56652 3068
rect 56508 3052 56560 3058
rect 56508 2994 56560 3000
rect 55312 2984 55364 2990
rect 55312 2926 55364 2932
rect 54760 2508 54812 2514
rect 54760 2450 54812 2456
rect 53656 2440 53708 2446
rect 53656 2382 53708 2388
rect 53668 800 53696 2382
rect 53932 2372 53984 2378
rect 53932 2314 53984 2320
rect 53944 800 53972 2314
rect 55680 2304 55732 2310
rect 55680 2246 55732 2252
rect 56416 2304 56468 2310
rect 56416 2246 56468 2252
rect 55692 2106 55720 2246
rect 55680 2100 55732 2106
rect 55680 2042 55732 2048
rect 56428 2038 56456 2246
rect 56416 2032 56468 2038
rect 56416 1974 56468 1980
rect 56520 1737 56548 2994
rect 57256 2446 57284 3334
rect 57992 3058 58020 4558
rect 58072 4140 58124 4146
rect 58072 4082 58124 4088
rect 58084 3913 58112 4082
rect 58070 3904 58126 3913
rect 58070 3839 58126 3848
rect 58176 3482 58204 4558
rect 58268 4282 58296 4966
rect 58256 4276 58308 4282
rect 58256 4218 58308 4224
rect 58256 3936 58308 3942
rect 58256 3878 58308 3884
rect 58268 3738 58296 3878
rect 58256 3732 58308 3738
rect 58256 3674 58308 3680
rect 58176 3454 58296 3482
rect 58162 3360 58218 3369
rect 58162 3295 58218 3304
rect 58176 3126 58204 3295
rect 58268 3194 58296 3454
rect 58256 3188 58308 3194
rect 58256 3130 58308 3136
rect 58164 3120 58216 3126
rect 58164 3062 58216 3068
rect 57980 3052 58032 3058
rect 57980 2994 58032 3000
rect 57992 2650 58020 2994
rect 58162 2816 58218 2825
rect 58162 2751 58218 2760
rect 57980 2644 58032 2650
rect 57980 2586 58032 2592
rect 58176 2446 58204 2751
rect 57244 2440 57296 2446
rect 57244 2382 57296 2388
rect 58164 2440 58216 2446
rect 58164 2382 58216 2388
rect 57336 2372 57388 2378
rect 57336 2314 57388 2320
rect 57348 2281 57376 2314
rect 57334 2272 57390 2281
rect 57334 2207 57390 2216
rect 56506 1728 56562 1737
rect 56506 1663 56562 1672
rect 56508 1352 56560 1358
rect 56508 1294 56560 1300
rect 56520 1193 56548 1294
rect 56506 1184 56562 1193
rect 56506 1119 56562 1128
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12806 0 12862 800
rect 13082 0 13138 800
rect 13358 0 13414 800
rect 13634 0 13690 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17222 0 17278 800
rect 17498 0 17554 800
rect 17774 0 17830 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 19982 0 20038 800
rect 20258 0 20314 800
rect 20534 0 20590 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25778 0 25834 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27710 0 27766 800
rect 27986 0 28042 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29366 0 29422 800
rect 29642 0 29698 800
rect 29918 0 29974 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32954 0 33010 800
rect 33230 0 33286 800
rect 33506 0 33562 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35162 0 35218 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43442 0 43498 800
rect 43718 0 43774 800
rect 43994 0 44050 800
rect 44270 0 44326 800
rect 44546 0 44602 800
rect 44822 0 44878 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50342 0 50398 800
rect 50618 0 50674 800
rect 50894 0 50950 800
rect 51170 0 51226 800
rect 51446 0 51502 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 53930 0 53986 800
<< via2 >>
rect 1674 60832 1730 60888
rect 1674 60152 1730 60208
rect 1582 59472 1638 59528
rect 2778 61512 2834 61568
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 1582 58792 1638 58848
rect 1674 58112 1730 58168
rect 1582 57432 1638 57488
rect 1674 56788 1676 56808
rect 1676 56788 1728 56808
rect 1728 56788 1730 56808
rect 1674 56752 1730 56788
rect 1674 56072 1730 56128
rect 1674 55392 1730 55448
rect 1582 54712 1638 54768
rect 1674 54032 1730 54088
rect 1582 53352 1638 53408
rect 1582 52672 1638 52728
rect 1674 51992 1730 52048
rect 1674 51332 1730 51368
rect 1674 51312 1676 51332
rect 1676 51312 1728 51332
rect 1728 51312 1730 51332
rect 1674 50632 1730 50688
rect 1674 49952 1730 50008
rect 1674 49272 1730 49328
rect 1674 48592 1730 48648
rect 1674 47912 1730 47968
rect 1398 40432 1454 40488
rect 1398 38392 1454 38448
rect 1398 35672 1454 35728
rect 1674 47232 1730 47288
rect 1674 46552 1730 46608
rect 1674 45892 1730 45928
rect 1674 45872 1676 45892
rect 1676 45872 1728 45892
rect 1728 45872 1730 45892
rect 1582 45192 1638 45248
rect 1674 44512 1730 44568
rect 1674 43832 1730 43888
rect 1582 43152 1638 43208
rect 1674 42472 1730 42528
rect 1674 41792 1730 41848
rect 1674 41112 1730 41168
rect 1674 39752 1730 39808
rect 1582 39072 1638 39128
rect 1674 37712 1730 37768
rect 1582 36352 1638 36408
rect 1674 34992 1730 35048
rect 1674 34312 1730 34368
rect 1674 33632 1730 33688
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 1674 32952 1730 33008
rect 1674 32272 1730 32328
rect 1674 31592 1730 31648
rect 1674 30912 1730 30968
rect 1674 30232 1730 30288
rect 1858 29572 1914 29608
rect 1858 29552 1860 29572
rect 1860 29552 1912 29572
rect 1912 29552 1914 29572
rect 1766 28872 1822 28928
rect 1858 28192 1914 28248
rect 1582 27512 1638 27568
rect 1766 26868 1768 26888
rect 1768 26868 1820 26888
rect 1820 26868 1822 26888
rect 1766 26832 1822 26868
rect 1858 26152 1914 26208
rect 1766 25472 1822 25528
rect 1858 24792 1914 24848
rect 1858 24132 1914 24168
rect 1858 24112 1860 24132
rect 1860 24112 1912 24132
rect 1912 24112 1914 24132
rect 1766 23432 1822 23488
rect 1858 22752 1914 22808
rect 1766 22072 1822 22128
rect 1858 21428 1860 21448
rect 1860 21428 1912 21448
rect 1912 21428 1914 21448
rect 1858 21392 1914 21428
rect 1858 20712 1914 20768
rect 1766 20032 1822 20088
rect 1858 19352 1914 19408
rect 1858 18692 1914 18728
rect 1858 18672 1860 18692
rect 1860 18672 1912 18692
rect 1912 18672 1914 18692
rect 1766 17992 1822 18048
rect 1858 17312 1914 17368
rect 1766 16632 1822 16688
rect 1766 15988 1768 16008
rect 1768 15988 1820 16008
rect 1820 15988 1822 16008
rect 1766 15952 1822 15988
rect 1858 15272 1914 15328
rect 1766 14592 1822 14648
rect 1858 13912 1914 13968
rect 1858 13268 1860 13288
rect 1860 13268 1912 13288
rect 1912 13268 1914 13288
rect 1858 13232 1914 13268
rect 1766 12552 1822 12608
rect 1858 11872 1914 11928
rect 1766 11192 1822 11248
rect 1766 10548 1768 10568
rect 1768 10548 1820 10568
rect 1820 10548 1822 10568
rect 1766 10512 1822 10548
rect 1858 9832 1914 9888
rect 1766 9152 1822 9208
rect 1858 8472 1914 8528
rect 1858 7812 1914 7848
rect 1858 7792 1860 7812
rect 1860 7792 1912 7812
rect 1912 7792 1914 7812
rect 1766 7112 1822 7168
rect 1858 6432 1914 6488
rect 1582 5888 1638 5944
rect 1766 5752 1822 5808
rect 2410 37032 2466 37088
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 7838 61140 7840 61160
rect 7840 61140 7892 61160
rect 7892 61140 7894 61160
rect 7838 61104 7894 61140
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 2042 6704 2098 6760
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 1950 5616 2006 5672
rect 1766 5108 1768 5128
rect 1768 5108 1820 5128
rect 1820 5108 1822 5128
rect 1766 5072 1822 5108
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 1858 4392 1914 4448
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 1766 3712 1822 3768
rect 1858 3032 1914 3088
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 1858 2388 1860 2408
rect 1860 2388 1912 2408
rect 1912 2388 1914 2408
rect 1858 2352 1914 2388
rect 8298 3848 8354 3904
rect 9954 3712 10010 3768
rect 9678 3188 9734 3224
rect 9678 3168 9680 3188
rect 9680 3168 9732 3188
rect 9732 3168 9734 3188
rect 9678 3052 9734 3088
rect 9678 3032 9680 3052
rect 9680 3032 9732 3052
rect 9732 3032 9734 3052
rect 9586 2760 9642 2816
rect 10598 3168 10654 3224
rect 11610 3440 11666 3496
rect 12346 3032 12402 3088
rect 11978 2760 12034 2816
rect 13542 17176 13598 17232
rect 13910 9016 13966 9072
rect 14094 8880 14150 8936
rect 13542 2916 13598 2952
rect 13542 2896 13544 2916
rect 13544 2896 13596 2916
rect 13596 2896 13598 2916
rect 13726 4004 13782 4040
rect 13726 3984 13728 4004
rect 13728 3984 13780 4004
rect 13780 3984 13782 4004
rect 13726 3596 13782 3632
rect 13726 3576 13728 3596
rect 13728 3576 13780 3596
rect 13780 3576 13782 3596
rect 16762 58540 16818 58576
rect 16762 58520 16764 58540
rect 16764 58520 16816 58540
rect 16816 58520 16818 58540
rect 17406 58540 17462 58576
rect 17406 58520 17408 58540
rect 17408 58520 17460 58540
rect 17460 58520 17462 58540
rect 15014 11736 15070 11792
rect 14738 4528 14794 4584
rect 16762 13368 16818 13424
rect 19580 60954 19636 60956
rect 19660 60954 19716 60956
rect 19740 60954 19796 60956
rect 19820 60954 19876 60956
rect 19580 60902 19626 60954
rect 19626 60902 19636 60954
rect 19660 60902 19690 60954
rect 19690 60902 19702 60954
rect 19702 60902 19716 60954
rect 19740 60902 19754 60954
rect 19754 60902 19766 60954
rect 19766 60902 19796 60954
rect 19820 60902 19830 60954
rect 19830 60902 19876 60954
rect 19580 60900 19636 60902
rect 19660 60900 19716 60902
rect 19740 60900 19796 60902
rect 19820 60900 19876 60902
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19706 37712 19762 37768
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19522 33088 19578 33144
rect 19614 32988 19616 33008
rect 19616 32988 19668 33008
rect 19668 32988 19670 33008
rect 19614 32952 19670 32988
rect 19890 32952 19946 33008
rect 19338 32716 19340 32736
rect 19340 32716 19392 32736
rect 19392 32716 19394 32736
rect 19338 32680 19394 32716
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 20074 33088 20130 33144
rect 19798 32020 19854 32056
rect 19798 32000 19800 32020
rect 19800 32000 19852 32020
rect 19852 32000 19854 32020
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 20350 32952 20406 33008
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19982 29960 20038 30016
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 17314 16496 17370 16552
rect 17130 14728 17186 14784
rect 17406 14728 17462 14784
rect 16946 6316 17002 6352
rect 16946 6296 16948 6316
rect 16948 6296 17000 6316
rect 17000 6296 17002 6316
rect 18142 16496 18198 16552
rect 18234 16108 18290 16144
rect 18234 16088 18236 16108
rect 18236 16088 18288 16108
rect 18288 16088 18290 16108
rect 17866 6452 17922 6488
rect 17866 6432 17868 6452
rect 17868 6432 17920 6452
rect 17920 6432 17922 6452
rect 17314 3168 17370 3224
rect 17866 3032 17922 3088
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 20902 32020 20958 32056
rect 20902 32000 20904 32020
rect 20904 32000 20956 32020
rect 20956 32000 20958 32020
rect 21178 32852 21180 32872
rect 21180 32852 21232 32872
rect 21232 32852 21234 32872
rect 21178 32816 21234 32852
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 18694 3884 18696 3904
rect 18696 3884 18748 3904
rect 18748 3884 18750 3904
rect 18694 3848 18750 3884
rect 19154 10104 19210 10160
rect 19062 8236 19064 8256
rect 19064 8236 19116 8256
rect 19116 8236 19118 8256
rect 19062 8200 19118 8236
rect 19982 16768 20038 16824
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19522 15444 19524 15464
rect 19524 15444 19576 15464
rect 19576 15444 19578 15464
rect 19522 15408 19578 15444
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19430 15000 19486 15056
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19890 12316 19892 12336
rect 19892 12316 19944 12336
rect 19944 12316 19946 12336
rect 19890 12280 19946 12316
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19798 11636 19800 11656
rect 19800 11636 19852 11656
rect 19852 11636 19854 11656
rect 19798 11600 19854 11636
rect 19338 11192 19394 11248
rect 19246 6432 19302 6488
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 20074 10240 20130 10296
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19798 7268 19854 7304
rect 19798 7248 19800 7268
rect 19800 7248 19852 7268
rect 19852 7248 19854 7268
rect 20534 16360 20590 16416
rect 20350 11192 20406 11248
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 20258 6568 20314 6624
rect 19154 4528 19210 4584
rect 18970 3884 18972 3904
rect 18972 3884 19024 3904
rect 19024 3884 19026 3904
rect 18970 3848 19026 3884
rect 19246 3848 19302 3904
rect 19246 3712 19302 3768
rect 18970 3304 19026 3360
rect 19154 3340 19156 3360
rect 19156 3340 19208 3360
rect 19208 3340 19210 3360
rect 19154 3304 19210 3340
rect 19246 3168 19302 3224
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19798 5208 19854 5264
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19430 3712 19486 3768
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20074 2624 20130 2680
rect 21086 17312 21142 17368
rect 21454 15952 21510 16008
rect 21362 14456 21418 14512
rect 22926 35264 22982 35320
rect 22742 29144 22798 29200
rect 21822 15408 21878 15464
rect 21362 12960 21418 13016
rect 20994 12316 20996 12336
rect 20996 12316 21048 12336
rect 21048 12316 21050 12336
rect 20994 12280 21050 12316
rect 20718 8200 20774 8256
rect 20442 2896 20498 2952
rect 21546 10376 21602 10432
rect 22650 17312 22706 17368
rect 22650 17040 22706 17096
rect 24766 36100 24822 36136
rect 24766 36080 24768 36100
rect 24768 36080 24820 36100
rect 24820 36080 24822 36100
rect 24122 35012 24178 35048
rect 24122 34992 24124 35012
rect 24124 34992 24176 35012
rect 24176 34992 24178 35012
rect 24122 29008 24178 29064
rect 22834 17584 22890 17640
rect 22006 10260 22062 10296
rect 22006 10240 22008 10260
rect 22008 10240 22060 10260
rect 22060 10240 22062 10260
rect 22098 10104 22154 10160
rect 22190 6976 22246 7032
rect 22098 6840 22154 6896
rect 21638 6432 21694 6488
rect 22006 6024 22062 6080
rect 22374 6704 22430 6760
rect 22466 5772 22522 5808
rect 22466 5752 22468 5772
rect 22468 5752 22520 5772
rect 22520 5752 22522 5772
rect 22466 4800 22522 4856
rect 22006 3712 22062 3768
rect 22282 3032 22338 3088
rect 23202 15952 23258 16008
rect 22834 6568 22890 6624
rect 22834 4664 22890 4720
rect 23570 15444 23572 15464
rect 23572 15444 23624 15464
rect 23624 15444 23626 15464
rect 23570 15408 23626 15444
rect 23754 10004 23756 10024
rect 23756 10004 23808 10024
rect 23808 10004 23810 10024
rect 23570 9716 23626 9752
rect 23754 9968 23810 10004
rect 23570 9696 23572 9716
rect 23572 9696 23624 9716
rect 23624 9696 23626 9716
rect 23570 6840 23626 6896
rect 24030 6432 24086 6488
rect 25226 35284 25282 35320
rect 25226 35264 25228 35284
rect 25228 35264 25280 35284
rect 25280 35264 25282 35284
rect 25502 35012 25558 35048
rect 25502 34992 25504 35012
rect 25504 34992 25556 35012
rect 25556 34992 25558 35012
rect 24582 18400 24638 18456
rect 24214 5208 24270 5264
rect 24490 11464 24546 11520
rect 24582 6860 24638 6896
rect 24582 6840 24584 6860
rect 24584 6840 24636 6860
rect 24636 6840 24638 6860
rect 24582 5636 24638 5672
rect 24582 5616 24584 5636
rect 24584 5616 24636 5636
rect 24636 5616 24638 5636
rect 24766 4700 24768 4720
rect 24768 4700 24820 4720
rect 24820 4700 24822 4720
rect 24766 4664 24822 4700
rect 25134 6740 25136 6760
rect 25136 6740 25188 6760
rect 25188 6740 25190 6760
rect 25134 6704 25190 6740
rect 25134 6024 25190 6080
rect 25502 17060 25558 17096
rect 25502 17040 25504 17060
rect 25504 17040 25556 17060
rect 25556 17040 25558 17060
rect 25410 16396 25412 16416
rect 25412 16396 25464 16416
rect 25464 16396 25466 16416
rect 25410 16360 25466 16396
rect 25410 14456 25466 14512
rect 25318 14320 25374 14376
rect 25870 18808 25926 18864
rect 26238 18264 26294 18320
rect 26514 30096 26570 30152
rect 26698 22888 26754 22944
rect 26606 18264 26662 18320
rect 26330 18128 26386 18184
rect 25134 4800 25190 4856
rect 24950 3848 25006 3904
rect 25502 9968 25558 10024
rect 27158 23160 27214 23216
rect 27526 38664 27582 38720
rect 27526 22072 27582 22128
rect 27802 22072 27858 22128
rect 27526 21936 27582 21992
rect 27802 20848 27858 20904
rect 27618 19252 27620 19272
rect 27620 19252 27672 19272
rect 27672 19252 27674 19272
rect 27618 19216 27674 19252
rect 26790 14728 26846 14784
rect 27158 17992 27214 18048
rect 27802 19352 27858 19408
rect 26790 10412 26792 10432
rect 26792 10412 26844 10432
rect 26844 10412 26846 10432
rect 26790 10376 26846 10412
rect 26054 8336 26110 8392
rect 25594 5772 25650 5808
rect 25594 5752 25596 5772
rect 25596 5752 25648 5772
rect 25648 5752 25650 5772
rect 25778 5652 25780 5672
rect 25780 5652 25832 5672
rect 25832 5652 25834 5672
rect 25778 5616 25834 5652
rect 26514 6432 26570 6488
rect 27066 10648 27122 10704
rect 26974 10376 27030 10432
rect 27434 9424 27490 9480
rect 26974 4020 26976 4040
rect 26976 4020 27028 4040
rect 27028 4020 27030 4040
rect 25962 3576 26018 3632
rect 26974 3984 27030 4020
rect 27158 7248 27214 7304
rect 28078 18828 28134 18864
rect 28078 18808 28080 18828
rect 28080 18808 28132 18828
rect 28132 18808 28134 18828
rect 27710 6432 27766 6488
rect 28262 19080 28318 19136
rect 28814 20884 28816 20904
rect 28816 20884 28868 20904
rect 28868 20884 28870 20904
rect 28814 20848 28870 20884
rect 28538 19508 28594 19544
rect 28538 19488 28540 19508
rect 28540 19488 28592 19508
rect 28592 19488 28594 19508
rect 28538 19372 28594 19408
rect 28538 19352 28540 19372
rect 28540 19352 28592 19372
rect 28592 19352 28594 19372
rect 28446 18536 28502 18592
rect 28354 17448 28410 17504
rect 28262 16360 28318 16416
rect 28538 17992 28594 18048
rect 28814 18400 28870 18456
rect 29182 19488 29238 19544
rect 29090 19352 29146 19408
rect 28998 18164 29000 18184
rect 29000 18164 29052 18184
rect 29052 18164 29054 18184
rect 28998 18128 29054 18164
rect 29182 17040 29238 17096
rect 29642 22888 29698 22944
rect 33322 60832 33378 60888
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 33230 60696 33286 60752
rect 35070 60696 35126 60752
rect 29918 23024 29974 23080
rect 30378 23060 30380 23080
rect 30380 23060 30432 23080
rect 30432 23060 30434 23080
rect 30378 23024 30434 23060
rect 29458 19488 29514 19544
rect 29458 17604 29514 17640
rect 29458 17584 29460 17604
rect 29460 17584 29512 17604
rect 29512 17584 29514 17604
rect 29366 16668 29368 16688
rect 29368 16668 29420 16688
rect 29420 16668 29422 16688
rect 29366 16632 29422 16668
rect 28170 9424 28226 9480
rect 28630 6976 28686 7032
rect 28630 5616 28686 5672
rect 29274 10668 29330 10704
rect 29274 10648 29276 10668
rect 29276 10648 29328 10668
rect 29328 10648 29330 10668
rect 29182 9696 29238 9752
rect 30010 21972 30012 21992
rect 30012 21972 30064 21992
rect 30064 21972 30066 21992
rect 30010 21936 30066 21972
rect 30562 19080 30618 19136
rect 29734 17720 29790 17776
rect 30746 18944 30802 19000
rect 30010 17584 30066 17640
rect 30102 17312 30158 17368
rect 30746 18400 30802 18456
rect 30838 18128 30894 18184
rect 30470 17992 30526 18048
rect 30286 16904 30342 16960
rect 30562 17856 30618 17912
rect 28906 3460 28962 3496
rect 28906 3440 28908 3460
rect 28908 3440 28960 3460
rect 28960 3440 28962 3460
rect 31022 17856 31078 17912
rect 30746 17312 30802 17368
rect 30930 16632 30986 16688
rect 31114 16496 31170 16552
rect 30746 13912 30802 13968
rect 31298 19252 31300 19272
rect 31300 19252 31352 19272
rect 31352 19252 31354 19272
rect 31298 19216 31354 19252
rect 31298 18672 31354 18728
rect 30010 9696 30066 9752
rect 30562 10376 30618 10432
rect 30378 9560 30434 9616
rect 30286 9460 30288 9480
rect 30288 9460 30340 9480
rect 30340 9460 30342 9480
rect 30286 9424 30342 9460
rect 31114 10648 31170 10704
rect 31206 9424 31262 9480
rect 31574 18572 31576 18592
rect 31576 18572 31628 18592
rect 31628 18572 31630 18592
rect 31574 18536 31630 18572
rect 31574 16632 31630 16688
rect 31482 14356 31484 14376
rect 31484 14356 31536 14376
rect 31536 14356 31538 14376
rect 31482 14320 31538 14356
rect 32034 20576 32090 20632
rect 32034 18944 32090 19000
rect 33138 29008 33194 29064
rect 32586 24676 32642 24712
rect 32586 24656 32588 24676
rect 32588 24656 32640 24676
rect 32640 24656 32642 24676
rect 33598 22752 33654 22808
rect 32034 17856 32090 17912
rect 32126 17584 32182 17640
rect 31942 17040 31998 17096
rect 32586 19488 32642 19544
rect 32678 17992 32734 18048
rect 33138 18400 33194 18456
rect 32862 17992 32918 18048
rect 33138 17856 33194 17912
rect 32494 16768 32550 16824
rect 32310 13912 32366 13968
rect 31574 12960 31630 13016
rect 31482 10376 31538 10432
rect 32126 8916 32128 8936
rect 32128 8916 32180 8936
rect 32180 8916 32182 8936
rect 32126 8880 32182 8916
rect 31574 8336 31630 8392
rect 31850 6452 31906 6488
rect 31850 6432 31852 6452
rect 31852 6432 31904 6452
rect 31904 6432 31906 6452
rect 33230 17448 33286 17504
rect 32862 8900 32918 8936
rect 32862 8880 32864 8900
rect 32864 8880 32916 8900
rect 32916 8880 32918 8900
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 35346 56616 35402 56672
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 33966 23568 34022 23624
rect 33874 23044 33930 23080
rect 33874 23024 33876 23044
rect 33876 23024 33928 23044
rect 33928 23024 33930 23044
rect 34150 22616 34206 22672
rect 33598 17176 33654 17232
rect 34150 22480 34206 22536
rect 33874 14864 33930 14920
rect 33414 11600 33470 11656
rect 33230 6296 33286 6352
rect 33690 11756 33746 11792
rect 33690 11736 33692 11756
rect 33692 11736 33744 11756
rect 33744 11736 33746 11756
rect 34334 18264 34390 18320
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35162 31184 35218 31240
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35070 23588 35126 23624
rect 35070 23568 35072 23588
rect 35072 23568 35124 23588
rect 35124 23568 35126 23588
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34702 19216 34758 19272
rect 34518 16904 34574 16960
rect 34334 15544 34390 15600
rect 33966 11756 34022 11792
rect 33966 11736 33968 11756
rect 33968 11736 34020 11756
rect 34020 11736 34022 11756
rect 33690 9696 33746 9752
rect 33782 7384 33838 7440
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34886 18400 34942 18456
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34702 11736 34758 11792
rect 34150 7948 34206 7984
rect 34150 7928 34152 7948
rect 34152 7928 34204 7948
rect 34204 7928 34206 7948
rect 35346 11600 35402 11656
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35070 9580 35126 9616
rect 35070 9560 35072 9580
rect 35072 9560 35124 9580
rect 35124 9560 35126 9580
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34886 8492 34942 8528
rect 34886 8472 34888 8492
rect 34888 8472 34940 8492
rect 34940 8472 34942 8492
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35714 31184 35770 31240
rect 35714 22888 35770 22944
rect 35714 22616 35770 22672
rect 35622 22480 35678 22536
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 38106 57296 38162 57352
rect 36450 23024 36506 23080
rect 36450 22752 36506 22808
rect 36358 18536 36414 18592
rect 36358 16496 36414 16552
rect 36542 19216 36598 19272
rect 37554 23568 37610 23624
rect 37002 18672 37058 18728
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36450 7384 36506 7440
rect 37278 8336 37334 8392
rect 38842 23044 38898 23080
rect 38842 23024 38844 23044
rect 38844 23024 38896 23044
rect 38896 23024 38898 23044
rect 38106 18128 38162 18184
rect 38198 17720 38254 17776
rect 38106 7928 38162 7984
rect 38658 16632 38714 16688
rect 38658 8492 38714 8528
rect 38658 8472 38660 8492
rect 38660 8472 38712 8492
rect 38712 8472 38714 8492
rect 42062 53080 42118 53136
rect 38658 7420 38660 7440
rect 38660 7420 38712 7440
rect 38712 7420 38714 7440
rect 38658 7384 38714 7420
rect 39118 3340 39120 3360
rect 39120 3340 39172 3360
rect 39172 3340 39174 3360
rect 39118 3304 39174 3340
rect 39486 5616 39542 5672
rect 39670 22924 39672 22944
rect 39672 22924 39724 22944
rect 39724 22924 39726 22944
rect 39670 22888 39726 22924
rect 39946 20576 40002 20632
rect 40222 22924 40224 22944
rect 40224 22924 40276 22944
rect 40276 22924 40278 22944
rect 40222 22888 40278 22924
rect 40314 21664 40370 21720
rect 40682 23024 40738 23080
rect 40682 22072 40738 22128
rect 40590 21528 40646 21584
rect 39946 7384 40002 7440
rect 41142 13640 41198 13696
rect 41050 3596 41106 3632
rect 41050 3576 41052 3596
rect 41052 3576 41104 3596
rect 41104 3576 41106 3596
rect 42522 23160 42578 23216
rect 42798 23060 42800 23080
rect 42800 23060 42852 23080
rect 42852 23060 42854 23080
rect 42798 23024 42854 23060
rect 42614 3712 42670 3768
rect 43074 3168 43130 3224
rect 43350 3304 43406 3360
rect 43350 3032 43406 3088
rect 43902 23060 43904 23080
rect 43904 23060 43956 23080
rect 43956 23060 43958 23080
rect 43902 23024 43958 23060
rect 43994 21800 44050 21856
rect 43902 21528 43958 21584
rect 43902 16632 43958 16688
rect 43718 3576 43774 3632
rect 45006 14864 45062 14920
rect 45374 22108 45376 22128
rect 45376 22108 45428 22128
rect 45428 22108 45430 22128
rect 45374 22072 45430 22108
rect 45374 21800 45430 21856
rect 45190 3476 45192 3496
rect 45192 3476 45244 3496
rect 45244 3476 45246 3496
rect 45190 3440 45246 3476
rect 44914 2896 44970 2952
rect 45098 3052 45154 3088
rect 45098 3032 45100 3052
rect 45100 3032 45152 3052
rect 45152 3032 45154 3052
rect 45742 3052 45798 3088
rect 45742 3032 45744 3052
rect 45744 3032 45796 3052
rect 45796 3032 45798 3052
rect 45650 2932 45652 2952
rect 45652 2932 45704 2952
rect 45704 2932 45706 2952
rect 45650 2896 45706 2932
rect 50300 60954 50356 60956
rect 50380 60954 50436 60956
rect 50460 60954 50516 60956
rect 50540 60954 50596 60956
rect 50300 60902 50346 60954
rect 50346 60902 50356 60954
rect 50380 60902 50410 60954
rect 50410 60902 50422 60954
rect 50422 60902 50436 60954
rect 50460 60902 50474 60954
rect 50474 60902 50486 60954
rect 50486 60902 50516 60954
rect 50540 60902 50550 60954
rect 50550 60902 50596 60954
rect 50300 60900 50356 60902
rect 50380 60900 50436 60902
rect 50460 60900 50516 60902
rect 50540 60900 50596 60902
rect 47858 21684 47914 21720
rect 47858 21664 47860 21684
rect 47860 21664 47912 21684
rect 47912 21664 47914 21684
rect 46846 3168 46902 3224
rect 47122 3712 47178 3768
rect 47950 2352 48006 2408
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 49698 19352 49754 19408
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 50894 3612 50896 3632
rect 50896 3612 50948 3632
rect 50948 3612 50950 3632
rect 50894 3576 50950 3612
rect 56046 62600 56102 62656
rect 56138 62056 56194 62112
rect 56138 60968 56194 61024
rect 56506 61512 56562 61568
rect 52458 3032 52514 3088
rect 57334 60424 57390 60480
rect 57978 59880 58034 59936
rect 57794 59336 57850 59392
rect 57886 58792 57942 58848
rect 57334 47912 57390 47968
rect 56966 42472 57022 42528
rect 57058 39208 57114 39264
rect 57242 44648 57298 44704
rect 57242 41384 57298 41440
rect 57242 38120 57298 38176
rect 57058 32680 57114 32736
rect 56322 21936 56378 21992
rect 57058 29416 57114 29472
rect 57150 21256 57206 21312
rect 57058 19624 57114 19680
rect 57886 49544 57942 49600
rect 57978 49000 58034 49056
rect 57978 47368 58034 47424
rect 57886 46280 57942 46336
rect 57978 45736 58034 45792
rect 57886 44104 57942 44160
rect 57886 41928 57942 41984
rect 57886 40840 57942 40896
rect 57886 39752 57942 39808
rect 57978 38664 58034 38720
rect 57886 37576 57942 37632
rect 57978 35944 58034 36000
rect 58162 58248 58218 58304
rect 58162 57704 58218 57760
rect 58162 57160 58218 57216
rect 58162 56616 58218 56672
rect 58346 56108 58348 56128
rect 58348 56108 58400 56128
rect 58400 56108 58402 56128
rect 58346 56072 58402 56108
rect 58346 54440 58402 54496
rect 58346 52844 58348 52864
rect 58348 52844 58400 52864
rect 58400 52844 58402 52864
rect 58346 52808 58402 52844
rect 58346 51176 58402 51232
rect 58162 43016 58218 43072
rect 58162 40296 58218 40352
rect 58162 36488 58218 36544
rect 58162 34856 58218 34912
rect 57978 34312 58034 34368
rect 58162 33224 58218 33280
rect 58162 31592 58218 31648
rect 57978 31048 58034 31104
rect 57978 27784 58034 27840
rect 58162 29960 58218 30016
rect 58162 28328 58218 28384
rect 58162 26696 58218 26752
rect 58070 26152 58126 26208
rect 58162 25064 58218 25120
rect 58070 24520 58126 24576
rect 58162 23432 58218 23488
rect 58070 22888 58126 22944
rect 58162 21800 58218 21856
rect 58162 20168 58218 20224
rect 57242 18808 57298 18864
rect 58162 18536 58218 18592
rect 57058 17992 57114 18048
rect 57334 16904 57390 16960
rect 57978 16360 58034 16416
rect 57242 15272 57298 15328
rect 57978 14728 58034 14784
rect 58070 14456 58126 14512
rect 57334 13640 57390 13696
rect 57978 13096 58034 13152
rect 57242 12008 57298 12064
rect 57150 11464 57206 11520
rect 57058 9832 57114 9888
rect 56230 8200 56286 8256
rect 58162 10376 58218 10432
rect 57334 8744 57390 8800
rect 56414 7112 56470 7168
rect 57978 6568 58034 6624
rect 57242 5480 57298 5536
rect 58070 4936 58126 4992
rect 58070 3848 58126 3904
rect 58162 3304 58218 3360
rect 58162 2760 58218 2816
rect 57334 2216 57390 2272
rect 56506 1672 56562 1728
rect 56506 1128 56562 1184
<< metal3 >>
rect 56041 62658 56107 62661
rect 59200 62658 60000 62688
rect 56041 62656 60000 62658
rect 56041 62600 56046 62656
rect 56102 62600 60000 62656
rect 56041 62598 60000 62600
rect 56041 62595 56107 62598
rect 59200 62568 60000 62598
rect 56133 62114 56199 62117
rect 59200 62114 60000 62144
rect 56133 62112 60000 62114
rect 56133 62056 56138 62112
rect 56194 62056 60000 62112
rect 56133 62054 60000 62056
rect 56133 62051 56199 62054
rect 59200 62024 60000 62054
rect 0 61570 800 61600
rect 2773 61570 2839 61573
rect 0 61568 2839 61570
rect 0 61512 2778 61568
rect 2834 61512 2839 61568
rect 0 61510 2839 61512
rect 0 61480 800 61510
rect 2773 61507 2839 61510
rect 56501 61570 56567 61573
rect 59200 61570 60000 61600
rect 56501 61568 60000 61570
rect 56501 61512 56506 61568
rect 56562 61512 60000 61568
rect 56501 61510 60000 61512
rect 56501 61507 56567 61510
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 34930 61504 35246 61505
rect 34930 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35246 61504
rect 59200 61480 60000 61510
rect 34930 61439 35246 61440
rect 7833 61162 7899 61165
rect 30966 61162 30972 61164
rect 7833 61160 30972 61162
rect 7833 61104 7838 61160
rect 7894 61104 30972 61160
rect 7833 61102 30972 61104
rect 7833 61099 7899 61102
rect 30966 61100 30972 61102
rect 31036 61100 31042 61164
rect 56133 61026 56199 61029
rect 59200 61026 60000 61056
rect 56133 61024 60000 61026
rect 56133 60968 56138 61024
rect 56194 60968 60000 61024
rect 56133 60966 60000 60968
rect 56133 60963 56199 60966
rect 19570 60960 19886 60961
rect 0 60890 800 60920
rect 19570 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19886 60960
rect 19570 60895 19886 60896
rect 50290 60960 50606 60961
rect 50290 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50606 60960
rect 59200 60936 60000 60966
rect 50290 60895 50606 60896
rect 1669 60890 1735 60893
rect 0 60888 1735 60890
rect 0 60832 1674 60888
rect 1730 60832 1735 60888
rect 0 60830 1735 60832
rect 0 60800 800 60830
rect 1669 60827 1735 60830
rect 32070 60828 32076 60892
rect 32140 60890 32146 60892
rect 33317 60890 33383 60893
rect 32140 60888 33383 60890
rect 32140 60832 33322 60888
rect 33378 60832 33383 60888
rect 32140 60830 33383 60832
rect 32140 60828 32146 60830
rect 33317 60827 33383 60830
rect 33225 60756 33291 60757
rect 33174 60754 33180 60756
rect 33134 60694 33180 60754
rect 33244 60752 33291 60756
rect 33286 60696 33291 60752
rect 33174 60692 33180 60694
rect 33244 60692 33291 60696
rect 34646 60692 34652 60756
rect 34716 60754 34722 60756
rect 35065 60754 35131 60757
rect 34716 60752 35131 60754
rect 34716 60696 35070 60752
rect 35126 60696 35131 60752
rect 34716 60694 35131 60696
rect 34716 60692 34722 60694
rect 33225 60691 33291 60692
rect 35065 60691 35131 60694
rect 57329 60482 57395 60485
rect 59200 60482 60000 60512
rect 57329 60480 60000 60482
rect 57329 60424 57334 60480
rect 57390 60424 60000 60480
rect 57329 60422 60000 60424
rect 57329 60419 57395 60422
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 34930 60416 35246 60417
rect 34930 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35246 60416
rect 59200 60392 60000 60422
rect 34930 60351 35246 60352
rect 0 60210 800 60240
rect 1669 60210 1735 60213
rect 0 60208 1735 60210
rect 0 60152 1674 60208
rect 1730 60152 1735 60208
rect 0 60150 1735 60152
rect 0 60120 800 60150
rect 1669 60147 1735 60150
rect 57973 59938 58039 59941
rect 59200 59938 60000 59968
rect 57973 59936 60000 59938
rect 57973 59880 57978 59936
rect 58034 59880 60000 59936
rect 57973 59878 60000 59880
rect 57973 59875 58039 59878
rect 19570 59872 19886 59873
rect 19570 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19886 59872
rect 19570 59807 19886 59808
rect 50290 59872 50606 59873
rect 50290 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50606 59872
rect 59200 59848 60000 59878
rect 50290 59807 50606 59808
rect 0 59530 800 59560
rect 1577 59530 1643 59533
rect 0 59528 1643 59530
rect 0 59472 1582 59528
rect 1638 59472 1643 59528
rect 0 59470 1643 59472
rect 0 59440 800 59470
rect 1577 59467 1643 59470
rect 57789 59394 57855 59397
rect 59200 59394 60000 59424
rect 57789 59392 60000 59394
rect 57789 59336 57794 59392
rect 57850 59336 60000 59392
rect 57789 59334 60000 59336
rect 57789 59331 57855 59334
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 34930 59328 35246 59329
rect 34930 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35246 59328
rect 59200 59304 60000 59334
rect 34930 59263 35246 59264
rect 0 58850 800 58880
rect 1577 58850 1643 58853
rect 0 58848 1643 58850
rect 0 58792 1582 58848
rect 1638 58792 1643 58848
rect 0 58790 1643 58792
rect 0 58760 800 58790
rect 1577 58787 1643 58790
rect 57881 58850 57947 58853
rect 59200 58850 60000 58880
rect 57881 58848 60000 58850
rect 57881 58792 57886 58848
rect 57942 58792 60000 58848
rect 57881 58790 60000 58792
rect 57881 58787 57947 58790
rect 19570 58784 19886 58785
rect 19570 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19886 58784
rect 19570 58719 19886 58720
rect 50290 58784 50606 58785
rect 50290 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50606 58784
rect 59200 58760 60000 58790
rect 50290 58719 50606 58720
rect 16757 58578 16823 58581
rect 17401 58578 17467 58581
rect 16757 58576 17467 58578
rect 16757 58520 16762 58576
rect 16818 58520 17406 58576
rect 17462 58520 17467 58576
rect 16757 58518 17467 58520
rect 16757 58515 16823 58518
rect 17401 58515 17467 58518
rect 58157 58306 58223 58309
rect 59200 58306 60000 58336
rect 58157 58304 60000 58306
rect 58157 58248 58162 58304
rect 58218 58248 60000 58304
rect 58157 58246 60000 58248
rect 58157 58243 58223 58246
rect 4210 58240 4526 58241
rect 0 58170 800 58200
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 34930 58240 35246 58241
rect 34930 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35246 58240
rect 59200 58216 60000 58246
rect 34930 58175 35246 58176
rect 1669 58170 1735 58173
rect 0 58168 1735 58170
rect 0 58112 1674 58168
rect 1730 58112 1735 58168
rect 0 58110 1735 58112
rect 0 58080 800 58110
rect 1669 58107 1735 58110
rect 58157 57762 58223 57765
rect 59200 57762 60000 57792
rect 58157 57760 60000 57762
rect 58157 57704 58162 57760
rect 58218 57704 60000 57760
rect 58157 57702 60000 57704
rect 58157 57699 58223 57702
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 59200 57672 60000 57702
rect 50290 57631 50606 57632
rect 0 57490 800 57520
rect 1577 57490 1643 57493
rect 0 57488 1643 57490
rect 0 57432 1582 57488
rect 1638 57432 1643 57488
rect 0 57430 1643 57432
rect 0 57400 800 57430
rect 1577 57427 1643 57430
rect 38101 57356 38167 57357
rect 38101 57354 38148 57356
rect 38056 57352 38148 57354
rect 38056 57296 38106 57352
rect 38056 57294 38148 57296
rect 38101 57292 38148 57294
rect 38212 57292 38218 57356
rect 38101 57291 38167 57292
rect 58157 57218 58223 57221
rect 59200 57218 60000 57248
rect 58157 57216 60000 57218
rect 58157 57160 58162 57216
rect 58218 57160 60000 57216
rect 58157 57158 60000 57160
rect 58157 57155 58223 57158
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 59200 57128 60000 57158
rect 34930 57087 35246 57088
rect 0 56810 800 56840
rect 1669 56810 1735 56813
rect 0 56808 1735 56810
rect 0 56752 1674 56808
rect 1730 56752 1735 56808
rect 0 56750 1735 56752
rect 0 56720 800 56750
rect 1669 56747 1735 56750
rect 35341 56674 35407 56677
rect 35566 56674 35572 56676
rect 35341 56672 35572 56674
rect 35341 56616 35346 56672
rect 35402 56616 35572 56672
rect 35341 56614 35572 56616
rect 35341 56611 35407 56614
rect 35566 56612 35572 56614
rect 35636 56612 35642 56676
rect 58157 56674 58223 56677
rect 59200 56674 60000 56704
rect 58157 56672 60000 56674
rect 58157 56616 58162 56672
rect 58218 56616 60000 56672
rect 58157 56614 60000 56616
rect 58157 56611 58223 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 59200 56584 60000 56614
rect 50290 56543 50606 56544
rect 0 56130 800 56160
rect 1669 56130 1735 56133
rect 0 56128 1735 56130
rect 0 56072 1674 56128
rect 1730 56072 1735 56128
rect 0 56070 1735 56072
rect 0 56040 800 56070
rect 1669 56067 1735 56070
rect 58341 56130 58407 56133
rect 59200 56130 60000 56160
rect 58341 56128 60000 56130
rect 58341 56072 58346 56128
rect 58402 56072 60000 56128
rect 58341 56070 60000 56072
rect 58341 56067 58407 56070
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 59200 56040 60000 56070
rect 34930 55999 35246 56000
rect 19570 55520 19886 55521
rect 0 55450 800 55480
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 59200 55496 60000 55616
rect 50290 55455 50606 55456
rect 1669 55450 1735 55453
rect 0 55448 1735 55450
rect 0 55392 1674 55448
rect 1730 55392 1735 55448
rect 0 55390 1735 55392
rect 0 55360 800 55390
rect 1669 55387 1735 55390
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 59200 54952 60000 55072
rect 34930 54911 35246 54912
rect 0 54770 800 54800
rect 1577 54770 1643 54773
rect 0 54768 1643 54770
rect 0 54712 1582 54768
rect 1638 54712 1643 54768
rect 0 54710 1643 54712
rect 0 54680 800 54710
rect 1577 54707 1643 54710
rect 58341 54498 58407 54501
rect 59200 54498 60000 54528
rect 58341 54496 60000 54498
rect 58341 54440 58346 54496
rect 58402 54440 60000 54496
rect 58341 54438 60000 54440
rect 58341 54435 58407 54438
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 59200 54408 60000 54438
rect 50290 54367 50606 54368
rect 0 54090 800 54120
rect 1669 54090 1735 54093
rect 0 54088 1735 54090
rect 0 54032 1674 54088
rect 1730 54032 1735 54088
rect 0 54030 1735 54032
rect 0 54000 800 54030
rect 1669 54027 1735 54030
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 59200 53864 60000 53984
rect 34930 53823 35246 53824
rect 0 53410 800 53440
rect 1577 53410 1643 53413
rect 0 53408 1643 53410
rect 0 53352 1582 53408
rect 1638 53352 1643 53408
rect 0 53350 1643 53352
rect 0 53320 800 53350
rect 1577 53347 1643 53350
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 59200 53320 60000 53440
rect 50290 53279 50606 53280
rect 18270 53076 18276 53140
rect 18340 53138 18346 53140
rect 42057 53138 42123 53141
rect 18340 53136 42123 53138
rect 18340 53080 42062 53136
rect 42118 53080 42123 53136
rect 18340 53078 42123 53080
rect 18340 53076 18346 53078
rect 42057 53075 42123 53078
rect 58341 52866 58407 52869
rect 59200 52866 60000 52896
rect 58341 52864 60000 52866
rect 58341 52808 58346 52864
rect 58402 52808 60000 52864
rect 58341 52806 60000 52808
rect 58341 52803 58407 52806
rect 4210 52800 4526 52801
rect 0 52730 800 52760
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 59200 52776 60000 52806
rect 34930 52735 35246 52736
rect 1577 52730 1643 52733
rect 0 52728 1643 52730
rect 0 52672 1582 52728
rect 1638 52672 1643 52728
rect 0 52670 1643 52672
rect 0 52640 800 52670
rect 1577 52667 1643 52670
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 59200 52232 60000 52352
rect 50290 52191 50606 52192
rect 0 52050 800 52080
rect 1669 52050 1735 52053
rect 0 52048 1735 52050
rect 0 51992 1674 52048
rect 1730 51992 1735 52048
rect 0 51990 1735 51992
rect 0 51960 800 51990
rect 1669 51987 1735 51990
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 59200 51688 60000 51808
rect 34930 51647 35246 51648
rect 0 51370 800 51400
rect 1669 51370 1735 51373
rect 0 51368 1735 51370
rect 0 51312 1674 51368
rect 1730 51312 1735 51368
rect 0 51310 1735 51312
rect 0 51280 800 51310
rect 1669 51307 1735 51310
rect 58341 51234 58407 51237
rect 59200 51234 60000 51264
rect 58341 51232 60000 51234
rect 58341 51176 58346 51232
rect 58402 51176 60000 51232
rect 58341 51174 60000 51176
rect 58341 51171 58407 51174
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 59200 51144 60000 51174
rect 50290 51103 50606 51104
rect 0 50690 800 50720
rect 1669 50690 1735 50693
rect 0 50688 1735 50690
rect 0 50632 1674 50688
rect 1730 50632 1735 50688
rect 0 50630 1735 50632
rect 0 50600 800 50630
rect 1669 50627 1735 50630
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 59200 50600 60000 50720
rect 34930 50559 35246 50560
rect 19570 50080 19886 50081
rect 0 50010 800 50040
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 59200 50056 60000 50176
rect 50290 50015 50606 50016
rect 1669 50010 1735 50013
rect 0 50008 1735 50010
rect 0 49952 1674 50008
rect 1730 49952 1735 50008
rect 0 49950 1735 49952
rect 0 49920 800 49950
rect 1669 49947 1735 49950
rect 57881 49602 57947 49605
rect 59200 49602 60000 49632
rect 57881 49600 60000 49602
rect 57881 49544 57886 49600
rect 57942 49544 60000 49600
rect 57881 49542 60000 49544
rect 57881 49539 57947 49542
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 59200 49512 60000 49542
rect 34930 49471 35246 49472
rect 0 49330 800 49360
rect 1669 49330 1735 49333
rect 0 49328 1735 49330
rect 0 49272 1674 49328
rect 1730 49272 1735 49328
rect 0 49270 1735 49272
rect 0 49240 800 49270
rect 1669 49267 1735 49270
rect 57973 49058 58039 49061
rect 59200 49058 60000 49088
rect 57973 49056 60000 49058
rect 57973 49000 57978 49056
rect 58034 49000 60000 49056
rect 57973 48998 60000 49000
rect 57973 48995 58039 48998
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 59200 48968 60000 48998
rect 50290 48927 50606 48928
rect 0 48650 800 48680
rect 1669 48650 1735 48653
rect 0 48648 1735 48650
rect 0 48592 1674 48648
rect 1730 48592 1735 48648
rect 0 48590 1735 48592
rect 0 48560 800 48590
rect 1669 48587 1735 48590
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 59200 48424 60000 48544
rect 34930 48383 35246 48384
rect 0 47970 800 48000
rect 1669 47970 1735 47973
rect 0 47968 1735 47970
rect 0 47912 1674 47968
rect 1730 47912 1735 47968
rect 0 47910 1735 47912
rect 0 47880 800 47910
rect 1669 47907 1735 47910
rect 57329 47970 57395 47973
rect 59200 47970 60000 48000
rect 57329 47968 60000 47970
rect 57329 47912 57334 47968
rect 57390 47912 60000 47968
rect 57329 47910 60000 47912
rect 57329 47907 57395 47910
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 59200 47880 60000 47910
rect 50290 47839 50606 47840
rect 57973 47426 58039 47429
rect 59200 47426 60000 47456
rect 57973 47424 60000 47426
rect 57973 47368 57978 47424
rect 58034 47368 60000 47424
rect 57973 47366 60000 47368
rect 57973 47363 58039 47366
rect 4210 47360 4526 47361
rect 0 47290 800 47320
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 59200 47336 60000 47366
rect 34930 47295 35246 47296
rect 1669 47290 1735 47293
rect 0 47288 1735 47290
rect 0 47232 1674 47288
rect 1730 47232 1735 47288
rect 0 47230 1735 47232
rect 0 47200 800 47230
rect 1669 47227 1735 47230
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 59200 46792 60000 46912
rect 50290 46751 50606 46752
rect 0 46610 800 46640
rect 1669 46610 1735 46613
rect 0 46608 1735 46610
rect 0 46552 1674 46608
rect 1730 46552 1735 46608
rect 0 46550 1735 46552
rect 0 46520 800 46550
rect 1669 46547 1735 46550
rect 57881 46338 57947 46341
rect 59200 46338 60000 46368
rect 57881 46336 60000 46338
rect 57881 46280 57886 46336
rect 57942 46280 60000 46336
rect 57881 46278 60000 46280
rect 57881 46275 57947 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 59200 46248 60000 46278
rect 34930 46207 35246 46208
rect 0 45930 800 45960
rect 1669 45930 1735 45933
rect 0 45928 1735 45930
rect 0 45872 1674 45928
rect 1730 45872 1735 45928
rect 0 45870 1735 45872
rect 0 45840 800 45870
rect 1669 45867 1735 45870
rect 57973 45794 58039 45797
rect 59200 45794 60000 45824
rect 57973 45792 60000 45794
rect 57973 45736 57978 45792
rect 58034 45736 60000 45792
rect 57973 45734 60000 45736
rect 57973 45731 58039 45734
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 59200 45704 60000 45734
rect 50290 45663 50606 45664
rect 0 45250 800 45280
rect 1577 45250 1643 45253
rect 0 45248 1643 45250
rect 0 45192 1582 45248
rect 1638 45192 1643 45248
rect 0 45190 1643 45192
rect 0 45160 800 45190
rect 1577 45187 1643 45190
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 59200 45160 60000 45280
rect 34930 45119 35246 45120
rect 57237 44706 57303 44709
rect 59200 44706 60000 44736
rect 57237 44704 60000 44706
rect 57237 44648 57242 44704
rect 57298 44648 60000 44704
rect 57237 44646 60000 44648
rect 57237 44643 57303 44646
rect 19570 44640 19886 44641
rect 0 44570 800 44600
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 59200 44616 60000 44646
rect 50290 44575 50606 44576
rect 1669 44570 1735 44573
rect 0 44568 1735 44570
rect 0 44512 1674 44568
rect 1730 44512 1735 44568
rect 0 44510 1735 44512
rect 0 44480 800 44510
rect 1669 44507 1735 44510
rect 57881 44162 57947 44165
rect 59200 44162 60000 44192
rect 57881 44160 60000 44162
rect 57881 44104 57886 44160
rect 57942 44104 60000 44160
rect 57881 44102 60000 44104
rect 57881 44099 57947 44102
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 59200 44072 60000 44102
rect 34930 44031 35246 44032
rect 0 43890 800 43920
rect 1669 43890 1735 43893
rect 0 43888 1735 43890
rect 0 43832 1674 43888
rect 1730 43832 1735 43888
rect 0 43830 1735 43832
rect 0 43800 800 43830
rect 1669 43827 1735 43830
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 59200 43528 60000 43648
rect 50290 43487 50606 43488
rect 0 43210 800 43240
rect 1577 43210 1643 43213
rect 0 43208 1643 43210
rect 0 43152 1582 43208
rect 1638 43152 1643 43208
rect 0 43150 1643 43152
rect 0 43120 800 43150
rect 1577 43147 1643 43150
rect 58157 43074 58223 43077
rect 59200 43074 60000 43104
rect 58157 43072 60000 43074
rect 58157 43016 58162 43072
rect 58218 43016 60000 43072
rect 58157 43014 60000 43016
rect 58157 43011 58223 43014
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 59200 42984 60000 43014
rect 34930 42943 35246 42944
rect 0 42530 800 42560
rect 1669 42530 1735 42533
rect 0 42528 1735 42530
rect 0 42472 1674 42528
rect 1730 42472 1735 42528
rect 0 42470 1735 42472
rect 0 42440 800 42470
rect 1669 42467 1735 42470
rect 56961 42530 57027 42533
rect 59200 42530 60000 42560
rect 56961 42528 60000 42530
rect 56961 42472 56966 42528
rect 57022 42472 60000 42528
rect 56961 42470 60000 42472
rect 56961 42467 57027 42470
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 59200 42440 60000 42470
rect 50290 42399 50606 42400
rect 57881 41986 57947 41989
rect 59200 41986 60000 42016
rect 57881 41984 60000 41986
rect 57881 41928 57886 41984
rect 57942 41928 60000 41984
rect 57881 41926 60000 41928
rect 57881 41923 57947 41926
rect 4210 41920 4526 41921
rect 0 41850 800 41880
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 59200 41896 60000 41926
rect 34930 41855 35246 41856
rect 1669 41850 1735 41853
rect 0 41848 1735 41850
rect 0 41792 1674 41848
rect 1730 41792 1735 41848
rect 0 41790 1735 41792
rect 0 41760 800 41790
rect 1669 41787 1735 41790
rect 57237 41442 57303 41445
rect 59200 41442 60000 41472
rect 57237 41440 60000 41442
rect 57237 41384 57242 41440
rect 57298 41384 60000 41440
rect 57237 41382 60000 41384
rect 57237 41379 57303 41382
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 59200 41352 60000 41382
rect 50290 41311 50606 41312
rect 0 41170 800 41200
rect 1669 41170 1735 41173
rect 0 41168 1735 41170
rect 0 41112 1674 41168
rect 1730 41112 1735 41168
rect 0 41110 1735 41112
rect 0 41080 800 41110
rect 1669 41107 1735 41110
rect 57881 40898 57947 40901
rect 59200 40898 60000 40928
rect 57881 40896 60000 40898
rect 57881 40840 57886 40896
rect 57942 40840 60000 40896
rect 57881 40838 60000 40840
rect 57881 40835 57947 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 59200 40808 60000 40838
rect 34930 40767 35246 40768
rect 0 40490 800 40520
rect 1393 40490 1459 40493
rect 0 40488 1459 40490
rect 0 40432 1398 40488
rect 1454 40432 1459 40488
rect 0 40430 1459 40432
rect 0 40400 800 40430
rect 1393 40427 1459 40430
rect 58157 40354 58223 40357
rect 59200 40354 60000 40384
rect 58157 40352 60000 40354
rect 58157 40296 58162 40352
rect 58218 40296 60000 40352
rect 58157 40294 60000 40296
rect 58157 40291 58223 40294
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 59200 40264 60000 40294
rect 50290 40223 50606 40224
rect 0 39810 800 39840
rect 1669 39810 1735 39813
rect 0 39808 1735 39810
rect 0 39752 1674 39808
rect 1730 39752 1735 39808
rect 0 39750 1735 39752
rect 0 39720 800 39750
rect 1669 39747 1735 39750
rect 57881 39810 57947 39813
rect 59200 39810 60000 39840
rect 57881 39808 60000 39810
rect 57881 39752 57886 39808
rect 57942 39752 60000 39808
rect 57881 39750 60000 39752
rect 57881 39747 57947 39750
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 59200 39720 60000 39750
rect 34930 39679 35246 39680
rect 57053 39266 57119 39269
rect 59200 39266 60000 39296
rect 57053 39264 60000 39266
rect 57053 39208 57058 39264
rect 57114 39208 60000 39264
rect 57053 39206 60000 39208
rect 57053 39203 57119 39206
rect 19570 39200 19886 39201
rect 0 39130 800 39160
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 59200 39176 60000 39206
rect 50290 39135 50606 39136
rect 1577 39130 1643 39133
rect 0 39128 1643 39130
rect 0 39072 1582 39128
rect 1638 39072 1643 39128
rect 0 39070 1643 39072
rect 0 39040 800 39070
rect 1577 39067 1643 39070
rect 27521 38722 27587 38725
rect 28758 38722 28764 38724
rect 27521 38720 28764 38722
rect 27521 38664 27526 38720
rect 27582 38664 28764 38720
rect 27521 38662 28764 38664
rect 27521 38659 27587 38662
rect 28758 38660 28764 38662
rect 28828 38660 28834 38724
rect 57973 38722 58039 38725
rect 59200 38722 60000 38752
rect 57973 38720 60000 38722
rect 57973 38664 57978 38720
rect 58034 38664 60000 38720
rect 57973 38662 60000 38664
rect 57973 38659 58039 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 59200 38632 60000 38662
rect 34930 38591 35246 38592
rect 0 38450 800 38480
rect 1393 38450 1459 38453
rect 0 38448 1459 38450
rect 0 38392 1398 38448
rect 1454 38392 1459 38448
rect 0 38390 1459 38392
rect 0 38360 800 38390
rect 1393 38387 1459 38390
rect 57237 38178 57303 38181
rect 59200 38178 60000 38208
rect 57237 38176 60000 38178
rect 57237 38120 57242 38176
rect 57298 38120 60000 38176
rect 57237 38118 60000 38120
rect 57237 38115 57303 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 59200 38088 60000 38118
rect 50290 38047 50606 38048
rect 0 37770 800 37800
rect 1669 37770 1735 37773
rect 0 37768 1735 37770
rect 0 37712 1674 37768
rect 1730 37712 1735 37768
rect 0 37710 1735 37712
rect 0 37680 800 37710
rect 1669 37707 1735 37710
rect 19701 37770 19767 37773
rect 20110 37770 20116 37772
rect 19701 37768 20116 37770
rect 19701 37712 19706 37768
rect 19762 37712 20116 37768
rect 19701 37710 20116 37712
rect 19701 37707 19767 37710
rect 20110 37708 20116 37710
rect 20180 37708 20186 37772
rect 57881 37634 57947 37637
rect 59200 37634 60000 37664
rect 57881 37632 60000 37634
rect 57881 37576 57886 37632
rect 57942 37576 60000 37632
rect 57881 37574 60000 37576
rect 57881 37571 57947 37574
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 59200 37544 60000 37574
rect 34930 37503 35246 37504
rect 0 37090 800 37120
rect 2405 37090 2471 37093
rect 0 37088 2471 37090
rect 0 37032 2410 37088
rect 2466 37032 2471 37088
rect 0 37030 2471 37032
rect 0 37000 800 37030
rect 2405 37027 2471 37030
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 59200 37000 60000 37120
rect 50290 36959 50606 36960
rect 58157 36546 58223 36549
rect 59200 36546 60000 36576
rect 58157 36544 60000 36546
rect 58157 36488 58162 36544
rect 58218 36488 60000 36544
rect 58157 36486 60000 36488
rect 58157 36483 58223 36486
rect 4210 36480 4526 36481
rect 0 36410 800 36440
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 59200 36456 60000 36486
rect 34930 36415 35246 36416
rect 1577 36410 1643 36413
rect 0 36408 1643 36410
rect 0 36352 1582 36408
rect 1638 36352 1643 36408
rect 0 36350 1643 36352
rect 0 36320 800 36350
rect 1577 36347 1643 36350
rect 20110 36076 20116 36140
rect 20180 36138 20186 36140
rect 24761 36138 24827 36141
rect 20180 36136 24827 36138
rect 20180 36080 24766 36136
rect 24822 36080 24827 36136
rect 20180 36078 24827 36080
rect 20180 36076 20186 36078
rect 24761 36075 24827 36078
rect 57973 36002 58039 36005
rect 59200 36002 60000 36032
rect 57973 36000 60000 36002
rect 57973 35944 57978 36000
rect 58034 35944 60000 36000
rect 57973 35942 60000 35944
rect 57973 35939 58039 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 59200 35912 60000 35942
rect 50290 35871 50606 35872
rect 0 35730 800 35760
rect 1393 35730 1459 35733
rect 0 35728 1459 35730
rect 0 35672 1398 35728
rect 1454 35672 1459 35728
rect 0 35670 1459 35672
rect 0 35640 800 35670
rect 1393 35667 1459 35670
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 59200 35368 60000 35488
rect 34930 35327 35246 35328
rect 22921 35322 22987 35325
rect 25221 35322 25287 35325
rect 22921 35320 25287 35322
rect 22921 35264 22926 35320
rect 22982 35264 25226 35320
rect 25282 35264 25287 35320
rect 22921 35262 25287 35264
rect 22921 35259 22987 35262
rect 25221 35259 25287 35262
rect 0 35050 800 35080
rect 1669 35050 1735 35053
rect 0 35048 1735 35050
rect 0 34992 1674 35048
rect 1730 34992 1735 35048
rect 0 34990 1735 34992
rect 0 34960 800 34990
rect 1669 34987 1735 34990
rect 24117 35050 24183 35053
rect 25497 35050 25563 35053
rect 24117 35048 25563 35050
rect 24117 34992 24122 35048
rect 24178 34992 25502 35048
rect 25558 34992 25563 35048
rect 24117 34990 25563 34992
rect 24117 34987 24183 34990
rect 25497 34987 25563 34990
rect 58157 34914 58223 34917
rect 59200 34914 60000 34944
rect 58157 34912 60000 34914
rect 58157 34856 58162 34912
rect 58218 34856 60000 34912
rect 58157 34854 60000 34856
rect 58157 34851 58223 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 59200 34824 60000 34854
rect 50290 34783 50606 34784
rect 0 34370 800 34400
rect 1669 34370 1735 34373
rect 0 34368 1735 34370
rect 0 34312 1674 34368
rect 1730 34312 1735 34368
rect 0 34310 1735 34312
rect 0 34280 800 34310
rect 1669 34307 1735 34310
rect 57973 34370 58039 34373
rect 59200 34370 60000 34400
rect 57973 34368 60000 34370
rect 57973 34312 57978 34368
rect 58034 34312 60000 34368
rect 57973 34310 60000 34312
rect 57973 34307 58039 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 59200 34280 60000 34310
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 0 33690 800 33720
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 59200 33736 60000 33856
rect 50290 33695 50606 33696
rect 1669 33690 1735 33693
rect 0 33688 1735 33690
rect 0 33632 1674 33688
rect 1730 33632 1735 33688
rect 0 33630 1735 33632
rect 0 33600 800 33630
rect 1669 33627 1735 33630
rect 58157 33282 58223 33285
rect 59200 33282 60000 33312
rect 58157 33280 60000 33282
rect 58157 33224 58162 33280
rect 58218 33224 60000 33280
rect 58157 33222 60000 33224
rect 58157 33219 58223 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 59200 33192 60000 33222
rect 34930 33151 35246 33152
rect 19517 33146 19583 33149
rect 20069 33146 20135 33149
rect 19517 33144 20135 33146
rect 19517 33088 19522 33144
rect 19578 33088 20074 33144
rect 20130 33088 20135 33144
rect 19517 33086 20135 33088
rect 19517 33083 19583 33086
rect 20069 33083 20135 33086
rect 0 33010 800 33040
rect 1669 33010 1735 33013
rect 0 33008 1735 33010
rect 0 32952 1674 33008
rect 1730 32952 1735 33008
rect 0 32950 1735 32952
rect 0 32920 800 32950
rect 1669 32947 1735 32950
rect 19609 33010 19675 33013
rect 19885 33010 19951 33013
rect 20345 33010 20411 33013
rect 19609 33008 20411 33010
rect 19609 32952 19614 33008
rect 19670 32952 19890 33008
rect 19946 32952 20350 33008
rect 20406 32952 20411 33008
rect 19609 32950 20411 32952
rect 19609 32947 19675 32950
rect 19885 32947 19951 32950
rect 20345 32947 20411 32950
rect 21173 32874 21239 32877
rect 19382 32872 21239 32874
rect 19382 32816 21178 32872
rect 21234 32816 21239 32872
rect 19382 32814 21239 32816
rect 19382 32741 19442 32814
rect 21173 32811 21239 32814
rect 19333 32736 19442 32741
rect 19333 32680 19338 32736
rect 19394 32680 19442 32736
rect 19333 32678 19442 32680
rect 57053 32738 57119 32741
rect 59200 32738 60000 32768
rect 57053 32736 60000 32738
rect 57053 32680 57058 32736
rect 57114 32680 60000 32736
rect 57053 32678 60000 32680
rect 19333 32675 19399 32678
rect 57053 32675 57119 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 59200 32648 60000 32678
rect 50290 32607 50606 32608
rect 0 32330 800 32360
rect 1669 32330 1735 32333
rect 0 32328 1735 32330
rect 0 32272 1674 32328
rect 1730 32272 1735 32328
rect 0 32270 1735 32272
rect 0 32240 800 32270
rect 1669 32267 1735 32270
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 59200 32104 60000 32224
rect 34930 32063 35246 32064
rect 19793 32058 19859 32061
rect 20897 32058 20963 32061
rect 19793 32056 20963 32058
rect 19793 32000 19798 32056
rect 19854 32000 20902 32056
rect 20958 32000 20963 32056
rect 19793 31998 20963 32000
rect 19793 31995 19859 31998
rect 20897 31995 20963 31998
rect 0 31650 800 31680
rect 1669 31650 1735 31653
rect 0 31648 1735 31650
rect 0 31592 1674 31648
rect 1730 31592 1735 31648
rect 0 31590 1735 31592
rect 0 31560 800 31590
rect 1669 31587 1735 31590
rect 58157 31650 58223 31653
rect 59200 31650 60000 31680
rect 58157 31648 60000 31650
rect 58157 31592 58162 31648
rect 58218 31592 60000 31648
rect 58157 31590 60000 31592
rect 58157 31587 58223 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 59200 31560 60000 31590
rect 50290 31519 50606 31520
rect 35157 31242 35223 31245
rect 35709 31242 35775 31245
rect 35157 31240 35775 31242
rect 35157 31184 35162 31240
rect 35218 31184 35714 31240
rect 35770 31184 35775 31240
rect 35157 31182 35775 31184
rect 35157 31179 35223 31182
rect 35709 31179 35775 31182
rect 57973 31106 58039 31109
rect 59200 31106 60000 31136
rect 57973 31104 60000 31106
rect 57973 31048 57978 31104
rect 58034 31048 60000 31104
rect 57973 31046 60000 31048
rect 57973 31043 58039 31046
rect 4210 31040 4526 31041
rect 0 30970 800 31000
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 59200 31016 60000 31046
rect 34930 30975 35246 30976
rect 1669 30970 1735 30973
rect 0 30968 1735 30970
rect 0 30912 1674 30968
rect 1730 30912 1735 30968
rect 0 30910 1735 30912
rect 0 30880 800 30910
rect 1669 30907 1735 30910
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 59200 30472 60000 30592
rect 50290 30431 50606 30432
rect 0 30290 800 30320
rect 1669 30290 1735 30293
rect 0 30288 1735 30290
rect 0 30232 1674 30288
rect 1730 30232 1735 30288
rect 0 30230 1735 30232
rect 0 30200 800 30230
rect 1669 30227 1735 30230
rect 26509 30154 26575 30157
rect 31886 30154 31892 30156
rect 26509 30152 31892 30154
rect 26509 30096 26514 30152
rect 26570 30096 31892 30152
rect 26509 30094 31892 30096
rect 26509 30091 26575 30094
rect 31886 30092 31892 30094
rect 31956 30092 31962 30156
rect 19977 30018 20043 30021
rect 20110 30018 20116 30020
rect 19977 30016 20116 30018
rect 19977 29960 19982 30016
rect 20038 29960 20116 30016
rect 19977 29958 20116 29960
rect 19977 29955 20043 29958
rect 20110 29956 20116 29958
rect 20180 29956 20186 30020
rect 58157 30018 58223 30021
rect 59200 30018 60000 30048
rect 58157 30016 60000 30018
rect 58157 29960 58162 30016
rect 58218 29960 60000 30016
rect 58157 29958 60000 29960
rect 58157 29955 58223 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 59200 29928 60000 29958
rect 34930 29887 35246 29888
rect 0 29610 800 29640
rect 1853 29610 1919 29613
rect 0 29608 1919 29610
rect 0 29552 1858 29608
rect 1914 29552 1919 29608
rect 0 29550 1919 29552
rect 0 29520 800 29550
rect 1853 29547 1919 29550
rect 57053 29474 57119 29477
rect 59200 29474 60000 29504
rect 57053 29472 60000 29474
rect 57053 29416 57058 29472
rect 57114 29416 60000 29472
rect 57053 29414 60000 29416
rect 57053 29411 57119 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 59200 29384 60000 29414
rect 50290 29343 50606 29344
rect 22737 29202 22803 29205
rect 28574 29202 28580 29204
rect 22737 29200 28580 29202
rect 22737 29144 22742 29200
rect 22798 29144 28580 29200
rect 22737 29142 28580 29144
rect 22737 29139 22803 29142
rect 28574 29140 28580 29142
rect 28644 29140 28650 29204
rect 24117 29068 24183 29069
rect 24117 29066 24164 29068
rect 24072 29064 24164 29066
rect 24072 29008 24122 29064
rect 24072 29006 24164 29008
rect 24117 29004 24164 29006
rect 24228 29004 24234 29068
rect 31518 29004 31524 29068
rect 31588 29066 31594 29068
rect 33133 29066 33199 29069
rect 31588 29064 33199 29066
rect 31588 29008 33138 29064
rect 33194 29008 33199 29064
rect 31588 29006 33199 29008
rect 31588 29004 31594 29006
rect 24117 29003 24183 29004
rect 33133 29003 33199 29006
rect 0 28930 800 28960
rect 1761 28930 1827 28933
rect 0 28928 1827 28930
rect 0 28872 1766 28928
rect 1822 28872 1827 28928
rect 0 28870 1827 28872
rect 0 28840 800 28870
rect 1761 28867 1827 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 59200 28840 60000 28960
rect 34930 28799 35246 28800
rect 58157 28386 58223 28389
rect 59200 28386 60000 28416
rect 58157 28384 60000 28386
rect 58157 28328 58162 28384
rect 58218 28328 60000 28384
rect 58157 28326 60000 28328
rect 58157 28323 58223 28326
rect 19570 28320 19886 28321
rect 0 28250 800 28280
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 59200 28296 60000 28326
rect 50290 28255 50606 28256
rect 1853 28250 1919 28253
rect 0 28248 1919 28250
rect 0 28192 1858 28248
rect 1914 28192 1919 28248
rect 0 28190 1919 28192
rect 0 28160 800 28190
rect 1853 28187 1919 28190
rect 57973 27842 58039 27845
rect 59200 27842 60000 27872
rect 57973 27840 60000 27842
rect 57973 27784 57978 27840
rect 58034 27784 60000 27840
rect 57973 27782 60000 27784
rect 57973 27779 58039 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 59200 27752 60000 27782
rect 34930 27711 35246 27712
rect 0 27570 800 27600
rect 1577 27570 1643 27573
rect 0 27568 1643 27570
rect 0 27512 1582 27568
rect 1638 27512 1643 27568
rect 0 27510 1643 27512
rect 0 27480 800 27510
rect 1577 27507 1643 27510
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 59200 27208 60000 27328
rect 50290 27167 50606 27168
rect 0 26890 800 26920
rect 1761 26890 1827 26893
rect 0 26888 1827 26890
rect 0 26832 1766 26888
rect 1822 26832 1827 26888
rect 0 26830 1827 26832
rect 0 26800 800 26830
rect 1761 26827 1827 26830
rect 58157 26754 58223 26757
rect 59200 26754 60000 26784
rect 58157 26752 60000 26754
rect 58157 26696 58162 26752
rect 58218 26696 60000 26752
rect 58157 26694 60000 26696
rect 58157 26691 58223 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 59200 26664 60000 26694
rect 34930 26623 35246 26624
rect 0 26210 800 26240
rect 1853 26210 1919 26213
rect 0 26208 1919 26210
rect 0 26152 1858 26208
rect 1914 26152 1919 26208
rect 0 26150 1919 26152
rect 0 26120 800 26150
rect 1853 26147 1919 26150
rect 58065 26210 58131 26213
rect 59200 26210 60000 26240
rect 58065 26208 60000 26210
rect 58065 26152 58070 26208
rect 58126 26152 60000 26208
rect 58065 26150 60000 26152
rect 58065 26147 58131 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 59200 26120 60000 26150
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 0 25530 800 25560
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 59200 25576 60000 25696
rect 34930 25535 35246 25536
rect 1761 25530 1827 25533
rect 0 25528 1827 25530
rect 0 25472 1766 25528
rect 1822 25472 1827 25528
rect 0 25470 1827 25472
rect 0 25440 800 25470
rect 1761 25467 1827 25470
rect 58157 25122 58223 25125
rect 59200 25122 60000 25152
rect 58157 25120 60000 25122
rect 58157 25064 58162 25120
rect 58218 25064 60000 25120
rect 58157 25062 60000 25064
rect 58157 25059 58223 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 59200 25032 60000 25062
rect 50290 24991 50606 24992
rect 0 24850 800 24880
rect 1853 24850 1919 24853
rect 0 24848 1919 24850
rect 0 24792 1858 24848
rect 1914 24792 1919 24848
rect 0 24790 1919 24792
rect 0 24760 800 24790
rect 1853 24787 1919 24790
rect 29494 24652 29500 24716
rect 29564 24714 29570 24716
rect 32581 24714 32647 24717
rect 29564 24712 32647 24714
rect 29564 24656 32586 24712
rect 32642 24656 32647 24712
rect 29564 24654 32647 24656
rect 29564 24652 29570 24654
rect 32581 24651 32647 24654
rect 58065 24578 58131 24581
rect 59200 24578 60000 24608
rect 58065 24576 60000 24578
rect 58065 24520 58070 24576
rect 58126 24520 60000 24576
rect 58065 24518 60000 24520
rect 58065 24515 58131 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 59200 24488 60000 24518
rect 34930 24447 35246 24448
rect 0 24170 800 24200
rect 1853 24170 1919 24173
rect 0 24168 1919 24170
rect 0 24112 1858 24168
rect 1914 24112 1919 24168
rect 0 24110 1919 24112
rect 0 24080 800 24110
rect 1853 24107 1919 24110
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 59200 23944 60000 24064
rect 50290 23903 50606 23904
rect 33961 23626 34027 23629
rect 35065 23626 35131 23629
rect 37549 23626 37615 23629
rect 33961 23624 37615 23626
rect 33961 23568 33966 23624
rect 34022 23568 35070 23624
rect 35126 23568 37554 23624
rect 37610 23568 37615 23624
rect 33961 23566 37615 23568
rect 33961 23563 34027 23566
rect 35065 23563 35131 23566
rect 37549 23563 37615 23566
rect 0 23490 800 23520
rect 1761 23490 1827 23493
rect 0 23488 1827 23490
rect 0 23432 1766 23488
rect 1822 23432 1827 23488
rect 0 23430 1827 23432
rect 0 23400 800 23430
rect 1761 23427 1827 23430
rect 58157 23490 58223 23493
rect 59200 23490 60000 23520
rect 58157 23488 60000 23490
rect 58157 23432 58162 23488
rect 58218 23432 60000 23488
rect 58157 23430 60000 23432
rect 58157 23427 58223 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 59200 23400 60000 23430
rect 34930 23359 35246 23360
rect 27153 23218 27219 23221
rect 42517 23218 42583 23221
rect 27153 23216 42583 23218
rect 27153 23160 27158 23216
rect 27214 23160 42522 23216
rect 42578 23160 42583 23216
rect 27153 23158 42583 23160
rect 27153 23155 27219 23158
rect 42517 23155 42583 23158
rect 29913 23082 29979 23085
rect 30373 23082 30439 23085
rect 29913 23080 30439 23082
rect 29913 23024 29918 23080
rect 29974 23024 30378 23080
rect 30434 23024 30439 23080
rect 29913 23022 30439 23024
rect 29913 23019 29979 23022
rect 30373 23019 30439 23022
rect 33869 23082 33935 23085
rect 36445 23082 36511 23085
rect 33869 23080 36511 23082
rect 33869 23024 33874 23080
rect 33930 23024 36450 23080
rect 36506 23024 36511 23080
rect 33869 23022 36511 23024
rect 33869 23019 33935 23022
rect 36445 23019 36511 23022
rect 38837 23082 38903 23085
rect 40677 23082 40743 23085
rect 38837 23080 40743 23082
rect 38837 23024 38842 23080
rect 38898 23024 40682 23080
rect 40738 23024 40743 23080
rect 38837 23022 40743 23024
rect 38837 23019 38903 23022
rect 40677 23019 40743 23022
rect 42793 23082 42859 23085
rect 43897 23082 43963 23085
rect 42793 23080 43963 23082
rect 42793 23024 42798 23080
rect 42854 23024 43902 23080
rect 43958 23024 43963 23080
rect 42793 23022 43963 23024
rect 42793 23019 42859 23022
rect 43897 23019 43963 23022
rect 26693 22946 26759 22949
rect 29637 22946 29703 22949
rect 35709 22946 35775 22949
rect 26693 22944 35775 22946
rect 26693 22888 26698 22944
rect 26754 22888 29642 22944
rect 29698 22888 35714 22944
rect 35770 22888 35775 22944
rect 26693 22886 35775 22888
rect 26693 22883 26759 22886
rect 29637 22883 29703 22886
rect 35709 22883 35775 22886
rect 39665 22946 39731 22949
rect 40217 22946 40283 22949
rect 39665 22944 40283 22946
rect 39665 22888 39670 22944
rect 39726 22888 40222 22944
rect 40278 22888 40283 22944
rect 39665 22886 40283 22888
rect 39665 22883 39731 22886
rect 40217 22883 40283 22886
rect 58065 22946 58131 22949
rect 59200 22946 60000 22976
rect 58065 22944 60000 22946
rect 58065 22888 58070 22944
rect 58126 22888 60000 22944
rect 58065 22886 60000 22888
rect 58065 22883 58131 22886
rect 19570 22880 19886 22881
rect 0 22810 800 22840
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 59200 22856 60000 22886
rect 50290 22815 50606 22816
rect 1853 22810 1919 22813
rect 0 22808 1919 22810
rect 0 22752 1858 22808
rect 1914 22752 1919 22808
rect 0 22750 1919 22752
rect 0 22720 800 22750
rect 1853 22747 1919 22750
rect 33593 22810 33659 22813
rect 36445 22810 36511 22813
rect 33593 22808 36511 22810
rect 33593 22752 33598 22808
rect 33654 22752 36450 22808
rect 36506 22752 36511 22808
rect 33593 22750 36511 22752
rect 33593 22747 33659 22750
rect 36445 22747 36511 22750
rect 34145 22674 34211 22677
rect 35709 22674 35775 22677
rect 34145 22672 35775 22674
rect 34145 22616 34150 22672
rect 34206 22616 35714 22672
rect 35770 22616 35775 22672
rect 34145 22614 35775 22616
rect 34145 22611 34211 22614
rect 35709 22611 35775 22614
rect 34145 22538 34211 22541
rect 35617 22538 35683 22541
rect 34145 22536 35683 22538
rect 34145 22480 34150 22536
rect 34206 22480 35622 22536
rect 35678 22480 35683 22536
rect 34145 22478 35683 22480
rect 34145 22475 34211 22478
rect 35617 22475 35683 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 59200 22312 60000 22432
rect 34930 22271 35246 22272
rect 0 22130 800 22160
rect 1761 22130 1827 22133
rect 0 22128 1827 22130
rect 0 22072 1766 22128
rect 1822 22072 1827 22128
rect 0 22070 1827 22072
rect 0 22040 800 22070
rect 1761 22067 1827 22070
rect 27521 22130 27587 22133
rect 27797 22130 27863 22133
rect 27521 22128 27863 22130
rect 27521 22072 27526 22128
rect 27582 22072 27802 22128
rect 27858 22072 27863 22128
rect 27521 22070 27863 22072
rect 27521 22067 27587 22070
rect 27797 22067 27863 22070
rect 40677 22130 40743 22133
rect 45369 22130 45435 22133
rect 40677 22128 45435 22130
rect 40677 22072 40682 22128
rect 40738 22072 45374 22128
rect 45430 22072 45435 22128
rect 40677 22070 45435 22072
rect 40677 22067 40743 22070
rect 45369 22067 45435 22070
rect 20110 21932 20116 21996
rect 20180 21994 20186 21996
rect 27521 21994 27587 21997
rect 20180 21992 27587 21994
rect 20180 21936 27526 21992
rect 27582 21936 27587 21992
rect 20180 21934 27587 21936
rect 20180 21932 20186 21934
rect 27521 21931 27587 21934
rect 30005 21994 30071 21997
rect 56317 21994 56383 21997
rect 30005 21992 56383 21994
rect 30005 21936 30010 21992
rect 30066 21936 56322 21992
rect 56378 21936 56383 21992
rect 30005 21934 56383 21936
rect 30005 21931 30071 21934
rect 56317 21931 56383 21934
rect 43989 21858 44055 21861
rect 45369 21858 45435 21861
rect 43989 21856 45435 21858
rect 43989 21800 43994 21856
rect 44050 21800 45374 21856
rect 45430 21800 45435 21856
rect 43989 21798 45435 21800
rect 43989 21795 44055 21798
rect 45369 21795 45435 21798
rect 58157 21858 58223 21861
rect 59200 21858 60000 21888
rect 58157 21856 60000 21858
rect 58157 21800 58162 21856
rect 58218 21800 60000 21856
rect 58157 21798 60000 21800
rect 58157 21795 58223 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 59200 21768 60000 21798
rect 50290 21727 50606 21728
rect 40309 21722 40375 21725
rect 47853 21722 47919 21725
rect 40309 21720 47919 21722
rect 40309 21664 40314 21720
rect 40370 21664 47858 21720
rect 47914 21664 47919 21720
rect 40309 21662 47919 21664
rect 40309 21659 40375 21662
rect 47853 21659 47919 21662
rect 40585 21586 40651 21589
rect 43897 21586 43963 21589
rect 40585 21584 43963 21586
rect 40585 21528 40590 21584
rect 40646 21528 43902 21584
rect 43958 21528 43963 21584
rect 40585 21526 43963 21528
rect 40585 21523 40651 21526
rect 43897 21523 43963 21526
rect 0 21450 800 21480
rect 1853 21450 1919 21453
rect 0 21448 1919 21450
rect 0 21392 1858 21448
rect 1914 21392 1919 21448
rect 0 21390 1919 21392
rect 0 21360 800 21390
rect 1853 21387 1919 21390
rect 57145 21314 57211 21317
rect 59200 21314 60000 21344
rect 57145 21312 60000 21314
rect 57145 21256 57150 21312
rect 57206 21256 60000 21312
rect 57145 21254 60000 21256
rect 57145 21251 57211 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 59200 21224 60000 21254
rect 34930 21183 35246 21184
rect 27797 20906 27863 20909
rect 28809 20908 28875 20909
rect 28758 20906 28764 20908
rect 27797 20904 28764 20906
rect 28828 20904 28875 20908
rect 27797 20848 27802 20904
rect 27858 20848 28764 20904
rect 28870 20848 28875 20904
rect 27797 20846 28764 20848
rect 27797 20843 27863 20846
rect 28758 20844 28764 20846
rect 28828 20844 28875 20848
rect 28809 20843 28875 20844
rect 0 20770 800 20800
rect 1853 20770 1919 20773
rect 0 20768 1919 20770
rect 0 20712 1858 20768
rect 1914 20712 1919 20768
rect 0 20710 1919 20712
rect 0 20680 800 20710
rect 1853 20707 1919 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 59200 20680 60000 20800
rect 50290 20639 50606 20640
rect 32029 20634 32095 20637
rect 39941 20634 40007 20637
rect 32029 20632 40007 20634
rect 32029 20576 32034 20632
rect 32090 20576 39946 20632
rect 40002 20576 40007 20632
rect 32029 20574 40007 20576
rect 32029 20571 32095 20574
rect 39941 20571 40007 20574
rect 58157 20226 58223 20229
rect 59200 20226 60000 20256
rect 58157 20224 60000 20226
rect 58157 20168 58162 20224
rect 58218 20168 60000 20224
rect 58157 20166 60000 20168
rect 58157 20163 58223 20166
rect 4210 20160 4526 20161
rect 0 20090 800 20120
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 59200 20136 60000 20166
rect 34930 20095 35246 20096
rect 1761 20090 1827 20093
rect 0 20088 1827 20090
rect 0 20032 1766 20088
rect 1822 20032 1827 20088
rect 0 20030 1827 20032
rect 0 20000 800 20030
rect 1761 20027 1827 20030
rect 57053 19682 57119 19685
rect 59200 19682 60000 19712
rect 57053 19680 60000 19682
rect 57053 19624 57058 19680
rect 57114 19624 60000 19680
rect 57053 19622 60000 19624
rect 57053 19619 57119 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 59200 19592 60000 19622
rect 50290 19551 50606 19552
rect 28533 19546 28599 19549
rect 29177 19546 29243 19549
rect 28533 19544 29243 19546
rect 28533 19488 28538 19544
rect 28594 19488 29182 19544
rect 29238 19488 29243 19544
rect 28533 19486 29243 19488
rect 28533 19483 28599 19486
rect 29177 19483 29243 19486
rect 29453 19546 29519 19549
rect 32581 19546 32647 19549
rect 29453 19544 32647 19546
rect 29453 19488 29458 19544
rect 29514 19488 32586 19544
rect 32642 19488 32647 19544
rect 29453 19486 32647 19488
rect 29453 19483 29519 19486
rect 32581 19483 32647 19486
rect 0 19410 800 19440
rect 1853 19410 1919 19413
rect 0 19408 1919 19410
rect 0 19352 1858 19408
rect 1914 19352 1919 19408
rect 0 19350 1919 19352
rect 0 19320 800 19350
rect 1853 19347 1919 19350
rect 27797 19410 27863 19413
rect 28533 19412 28599 19413
rect 28533 19410 28580 19412
rect 27797 19408 28580 19410
rect 27797 19352 27802 19408
rect 27858 19352 28538 19408
rect 27797 19350 28580 19352
rect 27797 19347 27863 19350
rect 28533 19348 28580 19350
rect 28644 19348 28650 19412
rect 29085 19410 29151 19413
rect 49693 19410 49759 19413
rect 29085 19408 49759 19410
rect 29085 19352 29090 19408
rect 29146 19352 49698 19408
rect 49754 19352 49759 19408
rect 29085 19350 49759 19352
rect 28533 19347 28599 19348
rect 29085 19347 29151 19350
rect 49693 19347 49759 19350
rect 27613 19274 27679 19277
rect 31293 19274 31359 19277
rect 27613 19272 31359 19274
rect 27613 19216 27618 19272
rect 27674 19216 31298 19272
rect 31354 19216 31359 19272
rect 27613 19214 31359 19216
rect 27613 19211 27679 19214
rect 31293 19211 31359 19214
rect 34697 19274 34763 19277
rect 36537 19274 36603 19277
rect 34697 19272 36603 19274
rect 34697 19216 34702 19272
rect 34758 19216 36542 19272
rect 36598 19216 36603 19272
rect 34697 19214 36603 19216
rect 34697 19211 34763 19214
rect 36537 19211 36603 19214
rect 28257 19138 28323 19141
rect 30557 19138 30623 19141
rect 28257 19136 30623 19138
rect 28257 19080 28262 19136
rect 28318 19080 30562 19136
rect 30618 19080 30623 19136
rect 28257 19078 30623 19080
rect 28257 19075 28323 19078
rect 30557 19075 30623 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 59200 19048 60000 19168
rect 34930 19007 35246 19008
rect 30741 19002 30807 19005
rect 32029 19002 32095 19005
rect 30741 19000 32095 19002
rect 30741 18944 30746 19000
rect 30802 18944 32034 19000
rect 32090 18944 32095 19000
rect 30741 18942 32095 18944
rect 30741 18939 30807 18942
rect 32029 18939 32095 18942
rect 25865 18866 25931 18869
rect 28073 18866 28139 18869
rect 57237 18866 57303 18869
rect 25865 18864 57303 18866
rect 25865 18808 25870 18864
rect 25926 18808 28078 18864
rect 28134 18808 57242 18864
rect 57298 18808 57303 18864
rect 25865 18806 57303 18808
rect 25865 18803 25931 18806
rect 28073 18803 28139 18806
rect 57237 18803 57303 18806
rect 0 18730 800 18760
rect 1853 18730 1919 18733
rect 0 18728 1919 18730
rect 0 18672 1858 18728
rect 1914 18672 1919 18728
rect 0 18670 1919 18672
rect 0 18640 800 18670
rect 1853 18667 1919 18670
rect 31293 18730 31359 18733
rect 36997 18730 37063 18733
rect 31293 18728 37063 18730
rect 31293 18672 31298 18728
rect 31354 18672 37002 18728
rect 37058 18672 37063 18728
rect 31293 18670 37063 18672
rect 31293 18667 31359 18670
rect 36997 18667 37063 18670
rect 28441 18594 28507 18597
rect 31569 18594 31635 18597
rect 36353 18594 36419 18597
rect 28441 18592 31635 18594
rect 28441 18536 28446 18592
rect 28502 18536 31574 18592
rect 31630 18536 31635 18592
rect 28441 18534 31635 18536
rect 28441 18531 28507 18534
rect 31569 18531 31635 18534
rect 31710 18592 36419 18594
rect 31710 18536 36358 18592
rect 36414 18536 36419 18592
rect 31710 18534 36419 18536
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 24577 18458 24643 18461
rect 28809 18458 28875 18461
rect 24577 18456 28875 18458
rect 24577 18400 24582 18456
rect 24638 18400 28814 18456
rect 28870 18400 28875 18456
rect 24577 18398 28875 18400
rect 24577 18395 24643 18398
rect 28809 18395 28875 18398
rect 30741 18458 30807 18461
rect 31710 18458 31770 18534
rect 36353 18531 36419 18534
rect 58157 18594 58223 18597
rect 59200 18594 60000 18624
rect 58157 18592 60000 18594
rect 58157 18536 58162 18592
rect 58218 18536 60000 18592
rect 58157 18534 60000 18536
rect 58157 18531 58223 18534
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 59200 18504 60000 18534
rect 50290 18463 50606 18464
rect 30741 18456 31770 18458
rect 30741 18400 30746 18456
rect 30802 18400 31770 18456
rect 30741 18398 31770 18400
rect 33133 18458 33199 18461
rect 34881 18458 34947 18461
rect 33133 18456 34947 18458
rect 33133 18400 33138 18456
rect 33194 18400 34886 18456
rect 34942 18400 34947 18456
rect 33133 18398 34947 18400
rect 30741 18395 30807 18398
rect 33133 18395 33199 18398
rect 34881 18395 34947 18398
rect 26233 18322 26299 18325
rect 26601 18322 26667 18325
rect 34329 18322 34395 18325
rect 26233 18320 34395 18322
rect 26233 18264 26238 18320
rect 26294 18264 26606 18320
rect 26662 18264 34334 18320
rect 34390 18264 34395 18320
rect 26233 18262 34395 18264
rect 26233 18259 26299 18262
rect 26601 18259 26667 18262
rect 34329 18259 34395 18262
rect 26325 18186 26391 18189
rect 28993 18186 29059 18189
rect 26325 18184 29059 18186
rect 26325 18128 26330 18184
rect 26386 18128 28998 18184
rect 29054 18128 29059 18184
rect 26325 18126 29059 18128
rect 26325 18123 26391 18126
rect 28993 18123 29059 18126
rect 30833 18186 30899 18189
rect 38101 18186 38167 18189
rect 30833 18184 38167 18186
rect 30833 18128 30838 18184
rect 30894 18128 38106 18184
rect 38162 18128 38167 18184
rect 30833 18126 38167 18128
rect 30833 18123 30899 18126
rect 38101 18123 38167 18126
rect 0 18050 800 18080
rect 1761 18050 1827 18053
rect 0 18048 1827 18050
rect 0 17992 1766 18048
rect 1822 17992 1827 18048
rect 0 17990 1827 17992
rect 0 17960 800 17990
rect 1761 17987 1827 17990
rect 27153 18050 27219 18053
rect 28533 18050 28599 18053
rect 27153 18048 28599 18050
rect 27153 17992 27158 18048
rect 27214 17992 28538 18048
rect 28594 17992 28599 18048
rect 27153 17990 28599 17992
rect 27153 17987 27219 17990
rect 28533 17987 28599 17990
rect 30465 18050 30531 18053
rect 32673 18050 32739 18053
rect 30465 18048 32739 18050
rect 30465 17992 30470 18048
rect 30526 17992 32678 18048
rect 32734 17992 32739 18048
rect 30465 17990 32739 17992
rect 30465 17987 30531 17990
rect 32673 17987 32739 17990
rect 32857 18050 32923 18053
rect 32990 18050 32996 18052
rect 32857 18048 32996 18050
rect 32857 17992 32862 18048
rect 32918 17992 32996 18048
rect 32857 17990 32996 17992
rect 32857 17987 32923 17990
rect 32990 17988 32996 17990
rect 33060 17988 33066 18052
rect 57053 18050 57119 18053
rect 59200 18050 60000 18080
rect 57053 18048 60000 18050
rect 57053 17992 57058 18048
rect 57114 17992 60000 18048
rect 57053 17990 60000 17992
rect 57053 17987 57119 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 59200 17960 60000 17990
rect 34930 17919 35246 17920
rect 30557 17914 30623 17917
rect 31017 17914 31083 17917
rect 30557 17912 31083 17914
rect 30557 17856 30562 17912
rect 30618 17856 31022 17912
rect 31078 17856 31083 17912
rect 30557 17854 31083 17856
rect 30557 17851 30623 17854
rect 31017 17851 31083 17854
rect 32029 17916 32095 17917
rect 33133 17916 33199 17917
rect 32029 17912 32076 17916
rect 32140 17914 32146 17916
rect 32029 17856 32034 17912
rect 32029 17852 32076 17856
rect 32140 17854 32186 17914
rect 33133 17912 33180 17916
rect 33244 17914 33250 17916
rect 33133 17856 33138 17912
rect 32140 17852 32146 17854
rect 33133 17852 33180 17856
rect 33244 17854 33290 17914
rect 33244 17852 33250 17854
rect 32029 17851 32095 17852
rect 33133 17851 33199 17852
rect 29729 17778 29795 17781
rect 38193 17778 38259 17781
rect 29729 17776 38259 17778
rect 29729 17720 29734 17776
rect 29790 17720 38198 17776
rect 38254 17720 38259 17776
rect 29729 17718 38259 17720
rect 29729 17715 29795 17718
rect 38193 17715 38259 17718
rect 22829 17642 22895 17645
rect 29453 17642 29519 17645
rect 22829 17640 29519 17642
rect 22829 17584 22834 17640
rect 22890 17584 29458 17640
rect 29514 17584 29519 17640
rect 22829 17582 29519 17584
rect 22829 17579 22895 17582
rect 29453 17579 29519 17582
rect 30005 17642 30071 17645
rect 32121 17642 32187 17645
rect 30005 17640 32187 17642
rect 30005 17584 30010 17640
rect 30066 17584 32126 17640
rect 32182 17584 32187 17640
rect 30005 17582 32187 17584
rect 30005 17579 30071 17582
rect 32121 17579 32187 17582
rect 28349 17506 28415 17509
rect 33225 17506 33291 17509
rect 28349 17504 33291 17506
rect 28349 17448 28354 17504
rect 28410 17448 33230 17504
rect 33286 17448 33291 17504
rect 28349 17446 33291 17448
rect 28349 17443 28415 17446
rect 33225 17443 33291 17446
rect 19570 17440 19886 17441
rect 0 17370 800 17400
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 59200 17416 60000 17536
rect 50290 17375 50606 17376
rect 1853 17370 1919 17373
rect 0 17368 1919 17370
rect 0 17312 1858 17368
rect 1914 17312 1919 17368
rect 0 17310 1919 17312
rect 0 17280 800 17310
rect 1853 17307 1919 17310
rect 21081 17370 21147 17373
rect 22645 17370 22711 17373
rect 21081 17368 22711 17370
rect 21081 17312 21086 17368
rect 21142 17312 22650 17368
rect 22706 17312 22711 17368
rect 21081 17310 22711 17312
rect 21081 17307 21147 17310
rect 22645 17307 22711 17310
rect 30097 17370 30163 17373
rect 30741 17370 30807 17373
rect 30097 17368 30807 17370
rect 30097 17312 30102 17368
rect 30158 17312 30746 17368
rect 30802 17312 30807 17368
rect 30097 17310 30807 17312
rect 30097 17307 30163 17310
rect 30741 17307 30807 17310
rect 13537 17234 13603 17237
rect 33593 17234 33659 17237
rect 13537 17232 33659 17234
rect 13537 17176 13542 17232
rect 13598 17176 33598 17232
rect 33654 17176 33659 17232
rect 13537 17174 33659 17176
rect 13537 17171 13603 17174
rect 33593 17171 33659 17174
rect 22645 17098 22711 17101
rect 25497 17098 25563 17101
rect 22645 17096 25563 17098
rect 22645 17040 22650 17096
rect 22706 17040 25502 17096
rect 25558 17040 25563 17096
rect 22645 17038 25563 17040
rect 22645 17035 22711 17038
rect 25497 17035 25563 17038
rect 29177 17098 29243 17101
rect 31937 17098 32003 17101
rect 29177 17096 32003 17098
rect 29177 17040 29182 17096
rect 29238 17040 31942 17096
rect 31998 17040 32003 17096
rect 29177 17038 32003 17040
rect 29177 17035 29243 17038
rect 31937 17035 32003 17038
rect 30281 16962 30347 16965
rect 34513 16962 34579 16965
rect 30281 16960 34579 16962
rect 30281 16904 30286 16960
rect 30342 16904 34518 16960
rect 34574 16904 34579 16960
rect 30281 16902 34579 16904
rect 30281 16899 30347 16902
rect 34513 16899 34579 16902
rect 57329 16962 57395 16965
rect 59200 16962 60000 16992
rect 57329 16960 60000 16962
rect 57329 16904 57334 16960
rect 57390 16904 60000 16960
rect 57329 16902 60000 16904
rect 57329 16899 57395 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 59200 16872 60000 16902
rect 34930 16831 35246 16832
rect 19977 16826 20043 16829
rect 32489 16826 32555 16829
rect 19977 16824 32555 16826
rect 19977 16768 19982 16824
rect 20038 16768 32494 16824
rect 32550 16768 32555 16824
rect 19977 16766 32555 16768
rect 19977 16763 20043 16766
rect 32489 16763 32555 16766
rect 0 16690 800 16720
rect 1761 16690 1827 16693
rect 0 16688 1827 16690
rect 0 16632 1766 16688
rect 1822 16632 1827 16688
rect 0 16630 1827 16632
rect 0 16600 800 16630
rect 1761 16627 1827 16630
rect 29361 16690 29427 16693
rect 30925 16690 30991 16693
rect 29361 16688 30991 16690
rect 29361 16632 29366 16688
rect 29422 16632 30930 16688
rect 30986 16632 30991 16688
rect 29361 16630 30991 16632
rect 29361 16627 29427 16630
rect 30925 16627 30991 16630
rect 31569 16690 31635 16693
rect 31886 16690 31892 16692
rect 31569 16688 31892 16690
rect 31569 16632 31574 16688
rect 31630 16632 31892 16688
rect 31569 16630 31892 16632
rect 31569 16627 31635 16630
rect 31886 16628 31892 16630
rect 31956 16628 31962 16692
rect 38653 16690 38719 16693
rect 43897 16690 43963 16693
rect 38653 16688 43963 16690
rect 38653 16632 38658 16688
rect 38714 16632 43902 16688
rect 43958 16632 43963 16688
rect 38653 16630 43963 16632
rect 38653 16627 38719 16630
rect 43897 16627 43963 16630
rect 17309 16554 17375 16557
rect 18137 16554 18203 16557
rect 17309 16552 18203 16554
rect 17309 16496 17314 16552
rect 17370 16496 18142 16552
rect 18198 16496 18203 16552
rect 17309 16494 18203 16496
rect 17309 16491 17375 16494
rect 18137 16491 18203 16494
rect 31109 16554 31175 16557
rect 36353 16554 36419 16557
rect 31109 16552 36419 16554
rect 31109 16496 31114 16552
rect 31170 16496 36358 16552
rect 36414 16496 36419 16552
rect 31109 16494 36419 16496
rect 31109 16491 31175 16494
rect 36353 16491 36419 16494
rect 20529 16418 20595 16421
rect 25405 16418 25471 16421
rect 28257 16418 28323 16421
rect 20529 16416 28323 16418
rect 20529 16360 20534 16416
rect 20590 16360 25410 16416
rect 25466 16360 28262 16416
rect 28318 16360 28323 16416
rect 20529 16358 28323 16360
rect 20529 16355 20595 16358
rect 25405 16355 25471 16358
rect 28257 16355 28323 16358
rect 57973 16418 58039 16421
rect 59200 16418 60000 16448
rect 57973 16416 60000 16418
rect 57973 16360 57978 16416
rect 58034 16360 60000 16416
rect 57973 16358 60000 16360
rect 57973 16355 58039 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 59200 16328 60000 16358
rect 50290 16287 50606 16288
rect 18229 16148 18295 16149
rect 18229 16146 18276 16148
rect 18184 16144 18276 16146
rect 18184 16088 18234 16144
rect 18184 16086 18276 16088
rect 18229 16084 18276 16086
rect 18340 16084 18346 16148
rect 18229 16083 18295 16084
rect 0 16010 800 16040
rect 1761 16010 1827 16013
rect 0 16008 1827 16010
rect 0 15952 1766 16008
rect 1822 15952 1827 16008
rect 0 15950 1827 15952
rect 0 15920 800 15950
rect 1761 15947 1827 15950
rect 21449 16010 21515 16013
rect 23197 16010 23263 16013
rect 21449 16008 23263 16010
rect 21449 15952 21454 16008
rect 21510 15952 23202 16008
rect 23258 15952 23263 16008
rect 21449 15950 23263 15952
rect 21449 15947 21515 15950
rect 23197 15947 23263 15950
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 59200 15784 60000 15904
rect 34930 15743 35246 15744
rect 34329 15602 34395 15605
rect 34646 15602 34652 15604
rect 34329 15600 34652 15602
rect 34329 15544 34334 15600
rect 34390 15544 34652 15600
rect 34329 15542 34652 15544
rect 34329 15539 34395 15542
rect 34646 15540 34652 15542
rect 34716 15540 34722 15604
rect 19517 15466 19583 15469
rect 21817 15466 21883 15469
rect 23565 15466 23631 15469
rect 19517 15464 23631 15466
rect 19517 15408 19522 15464
rect 19578 15408 21822 15464
rect 21878 15408 23570 15464
rect 23626 15408 23631 15464
rect 19517 15406 23631 15408
rect 19517 15403 19583 15406
rect 21817 15403 21883 15406
rect 23565 15403 23631 15406
rect 0 15330 800 15360
rect 1853 15330 1919 15333
rect 0 15328 1919 15330
rect 0 15272 1858 15328
rect 1914 15272 1919 15328
rect 0 15270 1919 15272
rect 0 15240 800 15270
rect 1853 15267 1919 15270
rect 57237 15330 57303 15333
rect 59200 15330 60000 15360
rect 57237 15328 60000 15330
rect 57237 15272 57242 15328
rect 57298 15272 60000 15328
rect 57237 15270 60000 15272
rect 57237 15267 57303 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 59200 15240 60000 15270
rect 50290 15199 50606 15200
rect 19425 15060 19491 15061
rect 19374 15058 19380 15060
rect 19334 14998 19380 15058
rect 19444 15056 19491 15060
rect 19486 15000 19491 15056
rect 19374 14996 19380 14998
rect 19444 14996 19491 15000
rect 19425 14995 19491 14996
rect 33869 14922 33935 14925
rect 45001 14922 45067 14925
rect 33869 14920 45067 14922
rect 33869 14864 33874 14920
rect 33930 14864 45006 14920
rect 45062 14864 45067 14920
rect 33869 14862 45067 14864
rect 33869 14859 33935 14862
rect 45001 14859 45067 14862
rect 17125 14786 17191 14789
rect 17401 14786 17467 14789
rect 26785 14786 26851 14789
rect 17125 14784 26851 14786
rect 17125 14728 17130 14784
rect 17186 14728 17406 14784
rect 17462 14728 26790 14784
rect 26846 14728 26851 14784
rect 17125 14726 26851 14728
rect 17125 14723 17191 14726
rect 17401 14723 17467 14726
rect 26785 14723 26851 14726
rect 57973 14786 58039 14789
rect 59200 14786 60000 14816
rect 57973 14784 60000 14786
rect 57973 14728 57978 14784
rect 58034 14728 60000 14784
rect 57973 14726 60000 14728
rect 57973 14723 58039 14726
rect 4210 14720 4526 14721
rect 0 14650 800 14680
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 59200 14696 60000 14726
rect 34930 14655 35246 14656
rect 1761 14650 1827 14653
rect 0 14648 1827 14650
rect 0 14592 1766 14648
rect 1822 14592 1827 14648
rect 0 14590 1827 14592
rect 0 14560 800 14590
rect 1761 14587 1827 14590
rect 21357 14514 21423 14517
rect 25405 14514 25471 14517
rect 58065 14514 58131 14517
rect 21357 14512 25471 14514
rect 21357 14456 21362 14512
rect 21418 14456 25410 14512
rect 25466 14456 25471 14512
rect 21357 14454 25471 14456
rect 21357 14451 21423 14454
rect 25405 14451 25471 14454
rect 31710 14512 58131 14514
rect 31710 14456 58070 14512
rect 58126 14456 58131 14512
rect 31710 14454 58131 14456
rect 25313 14378 25379 14381
rect 31477 14378 31543 14381
rect 31710 14378 31770 14454
rect 58065 14451 58131 14454
rect 25313 14376 31770 14378
rect 25313 14320 25318 14376
rect 25374 14320 31482 14376
rect 31538 14320 31770 14376
rect 25313 14318 31770 14320
rect 25313 14315 25379 14318
rect 31477 14315 31543 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 59200 14152 60000 14272
rect 50290 14111 50606 14112
rect 0 13970 800 14000
rect 1853 13970 1919 13973
rect 0 13968 1919 13970
rect 0 13912 1858 13968
rect 1914 13912 1919 13968
rect 0 13910 1919 13912
rect 0 13880 800 13910
rect 1853 13907 1919 13910
rect 30741 13970 30807 13973
rect 32305 13970 32371 13973
rect 30741 13968 32371 13970
rect 30741 13912 30746 13968
rect 30802 13912 32310 13968
rect 32366 13912 32371 13968
rect 30741 13910 32371 13912
rect 30741 13907 30807 13910
rect 32305 13907 32371 13910
rect 38142 13636 38148 13700
rect 38212 13698 38218 13700
rect 41137 13698 41203 13701
rect 38212 13696 41203 13698
rect 38212 13640 41142 13696
rect 41198 13640 41203 13696
rect 38212 13638 41203 13640
rect 38212 13636 38218 13638
rect 41137 13635 41203 13638
rect 57329 13698 57395 13701
rect 59200 13698 60000 13728
rect 57329 13696 60000 13698
rect 57329 13640 57334 13696
rect 57390 13640 60000 13696
rect 57329 13638 60000 13640
rect 57329 13635 57395 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 59200 13608 60000 13638
rect 34930 13567 35246 13568
rect 16757 13426 16823 13429
rect 23606 13426 23612 13428
rect 16757 13424 23612 13426
rect 16757 13368 16762 13424
rect 16818 13368 23612 13424
rect 16757 13366 23612 13368
rect 16757 13363 16823 13366
rect 23606 13364 23612 13366
rect 23676 13364 23682 13428
rect 0 13290 800 13320
rect 1853 13290 1919 13293
rect 0 13288 1919 13290
rect 0 13232 1858 13288
rect 1914 13232 1919 13288
rect 0 13230 1919 13232
rect 0 13200 800 13230
rect 1853 13227 1919 13230
rect 57973 13154 58039 13157
rect 59200 13154 60000 13184
rect 57973 13152 60000 13154
rect 57973 13096 57978 13152
rect 58034 13096 60000 13152
rect 57973 13094 60000 13096
rect 57973 13091 58039 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 59200 13064 60000 13094
rect 50290 13023 50606 13024
rect 21357 13018 21423 13021
rect 31569 13018 31635 13021
rect 21357 13016 31635 13018
rect 21357 12960 21362 13016
rect 21418 12960 31574 13016
rect 31630 12960 31635 13016
rect 21357 12958 31635 12960
rect 21357 12955 21423 12958
rect 31569 12955 31635 12958
rect 0 12610 800 12640
rect 1761 12610 1827 12613
rect 0 12608 1827 12610
rect 0 12552 1766 12608
rect 1822 12552 1827 12608
rect 0 12550 1827 12552
rect 0 12520 800 12550
rect 1761 12547 1827 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 59200 12520 60000 12640
rect 34930 12479 35246 12480
rect 19885 12338 19951 12341
rect 20989 12338 21055 12341
rect 19885 12336 21055 12338
rect 19885 12280 19890 12336
rect 19946 12280 20994 12336
rect 21050 12280 21055 12336
rect 19885 12278 21055 12280
rect 19885 12275 19951 12278
rect 20989 12275 21055 12278
rect 57237 12066 57303 12069
rect 59200 12066 60000 12096
rect 57237 12064 60000 12066
rect 57237 12008 57242 12064
rect 57298 12008 60000 12064
rect 57237 12006 60000 12008
rect 57237 12003 57303 12006
rect 19570 12000 19886 12001
rect 0 11930 800 11960
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 59200 11976 60000 12006
rect 50290 11935 50606 11936
rect 1853 11930 1919 11933
rect 0 11928 1919 11930
rect 0 11872 1858 11928
rect 1914 11872 1919 11928
rect 0 11870 1919 11872
rect 0 11840 800 11870
rect 1853 11867 1919 11870
rect 15009 11794 15075 11797
rect 33685 11794 33751 11797
rect 15009 11792 33751 11794
rect 15009 11736 15014 11792
rect 15070 11736 33690 11792
rect 33746 11736 33751 11792
rect 15009 11734 33751 11736
rect 15009 11731 15075 11734
rect 33685 11731 33751 11734
rect 33961 11794 34027 11797
rect 34697 11794 34763 11797
rect 33961 11792 34763 11794
rect 33961 11736 33966 11792
rect 34022 11736 34702 11792
rect 34758 11736 34763 11792
rect 33961 11734 34763 11736
rect 33961 11731 34027 11734
rect 34697 11731 34763 11734
rect 19374 11596 19380 11660
rect 19444 11658 19450 11660
rect 19793 11658 19859 11661
rect 19444 11656 19859 11658
rect 19444 11600 19798 11656
rect 19854 11600 19859 11656
rect 19444 11598 19859 11600
rect 19444 11596 19450 11598
rect 19793 11595 19859 11598
rect 30966 11596 30972 11660
rect 31036 11658 31042 11660
rect 33409 11658 33475 11661
rect 35341 11658 35407 11661
rect 31036 11656 33475 11658
rect 31036 11600 33414 11656
rect 33470 11600 33475 11656
rect 31036 11598 33475 11600
rect 31036 11596 31042 11598
rect 33409 11595 33475 11598
rect 33550 11656 35407 11658
rect 33550 11600 35346 11656
rect 35402 11600 35407 11656
rect 33550 11598 35407 11600
rect 24485 11522 24551 11525
rect 33550 11522 33610 11598
rect 35341 11595 35407 11598
rect 24485 11520 33610 11522
rect 24485 11464 24490 11520
rect 24546 11464 33610 11520
rect 24485 11462 33610 11464
rect 57145 11522 57211 11525
rect 59200 11522 60000 11552
rect 57145 11520 60000 11522
rect 57145 11464 57150 11520
rect 57206 11464 60000 11520
rect 57145 11462 60000 11464
rect 24485 11459 24551 11462
rect 57145 11459 57211 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 59200 11432 60000 11462
rect 34930 11391 35246 11392
rect 0 11250 800 11280
rect 1761 11250 1827 11253
rect 0 11248 1827 11250
rect 0 11192 1766 11248
rect 1822 11192 1827 11248
rect 0 11190 1827 11192
rect 0 11160 800 11190
rect 1761 11187 1827 11190
rect 19333 11250 19399 11253
rect 20345 11250 20411 11253
rect 19333 11248 20411 11250
rect 19333 11192 19338 11248
rect 19394 11192 20350 11248
rect 20406 11192 20411 11248
rect 19333 11190 20411 11192
rect 19333 11187 19399 11190
rect 20345 11187 20411 11190
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 59200 10888 60000 11008
rect 50290 10847 50606 10848
rect 27061 10706 27127 10709
rect 29269 10706 29335 10709
rect 31109 10706 31175 10709
rect 27061 10704 31175 10706
rect 27061 10648 27066 10704
rect 27122 10648 29274 10704
rect 29330 10648 31114 10704
rect 31170 10648 31175 10704
rect 27061 10646 31175 10648
rect 27061 10643 27127 10646
rect 29269 10643 29335 10646
rect 31109 10643 31175 10646
rect 0 10570 800 10600
rect 1761 10570 1827 10573
rect 0 10568 1827 10570
rect 0 10512 1766 10568
rect 1822 10512 1827 10568
rect 0 10510 1827 10512
rect 0 10480 800 10510
rect 1761 10507 1827 10510
rect 21541 10434 21607 10437
rect 26785 10434 26851 10437
rect 21541 10432 26851 10434
rect 21541 10376 21546 10432
rect 21602 10376 26790 10432
rect 26846 10376 26851 10432
rect 21541 10374 26851 10376
rect 21541 10371 21607 10374
rect 26785 10371 26851 10374
rect 26969 10434 27035 10437
rect 30557 10434 30623 10437
rect 31477 10434 31543 10437
rect 26969 10432 31543 10434
rect 26969 10376 26974 10432
rect 27030 10376 30562 10432
rect 30618 10376 31482 10432
rect 31538 10376 31543 10432
rect 26969 10374 31543 10376
rect 26969 10371 27035 10374
rect 30557 10371 30623 10374
rect 31477 10371 31543 10374
rect 58157 10434 58223 10437
rect 59200 10434 60000 10464
rect 58157 10432 60000 10434
rect 58157 10376 58162 10432
rect 58218 10376 60000 10432
rect 58157 10374 60000 10376
rect 58157 10371 58223 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 59200 10344 60000 10374
rect 34930 10303 35246 10304
rect 20069 10298 20135 10301
rect 22001 10298 22067 10301
rect 20069 10296 22067 10298
rect 20069 10240 20074 10296
rect 20130 10240 22006 10296
rect 22062 10240 22067 10296
rect 20069 10238 22067 10240
rect 20069 10235 20135 10238
rect 22001 10235 22067 10238
rect 19149 10162 19215 10165
rect 22093 10162 22159 10165
rect 19149 10160 22159 10162
rect 19149 10104 19154 10160
rect 19210 10104 22098 10160
rect 22154 10104 22159 10160
rect 19149 10102 22159 10104
rect 19149 10099 19215 10102
rect 22093 10099 22159 10102
rect 23749 10026 23815 10029
rect 25497 10026 25563 10029
rect 23749 10024 25563 10026
rect 23749 9968 23754 10024
rect 23810 9968 25502 10024
rect 25558 9968 25563 10024
rect 23749 9966 25563 9968
rect 23749 9963 23815 9966
rect 25497 9963 25563 9966
rect 0 9890 800 9920
rect 1853 9890 1919 9893
rect 0 9888 1919 9890
rect 0 9832 1858 9888
rect 1914 9832 1919 9888
rect 0 9830 1919 9832
rect 0 9800 800 9830
rect 1853 9827 1919 9830
rect 57053 9890 57119 9893
rect 59200 9890 60000 9920
rect 57053 9888 60000 9890
rect 57053 9832 57058 9888
rect 57114 9832 60000 9888
rect 57053 9830 60000 9832
rect 57053 9827 57119 9830
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 59200 9800 60000 9830
rect 50290 9759 50606 9760
rect 23565 9754 23631 9757
rect 29177 9754 29243 9757
rect 23565 9752 29243 9754
rect 23565 9696 23570 9752
rect 23626 9696 29182 9752
rect 29238 9696 29243 9752
rect 23565 9694 29243 9696
rect 23565 9691 23631 9694
rect 29177 9691 29243 9694
rect 30005 9754 30071 9757
rect 33685 9754 33751 9757
rect 30005 9752 33751 9754
rect 30005 9696 30010 9752
rect 30066 9696 33690 9752
rect 33746 9696 33751 9752
rect 30005 9694 33751 9696
rect 30005 9691 30071 9694
rect 33685 9691 33751 9694
rect 30373 9618 30439 9621
rect 31518 9618 31524 9620
rect 30373 9616 31524 9618
rect 30373 9560 30378 9616
rect 30434 9560 31524 9616
rect 30373 9558 31524 9560
rect 30373 9555 30439 9558
rect 31518 9556 31524 9558
rect 31588 9556 31594 9620
rect 35065 9618 35131 9621
rect 35566 9618 35572 9620
rect 35065 9616 35572 9618
rect 35065 9560 35070 9616
rect 35126 9560 35572 9616
rect 35065 9558 35572 9560
rect 35065 9555 35131 9558
rect 35566 9556 35572 9558
rect 35636 9556 35642 9620
rect 27429 9482 27495 9485
rect 28165 9482 28231 9485
rect 27429 9480 28231 9482
rect 27429 9424 27434 9480
rect 27490 9424 28170 9480
rect 28226 9424 28231 9480
rect 27429 9422 28231 9424
rect 27429 9419 27495 9422
rect 28165 9419 28231 9422
rect 30281 9482 30347 9485
rect 31201 9482 31267 9485
rect 30281 9480 31267 9482
rect 30281 9424 30286 9480
rect 30342 9424 31206 9480
rect 31262 9424 31267 9480
rect 30281 9422 31267 9424
rect 30281 9419 30347 9422
rect 31201 9419 31267 9422
rect 4210 9280 4526 9281
rect 0 9210 800 9240
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 59200 9256 60000 9376
rect 34930 9215 35246 9216
rect 1761 9210 1827 9213
rect 0 9208 1827 9210
rect 0 9152 1766 9208
rect 1822 9152 1827 9208
rect 0 9150 1827 9152
rect 0 9120 800 9150
rect 1761 9147 1827 9150
rect 13905 9074 13971 9077
rect 24526 9074 24532 9076
rect 13905 9072 24532 9074
rect 13905 9016 13910 9072
rect 13966 9016 24532 9072
rect 13905 9014 24532 9016
rect 13905 9011 13971 9014
rect 24526 9012 24532 9014
rect 24596 9012 24602 9076
rect 14089 8938 14155 8941
rect 25446 8938 25452 8940
rect 14089 8936 25452 8938
rect 14089 8880 14094 8936
rect 14150 8880 25452 8936
rect 14089 8878 25452 8880
rect 14089 8875 14155 8878
rect 25446 8876 25452 8878
rect 25516 8876 25522 8940
rect 32121 8938 32187 8941
rect 32857 8938 32923 8941
rect 32121 8936 32923 8938
rect 32121 8880 32126 8936
rect 32182 8880 32862 8936
rect 32918 8880 32923 8936
rect 32121 8878 32923 8880
rect 32121 8875 32187 8878
rect 32857 8875 32923 8878
rect 57329 8802 57395 8805
rect 59200 8802 60000 8832
rect 57329 8800 60000 8802
rect 57329 8744 57334 8800
rect 57390 8744 60000 8800
rect 57329 8742 60000 8744
rect 57329 8739 57395 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 59200 8712 60000 8742
rect 50290 8671 50606 8672
rect 0 8530 800 8560
rect 1853 8530 1919 8533
rect 0 8528 1919 8530
rect 0 8472 1858 8528
rect 1914 8472 1919 8528
rect 0 8470 1919 8472
rect 0 8440 800 8470
rect 1853 8467 1919 8470
rect 34881 8530 34947 8533
rect 38653 8530 38719 8533
rect 34881 8528 38719 8530
rect 34881 8472 34886 8528
rect 34942 8472 38658 8528
rect 38714 8472 38719 8528
rect 34881 8470 38719 8472
rect 34881 8467 34947 8470
rect 38653 8467 38719 8470
rect 26049 8394 26115 8397
rect 29494 8394 29500 8396
rect 26049 8392 29500 8394
rect 26049 8336 26054 8392
rect 26110 8336 29500 8392
rect 26049 8334 29500 8336
rect 26049 8331 26115 8334
rect 29494 8332 29500 8334
rect 29564 8332 29570 8396
rect 31569 8394 31635 8397
rect 37273 8394 37339 8397
rect 31569 8392 37339 8394
rect 31569 8336 31574 8392
rect 31630 8336 37278 8392
rect 37334 8336 37339 8392
rect 31569 8334 37339 8336
rect 31569 8331 31635 8334
rect 37273 8331 37339 8334
rect 19057 8258 19123 8261
rect 20713 8258 20779 8261
rect 19057 8256 20779 8258
rect 19057 8200 19062 8256
rect 19118 8200 20718 8256
rect 20774 8200 20779 8256
rect 19057 8198 20779 8200
rect 19057 8195 19123 8198
rect 20713 8195 20779 8198
rect 56225 8258 56291 8261
rect 59200 8258 60000 8288
rect 56225 8256 60000 8258
rect 56225 8200 56230 8256
rect 56286 8200 60000 8256
rect 56225 8198 60000 8200
rect 56225 8195 56291 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 59200 8168 60000 8198
rect 34930 8127 35246 8128
rect 34145 7986 34211 7989
rect 38101 7986 38167 7989
rect 34145 7984 38167 7986
rect 34145 7928 34150 7984
rect 34206 7928 38106 7984
rect 38162 7928 38167 7984
rect 34145 7926 38167 7928
rect 34145 7923 34211 7926
rect 38101 7923 38167 7926
rect 0 7850 800 7880
rect 1853 7850 1919 7853
rect 0 7848 1919 7850
rect 0 7792 1858 7848
rect 1914 7792 1919 7848
rect 0 7790 1919 7792
rect 0 7760 800 7790
rect 1853 7787 1919 7790
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 59200 7624 60000 7744
rect 50290 7583 50606 7584
rect 33777 7442 33843 7445
rect 36445 7442 36511 7445
rect 33777 7440 36511 7442
rect 33777 7384 33782 7440
rect 33838 7384 36450 7440
rect 36506 7384 36511 7440
rect 33777 7382 36511 7384
rect 33777 7379 33843 7382
rect 36445 7379 36511 7382
rect 38653 7442 38719 7445
rect 39941 7442 40007 7445
rect 38653 7440 40007 7442
rect 38653 7384 38658 7440
rect 38714 7384 39946 7440
rect 40002 7384 40007 7440
rect 38653 7382 40007 7384
rect 38653 7379 38719 7382
rect 39941 7379 40007 7382
rect 19793 7306 19859 7309
rect 27153 7306 27219 7309
rect 19793 7304 27219 7306
rect 19793 7248 19798 7304
rect 19854 7248 27158 7304
rect 27214 7248 27219 7304
rect 19793 7246 27219 7248
rect 19793 7243 19859 7246
rect 27153 7243 27219 7246
rect 0 7170 800 7200
rect 1761 7170 1827 7173
rect 0 7168 1827 7170
rect 0 7112 1766 7168
rect 1822 7112 1827 7168
rect 0 7110 1827 7112
rect 0 7080 800 7110
rect 1761 7107 1827 7110
rect 56409 7170 56475 7173
rect 59200 7170 60000 7200
rect 56409 7168 60000 7170
rect 56409 7112 56414 7168
rect 56470 7112 60000 7168
rect 56409 7110 60000 7112
rect 56409 7107 56475 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 59200 7080 60000 7110
rect 34930 7039 35246 7040
rect 22185 7034 22251 7037
rect 28625 7034 28691 7037
rect 22185 7032 28691 7034
rect 22185 6976 22190 7032
rect 22246 6976 28630 7032
rect 28686 6976 28691 7032
rect 22185 6974 28691 6976
rect 22185 6971 22251 6974
rect 28625 6971 28691 6974
rect 22093 6898 22159 6901
rect 23565 6900 23631 6901
rect 24577 6900 24643 6901
rect 22093 6896 22570 6898
rect 22093 6840 22098 6896
rect 22154 6840 22570 6896
rect 22093 6838 22570 6840
rect 22093 6835 22159 6838
rect 2037 6762 2103 6765
rect 22369 6762 22435 6765
rect 2037 6760 22435 6762
rect 2037 6704 2042 6760
rect 2098 6704 22374 6760
rect 22430 6704 22435 6760
rect 2037 6702 22435 6704
rect 22510 6762 22570 6838
rect 23565 6896 23612 6900
rect 23676 6898 23682 6900
rect 23565 6840 23570 6896
rect 23565 6836 23612 6840
rect 23676 6838 23722 6898
rect 23676 6836 23682 6838
rect 24526 6836 24532 6900
rect 24596 6898 24643 6900
rect 24596 6896 24688 6898
rect 24638 6840 24688 6896
rect 24596 6838 24688 6840
rect 24596 6836 24643 6838
rect 23565 6835 23631 6836
rect 24577 6835 24643 6836
rect 25129 6762 25195 6765
rect 22510 6760 25195 6762
rect 22510 6704 25134 6760
rect 25190 6704 25195 6760
rect 22510 6702 25195 6704
rect 2037 6699 2103 6702
rect 22369 6699 22435 6702
rect 25129 6699 25195 6702
rect 20253 6626 20319 6629
rect 22829 6626 22895 6629
rect 20253 6624 22895 6626
rect 20253 6568 20258 6624
rect 20314 6568 22834 6624
rect 22890 6568 22895 6624
rect 20253 6566 22895 6568
rect 20253 6563 20319 6566
rect 22829 6563 22895 6566
rect 57973 6626 58039 6629
rect 59200 6626 60000 6656
rect 57973 6624 60000 6626
rect 57973 6568 57978 6624
rect 58034 6568 60000 6624
rect 57973 6566 60000 6568
rect 57973 6563 58039 6566
rect 19570 6560 19886 6561
rect 0 6490 800 6520
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 59200 6536 60000 6566
rect 50290 6495 50606 6496
rect 1853 6490 1919 6493
rect 0 6488 1919 6490
rect 0 6432 1858 6488
rect 1914 6432 1919 6488
rect 0 6430 1919 6432
rect 0 6400 800 6430
rect 1853 6427 1919 6430
rect 17861 6490 17927 6493
rect 19241 6490 19307 6493
rect 17861 6488 19307 6490
rect 17861 6432 17866 6488
rect 17922 6432 19246 6488
rect 19302 6432 19307 6488
rect 17861 6430 19307 6432
rect 17861 6427 17927 6430
rect 19241 6427 19307 6430
rect 21633 6490 21699 6493
rect 24025 6490 24091 6493
rect 21633 6488 24091 6490
rect 21633 6432 21638 6488
rect 21694 6432 24030 6488
rect 24086 6432 24091 6488
rect 21633 6430 24091 6432
rect 21633 6427 21699 6430
rect 24025 6427 24091 6430
rect 26509 6490 26575 6493
rect 27705 6490 27771 6493
rect 31845 6490 31911 6493
rect 26509 6488 31911 6490
rect 26509 6432 26514 6488
rect 26570 6432 27710 6488
rect 27766 6432 31850 6488
rect 31906 6432 31911 6488
rect 26509 6430 31911 6432
rect 26509 6427 26575 6430
rect 27705 6427 27771 6430
rect 31845 6427 31911 6430
rect 16941 6354 17007 6357
rect 33225 6354 33291 6357
rect 16941 6352 33291 6354
rect 16941 6296 16946 6352
rect 17002 6296 33230 6352
rect 33286 6296 33291 6352
rect 16941 6294 33291 6296
rect 16941 6291 17007 6294
rect 33225 6291 33291 6294
rect 22001 6082 22067 6085
rect 25129 6082 25195 6085
rect 22001 6080 25195 6082
rect 22001 6024 22006 6080
rect 22062 6024 25134 6080
rect 25190 6024 25195 6080
rect 22001 6022 25195 6024
rect 22001 6019 22067 6022
rect 25129 6019 25195 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 59200 5992 60000 6112
rect 34930 5951 35246 5952
rect 1577 5946 1643 5949
rect 1577 5944 1962 5946
rect 1577 5888 1582 5944
rect 1638 5888 1962 5944
rect 1577 5886 1962 5888
rect 1577 5883 1643 5886
rect 0 5810 800 5840
rect 1761 5810 1827 5813
rect 0 5808 1827 5810
rect 0 5752 1766 5808
rect 1822 5752 1827 5808
rect 0 5750 1827 5752
rect 1902 5810 1962 5886
rect 22461 5810 22527 5813
rect 1902 5808 22527 5810
rect 1902 5752 22466 5808
rect 22522 5752 22527 5808
rect 1902 5750 22527 5752
rect 0 5720 800 5750
rect 1761 5747 1827 5750
rect 22461 5747 22527 5750
rect 25446 5748 25452 5812
rect 25516 5810 25522 5812
rect 25589 5810 25655 5813
rect 25516 5808 25655 5810
rect 25516 5752 25594 5808
rect 25650 5752 25655 5808
rect 25516 5750 25655 5752
rect 25516 5748 25522 5750
rect 25589 5747 25655 5750
rect 1945 5674 2011 5677
rect 24577 5674 24643 5677
rect 1945 5672 24643 5674
rect 1945 5616 1950 5672
rect 2006 5616 24582 5672
rect 24638 5616 24643 5672
rect 1945 5614 24643 5616
rect 1945 5611 2011 5614
rect 24577 5611 24643 5614
rect 25773 5674 25839 5677
rect 28625 5674 28691 5677
rect 25773 5672 28691 5674
rect 25773 5616 25778 5672
rect 25834 5616 28630 5672
rect 28686 5616 28691 5672
rect 25773 5614 28691 5616
rect 25773 5611 25839 5614
rect 28625 5611 28691 5614
rect 39481 5674 39547 5677
rect 40902 5674 40908 5676
rect 39481 5672 40908 5674
rect 39481 5616 39486 5672
rect 39542 5616 40908 5672
rect 39481 5614 40908 5616
rect 39481 5611 39547 5614
rect 40902 5612 40908 5614
rect 40972 5612 40978 5676
rect 57237 5538 57303 5541
rect 59200 5538 60000 5568
rect 57237 5536 60000 5538
rect 57237 5480 57242 5536
rect 57298 5480 60000 5536
rect 57237 5478 60000 5480
rect 57237 5475 57303 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 59200 5448 60000 5478
rect 50290 5407 50606 5408
rect 19793 5266 19859 5269
rect 24209 5266 24275 5269
rect 19793 5264 24275 5266
rect 19793 5208 19798 5264
rect 19854 5208 24214 5264
rect 24270 5208 24275 5264
rect 19793 5206 24275 5208
rect 19793 5203 19859 5206
rect 24209 5203 24275 5206
rect 0 5130 800 5160
rect 1761 5130 1827 5133
rect 0 5128 1827 5130
rect 0 5072 1766 5128
rect 1822 5072 1827 5128
rect 0 5070 1827 5072
rect 0 5040 800 5070
rect 1761 5067 1827 5070
rect 58065 4994 58131 4997
rect 59200 4994 60000 5024
rect 58065 4992 60000 4994
rect 58065 4936 58070 4992
rect 58126 4936 60000 4992
rect 58065 4934 60000 4936
rect 58065 4931 58131 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 59200 4904 60000 4934
rect 34930 4863 35246 4864
rect 22461 4858 22527 4861
rect 25129 4858 25195 4861
rect 22461 4856 25195 4858
rect 22461 4800 22466 4856
rect 22522 4800 25134 4856
rect 25190 4800 25195 4856
rect 22461 4798 25195 4800
rect 22461 4795 22527 4798
rect 25129 4795 25195 4798
rect 22829 4722 22895 4725
rect 24761 4722 24827 4725
rect 22829 4720 24827 4722
rect 22829 4664 22834 4720
rect 22890 4664 24766 4720
rect 24822 4664 24827 4720
rect 22829 4662 24827 4664
rect 22829 4659 22895 4662
rect 24761 4659 24827 4662
rect 14733 4586 14799 4589
rect 19149 4586 19215 4589
rect 14733 4584 19215 4586
rect 14733 4528 14738 4584
rect 14794 4528 19154 4584
rect 19210 4528 19215 4584
rect 14733 4526 19215 4528
rect 14733 4523 14799 4526
rect 19149 4523 19215 4526
rect 0 4450 800 4480
rect 1853 4450 1919 4453
rect 0 4448 1919 4450
rect 0 4392 1858 4448
rect 1914 4392 1919 4448
rect 0 4390 1919 4392
rect 0 4360 800 4390
rect 1853 4387 1919 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 59200 4360 60000 4480
rect 50290 4319 50606 4320
rect 13721 4042 13787 4045
rect 26969 4042 27035 4045
rect 13721 4040 27035 4042
rect 13721 3984 13726 4040
rect 13782 3984 26974 4040
rect 27030 3984 27035 4040
rect 13721 3982 27035 3984
rect 13721 3979 13787 3982
rect 26969 3979 27035 3982
rect 8293 3906 8359 3909
rect 18689 3906 18755 3909
rect 8293 3904 18755 3906
rect 8293 3848 8298 3904
rect 8354 3848 18694 3904
rect 18750 3848 18755 3904
rect 8293 3846 18755 3848
rect 8293 3843 8359 3846
rect 18689 3843 18755 3846
rect 18965 3906 19031 3909
rect 19241 3906 19307 3909
rect 24945 3906 25011 3909
rect 18965 3904 25011 3906
rect 18965 3848 18970 3904
rect 19026 3848 19246 3904
rect 19302 3848 24950 3904
rect 25006 3848 25011 3904
rect 18965 3846 25011 3848
rect 18965 3843 19031 3846
rect 19241 3843 19307 3846
rect 24945 3843 25011 3846
rect 58065 3906 58131 3909
rect 59200 3906 60000 3936
rect 58065 3904 60000 3906
rect 58065 3848 58070 3904
rect 58126 3848 60000 3904
rect 58065 3846 60000 3848
rect 58065 3843 58131 3846
rect 4210 3840 4526 3841
rect 0 3770 800 3800
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 59200 3816 60000 3846
rect 34930 3775 35246 3776
rect 1761 3770 1827 3773
rect 0 3768 1827 3770
rect 0 3712 1766 3768
rect 1822 3712 1827 3768
rect 0 3710 1827 3712
rect 0 3680 800 3710
rect 1761 3707 1827 3710
rect 9949 3770 10015 3773
rect 19241 3770 19307 3773
rect 9949 3768 19307 3770
rect 9949 3712 9954 3768
rect 10010 3712 19246 3768
rect 19302 3712 19307 3768
rect 9949 3710 19307 3712
rect 9949 3707 10015 3710
rect 19241 3707 19307 3710
rect 19425 3770 19491 3773
rect 22001 3770 22067 3773
rect 19425 3768 22067 3770
rect 19425 3712 19430 3768
rect 19486 3712 22006 3768
rect 22062 3712 22067 3768
rect 19425 3710 22067 3712
rect 19425 3707 19491 3710
rect 22001 3707 22067 3710
rect 42609 3770 42675 3773
rect 47117 3770 47183 3773
rect 42609 3768 47183 3770
rect 42609 3712 42614 3768
rect 42670 3712 47122 3768
rect 47178 3712 47183 3768
rect 42609 3710 47183 3712
rect 42609 3707 42675 3710
rect 47117 3707 47183 3710
rect 13721 3634 13787 3637
rect 25957 3634 26023 3637
rect 13721 3632 26023 3634
rect 13721 3576 13726 3632
rect 13782 3576 25962 3632
rect 26018 3576 26023 3632
rect 13721 3574 26023 3576
rect 13721 3571 13787 3574
rect 25957 3571 26023 3574
rect 40902 3572 40908 3636
rect 40972 3634 40978 3636
rect 41045 3634 41111 3637
rect 40972 3632 41111 3634
rect 40972 3576 41050 3632
rect 41106 3576 41111 3632
rect 40972 3574 41111 3576
rect 40972 3572 40978 3574
rect 41045 3571 41111 3574
rect 43713 3634 43779 3637
rect 50889 3634 50955 3637
rect 43713 3632 50955 3634
rect 43713 3576 43718 3632
rect 43774 3576 50894 3632
rect 50950 3576 50955 3632
rect 43713 3574 50955 3576
rect 43713 3571 43779 3574
rect 50889 3571 50955 3574
rect 11605 3498 11671 3501
rect 28901 3498 28967 3501
rect 11605 3496 28967 3498
rect 11605 3440 11610 3496
rect 11666 3440 28906 3496
rect 28962 3440 28967 3496
rect 11605 3438 28967 3440
rect 11605 3435 11671 3438
rect 28901 3435 28967 3438
rect 32990 3436 32996 3500
rect 33060 3498 33066 3500
rect 45185 3498 45251 3501
rect 33060 3496 45251 3498
rect 33060 3440 45190 3496
rect 45246 3440 45251 3496
rect 33060 3438 45251 3440
rect 33060 3436 33066 3438
rect 45185 3435 45251 3438
rect 18965 3362 19031 3365
rect 19149 3362 19215 3365
rect 18965 3360 19215 3362
rect 18965 3304 18970 3360
rect 19026 3304 19154 3360
rect 19210 3304 19215 3360
rect 18965 3302 19215 3304
rect 18965 3299 19031 3302
rect 19149 3299 19215 3302
rect 39113 3362 39179 3365
rect 43345 3362 43411 3365
rect 39113 3360 43411 3362
rect 39113 3304 39118 3360
rect 39174 3304 43350 3360
rect 43406 3304 43411 3360
rect 39113 3302 43411 3304
rect 39113 3299 39179 3302
rect 43345 3299 43411 3302
rect 58157 3362 58223 3365
rect 59200 3362 60000 3392
rect 58157 3360 60000 3362
rect 58157 3304 58162 3360
rect 58218 3304 60000 3360
rect 58157 3302 60000 3304
rect 58157 3299 58223 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 59200 3272 60000 3302
rect 50290 3231 50606 3232
rect 9673 3226 9739 3229
rect 10593 3226 10659 3229
rect 9673 3224 10659 3226
rect 9673 3168 9678 3224
rect 9734 3168 10598 3224
rect 10654 3168 10659 3224
rect 9673 3166 10659 3168
rect 9673 3163 9739 3166
rect 10593 3163 10659 3166
rect 17309 3226 17375 3229
rect 19241 3226 19307 3229
rect 17309 3224 19307 3226
rect 17309 3168 17314 3224
rect 17370 3168 19246 3224
rect 19302 3168 19307 3224
rect 17309 3166 19307 3168
rect 17309 3163 17375 3166
rect 19241 3163 19307 3166
rect 43069 3226 43135 3229
rect 46841 3226 46907 3229
rect 43069 3224 46907 3226
rect 43069 3168 43074 3224
rect 43130 3168 46846 3224
rect 46902 3168 46907 3224
rect 43069 3166 46907 3168
rect 43069 3163 43135 3166
rect 46841 3163 46907 3166
rect 0 3090 800 3120
rect 1853 3090 1919 3093
rect 0 3088 1919 3090
rect 0 3032 1858 3088
rect 1914 3032 1919 3088
rect 0 3030 1919 3032
rect 0 3000 800 3030
rect 1853 3027 1919 3030
rect 9673 3090 9739 3093
rect 12341 3090 12407 3093
rect 9673 3088 12407 3090
rect 9673 3032 9678 3088
rect 9734 3032 12346 3088
rect 12402 3032 12407 3088
rect 9673 3030 12407 3032
rect 9673 3027 9739 3030
rect 12341 3027 12407 3030
rect 17861 3090 17927 3093
rect 22277 3090 22343 3093
rect 17861 3088 22343 3090
rect 17861 3032 17866 3088
rect 17922 3032 22282 3088
rect 22338 3032 22343 3088
rect 17861 3030 22343 3032
rect 17861 3027 17927 3030
rect 22277 3027 22343 3030
rect 43345 3090 43411 3093
rect 45093 3090 45159 3093
rect 43345 3088 45159 3090
rect 43345 3032 43350 3088
rect 43406 3032 45098 3088
rect 45154 3032 45159 3088
rect 43345 3030 45159 3032
rect 43345 3027 43411 3030
rect 45093 3027 45159 3030
rect 45737 3090 45803 3093
rect 52453 3090 52519 3093
rect 45737 3088 52519 3090
rect 45737 3032 45742 3088
rect 45798 3032 52458 3088
rect 52514 3032 52519 3088
rect 45737 3030 52519 3032
rect 45737 3027 45803 3030
rect 52453 3027 52519 3030
rect 13537 2954 13603 2957
rect 20437 2954 20503 2957
rect 13537 2952 20503 2954
rect 13537 2896 13542 2952
rect 13598 2896 20442 2952
rect 20498 2896 20503 2952
rect 13537 2894 20503 2896
rect 13537 2891 13603 2894
rect 20437 2891 20503 2894
rect 44909 2954 44975 2957
rect 45645 2954 45711 2957
rect 44909 2952 45711 2954
rect 44909 2896 44914 2952
rect 44970 2896 45650 2952
rect 45706 2896 45711 2952
rect 44909 2894 45711 2896
rect 44909 2891 44975 2894
rect 45645 2891 45711 2894
rect 9581 2818 9647 2821
rect 11973 2818 12039 2821
rect 9581 2816 12039 2818
rect 9581 2760 9586 2816
rect 9642 2760 11978 2816
rect 12034 2760 12039 2816
rect 9581 2758 12039 2760
rect 9581 2755 9647 2758
rect 11973 2755 12039 2758
rect 58157 2818 58223 2821
rect 59200 2818 60000 2848
rect 58157 2816 60000 2818
rect 58157 2760 58162 2816
rect 58218 2760 60000 2816
rect 58157 2758 60000 2760
rect 58157 2755 58223 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 59200 2728 60000 2758
rect 34930 2687 35246 2688
rect 20069 2684 20135 2685
rect 20069 2680 20116 2684
rect 20180 2682 20186 2684
rect 20069 2624 20074 2680
rect 20069 2620 20116 2624
rect 20180 2622 20226 2682
rect 20180 2620 20186 2622
rect 20069 2619 20135 2620
rect 0 2410 800 2440
rect 1853 2410 1919 2413
rect 0 2408 1919 2410
rect 0 2352 1858 2408
rect 1914 2352 1919 2408
rect 0 2350 1919 2352
rect 0 2320 800 2350
rect 1853 2347 1919 2350
rect 24158 2348 24164 2412
rect 24228 2410 24234 2412
rect 47945 2410 48011 2413
rect 24228 2408 48011 2410
rect 24228 2352 47950 2408
rect 48006 2352 48011 2408
rect 24228 2350 48011 2352
rect 24228 2348 24234 2350
rect 47945 2347 48011 2350
rect 57329 2274 57395 2277
rect 59200 2274 60000 2304
rect 57329 2272 60000 2274
rect 57329 2216 57334 2272
rect 57390 2216 60000 2272
rect 57329 2214 60000 2216
rect 57329 2211 57395 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 59200 2184 60000 2214
rect 50290 2143 50606 2144
rect 56501 1730 56567 1733
rect 59200 1730 60000 1760
rect 56501 1728 60000 1730
rect 56501 1672 56506 1728
rect 56562 1672 60000 1728
rect 56501 1670 60000 1672
rect 56501 1667 56567 1670
rect 59200 1640 60000 1670
rect 56501 1186 56567 1189
rect 59200 1186 60000 1216
rect 56501 1184 60000 1186
rect 56501 1128 56506 1184
rect 56562 1128 60000 1184
rect 56501 1126 60000 1128
rect 56501 1123 56567 1126
rect 59200 1096 60000 1126
<< via3 >>
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 30972 61100 31036 61164
rect 19576 60956 19640 60960
rect 19576 60900 19580 60956
rect 19580 60900 19636 60956
rect 19636 60900 19640 60956
rect 19576 60896 19640 60900
rect 19656 60956 19720 60960
rect 19656 60900 19660 60956
rect 19660 60900 19716 60956
rect 19716 60900 19720 60956
rect 19656 60896 19720 60900
rect 19736 60956 19800 60960
rect 19736 60900 19740 60956
rect 19740 60900 19796 60956
rect 19796 60900 19800 60956
rect 19736 60896 19800 60900
rect 19816 60956 19880 60960
rect 19816 60900 19820 60956
rect 19820 60900 19876 60956
rect 19876 60900 19880 60956
rect 19816 60896 19880 60900
rect 50296 60956 50360 60960
rect 50296 60900 50300 60956
rect 50300 60900 50356 60956
rect 50356 60900 50360 60956
rect 50296 60896 50360 60900
rect 50376 60956 50440 60960
rect 50376 60900 50380 60956
rect 50380 60900 50436 60956
rect 50436 60900 50440 60956
rect 50376 60896 50440 60900
rect 50456 60956 50520 60960
rect 50456 60900 50460 60956
rect 50460 60900 50516 60956
rect 50516 60900 50520 60956
rect 50456 60896 50520 60900
rect 50536 60956 50600 60960
rect 50536 60900 50540 60956
rect 50540 60900 50596 60956
rect 50596 60900 50600 60956
rect 50536 60896 50600 60900
rect 32076 60828 32140 60892
rect 33180 60752 33244 60756
rect 33180 60696 33230 60752
rect 33230 60696 33244 60752
rect 33180 60692 33244 60696
rect 34652 60692 34716 60756
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 38148 57352 38212 57356
rect 38148 57296 38162 57352
rect 38162 57296 38212 57352
rect 38148 57292 38212 57296
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 35572 56612 35636 56676
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 18276 53076 18340 53140
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 28764 38660 28828 38724
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 20116 37708 20180 37772
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 20116 36076 20180 36140
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 31892 30092 31956 30156
rect 20116 29956 20180 30020
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 28580 29140 28644 29204
rect 24164 29064 24228 29068
rect 24164 29008 24178 29064
rect 24178 29008 24228 29064
rect 24164 29004 24228 29008
rect 31524 29004 31588 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 29500 24652 29564 24716
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 20116 21932 20180 21996
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 28764 20904 28828 20908
rect 28764 20848 28814 20904
rect 28814 20848 28828 20904
rect 28764 20844 28828 20848
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 28580 19408 28644 19412
rect 28580 19352 28594 19408
rect 28594 19352 28644 19408
rect 28580 19348 28644 19352
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 32996 17988 33060 18052
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 32076 17912 32140 17916
rect 32076 17856 32090 17912
rect 32090 17856 32140 17912
rect 32076 17852 32140 17856
rect 33180 17912 33244 17916
rect 33180 17856 33194 17912
rect 33194 17856 33244 17912
rect 33180 17852 33244 17856
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 31892 16628 31956 16692
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 18276 16144 18340 16148
rect 18276 16088 18290 16144
rect 18290 16088 18340 16144
rect 18276 16084 18340 16088
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 34652 15540 34716 15604
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 19380 15056 19444 15060
rect 19380 15000 19430 15056
rect 19430 15000 19444 15056
rect 19380 14996 19444 15000
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 38148 13636 38212 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 23612 13364 23676 13428
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 19380 11596 19444 11660
rect 30972 11596 31036 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 31524 9556 31588 9620
rect 35572 9556 35636 9620
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 24532 9012 24596 9076
rect 25452 8876 25516 8940
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 29500 8332 29564 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 23612 6896 23676 6900
rect 23612 6840 23626 6896
rect 23626 6840 23676 6896
rect 23612 6836 23676 6840
rect 24532 6896 24596 6900
rect 24532 6840 24582 6896
rect 24582 6840 24596 6896
rect 24532 6836 24596 6840
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 25452 5748 25516 5812
rect 40908 5612 40972 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 40908 3572 40972 3636
rect 32996 3436 33060 3500
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 20116 2680 20180 2684
rect 20116 2624 20130 2680
rect 20130 2624 20180 2680
rect 20116 2620 20180 2624
rect 24164 2348 24228 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 61504 4528 61520
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 19568 60960 19888 61520
rect 34928 61504 35248 61520
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 30971 61164 31037 61165
rect 30971 61100 30972 61164
rect 31036 61100 31037 61164
rect 30971 61099 31037 61100
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 59872 19888 60896
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 58784 19888 59808
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 18275 53140 18341 53141
rect 18275 53076 18276 53140
rect 18340 53076 18341 53140
rect 18275 53075 18341 53076
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 18278 16149 18338 53075
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 28763 38724 28829 38725
rect 28763 38660 28764 38724
rect 28828 38660 28829 38724
rect 28763 38659 28829 38660
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 20115 37772 20181 37773
rect 20115 37708 20116 37772
rect 20180 37708 20181 37772
rect 20115 37707 20181 37708
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 20118 36141 20178 37707
rect 20115 36140 20181 36141
rect 20115 36076 20116 36140
rect 20180 36076 20181 36140
rect 20115 36075 20181 36076
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 20118 30021 20178 36075
rect 20115 30020 20181 30021
rect 20115 29956 20116 30020
rect 20180 29956 20181 30020
rect 20115 29955 20181 29956
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 28579 29204 28645 29205
rect 28579 29140 28580 29204
rect 28644 29140 28645 29204
rect 28579 29139 28645 29140
rect 24163 29068 24229 29069
rect 24163 29004 24164 29068
rect 24228 29004 24229 29068
rect 24163 29003 24229 29004
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 20115 21996 20181 21997
rect 20115 21932 20116 21996
rect 20180 21932 20181 21996
rect 20115 21931 20181 21932
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 18275 16148 18341 16149
rect 18275 16084 18276 16148
rect 18340 16084 18341 16148
rect 18275 16083 18341 16084
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19379 15060 19445 15061
rect 19379 14996 19380 15060
rect 19444 14996 19445 15060
rect 19379 14995 19445 14996
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 19382 11661 19442 14995
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19379 11660 19445 11661
rect 19379 11596 19380 11660
rect 19444 11596 19445 11660
rect 19379 11595 19445 11596
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 20118 2685 20178 21931
rect 23611 13428 23677 13429
rect 23611 13364 23612 13428
rect 23676 13364 23677 13428
rect 23611 13363 23677 13364
rect 23614 6901 23674 13363
rect 23611 6900 23677 6901
rect 23611 6836 23612 6900
rect 23676 6836 23677 6900
rect 23611 6835 23677 6836
rect 20115 2684 20181 2685
rect 20115 2620 20116 2684
rect 20180 2620 20181 2684
rect 20115 2619 20181 2620
rect 24166 2413 24226 29003
rect 28582 19413 28642 29139
rect 28766 20909 28826 38659
rect 29499 24716 29565 24717
rect 29499 24652 29500 24716
rect 29564 24652 29565 24716
rect 29499 24651 29565 24652
rect 28763 20908 28829 20909
rect 28763 20844 28764 20908
rect 28828 20844 28829 20908
rect 28763 20843 28829 20844
rect 28579 19412 28645 19413
rect 28579 19348 28580 19412
rect 28644 19348 28645 19412
rect 28579 19347 28645 19348
rect 24531 9076 24597 9077
rect 24531 9012 24532 9076
rect 24596 9012 24597 9076
rect 24531 9011 24597 9012
rect 24534 6901 24594 9011
rect 25451 8940 25517 8941
rect 25451 8876 25452 8940
rect 25516 8876 25517 8940
rect 25451 8875 25517 8876
rect 24531 6900 24597 6901
rect 24531 6836 24532 6900
rect 24596 6836 24597 6900
rect 24531 6835 24597 6836
rect 25454 5813 25514 8875
rect 29502 8397 29562 24651
rect 30974 11661 31034 61099
rect 32075 60892 32141 60893
rect 32075 60828 32076 60892
rect 32140 60828 32141 60892
rect 32075 60827 32141 60828
rect 31891 30156 31957 30157
rect 31891 30092 31892 30156
rect 31956 30092 31957 30156
rect 31891 30091 31957 30092
rect 31523 29068 31589 29069
rect 31523 29004 31524 29068
rect 31588 29004 31589 29068
rect 31523 29003 31589 29004
rect 30971 11660 31037 11661
rect 30971 11596 30972 11660
rect 31036 11596 31037 11660
rect 30971 11595 31037 11596
rect 31526 9621 31586 29003
rect 31894 16693 31954 30091
rect 32078 17917 32138 60827
rect 33179 60756 33245 60757
rect 33179 60692 33180 60756
rect 33244 60692 33245 60756
rect 33179 60691 33245 60692
rect 34651 60756 34717 60757
rect 34651 60692 34652 60756
rect 34716 60692 34717 60756
rect 34651 60691 34717 60692
rect 32995 18052 33061 18053
rect 32995 17988 32996 18052
rect 33060 17988 33061 18052
rect 32995 17987 33061 17988
rect 32075 17916 32141 17917
rect 32075 17852 32076 17916
rect 32140 17852 32141 17916
rect 32075 17851 32141 17852
rect 31891 16692 31957 16693
rect 31891 16628 31892 16692
rect 31956 16628 31957 16692
rect 31891 16627 31957 16628
rect 31523 9620 31589 9621
rect 31523 9556 31524 9620
rect 31588 9556 31589 9620
rect 31523 9555 31589 9556
rect 29499 8396 29565 8397
rect 29499 8332 29500 8396
rect 29564 8332 29565 8396
rect 29499 8331 29565 8332
rect 25451 5812 25517 5813
rect 25451 5748 25452 5812
rect 25516 5748 25517 5812
rect 25451 5747 25517 5748
rect 32998 3501 33058 17987
rect 33182 17917 33242 60691
rect 33179 17916 33245 17917
rect 33179 17852 33180 17916
rect 33244 17852 33245 17916
rect 33179 17851 33245 17852
rect 34654 15605 34714 60691
rect 34928 60416 35248 61440
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 59328 35248 60352
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 57152 35248 58176
rect 50288 60960 50608 61520
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 59872 50608 60896
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 38147 57356 38213 57357
rect 38147 57292 38148 57356
rect 38212 57292 38213 57356
rect 38147 57291 38213 57292
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 35571 56676 35637 56677
rect 35571 56612 35572 56676
rect 35636 56612 35637 56676
rect 35571 56611 35637 56612
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34651 15604 34717 15605
rect 34651 15540 34652 15604
rect 34716 15540 34717 15604
rect 34651 15539 34717 15540
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 35574 9621 35634 56611
rect 38150 13701 38210 57291
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 38147 13700 38213 13701
rect 38147 13636 38148 13700
rect 38212 13636 38213 13700
rect 38147 13635 38213 13636
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 35571 9620 35637 9621
rect 35571 9556 35572 9620
rect 35636 9556 35637 9620
rect 35571 9555 35637 9556
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 40907 5676 40973 5677
rect 40907 5612 40908 5676
rect 40972 5612 40973 5676
rect 40907 5611 40973 5612
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 32995 3500 33061 3501
rect 32995 3436 32996 3500
rect 33060 3436 33061 3500
rect 32995 3435 33061 3436
rect 34928 2752 35248 3776
rect 40910 3637 40970 5611
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 40907 3636 40973 3637
rect 40907 3572 40908 3636
rect 40972 3572 40973 3636
rect 40907 3571 40973 3572
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 24163 2412 24229 2413
rect 24163 2348 24164 2412
rect 24228 2348 24229 2412
rect 24163 2347 24229 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2116 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1666464484
transform 1 0 43424 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1666464484
transform 1 0 18032 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1666464484
transform 1 0 22908 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1666464484
transform 1 0 19780 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1666464484
transform 1 0 14444 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1666464484
transform 1 0 22448 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1666464484
transform 1 0 23644 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1666464484
transform 1 0 18308 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1666464484
transform 1 0 20424 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1666464484
transform 1 0 20332 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1666464484
transform 1 0 1748 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1666464484
transform 1 0 23368 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1666464484
transform 1 0 38456 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1666464484
transform 1 0 25208 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1666464484
transform 1 0 33212 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1666464484
transform 1 0 25208 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1666464484
transform 1 0 25300 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1666464484
transform 1 0 20976 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1666464484
transform 1 0 19780 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1666464484
transform 1 0 28060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1666464484
transform 1 0 25392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1666464484
transform 1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1666464484
transform 1 0 53360 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1666464484
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1666464484
transform 1 0 46092 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1666464484
transform 1 0 20792 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1666464484
transform 1 0 28152 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1666464484
transform 1 0 34592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 2116 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41
timestamp 1666464484
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46
timestamp 1666464484
transform 1 0 5336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1666464484
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1666464484
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1666464484
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74
timestamp 1666464484
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1666464484
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1666464484
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1666464484
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1666464484
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122
timestamp 1666464484
transform 1 0 12328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_130
timestamp 1666464484
transform 1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1666464484
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1666464484
transform 1 0 14536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1666464484
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666464484
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174
timestamp 1666464484
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1666464484
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666464484
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1666464484
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1666464484
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666464484
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1666464484
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1666464484
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1666464484
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_258
timestamp 1666464484
transform 1 0 24840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_268
timestamp 1666464484
transform 1 0 25760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1666464484
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_289
timestamp 1666464484
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_296
timestamp 1666464484
transform 1 0 28336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1666464484
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_315
timestamp 1666464484
transform 1 0 30084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_322
timestamp 1666464484
transform 1 0 30728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1666464484
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_345
timestamp 1666464484
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1666464484
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1666464484
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1666464484
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1666464484
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1666464484
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1666464484
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1666464484
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_401
timestamp 1666464484
transform 1 0 37996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_411
timestamp 1666464484
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1666464484
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666464484
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_429
timestamp 1666464484
transform 1 0 40572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_439
timestamp 1666464484
transform 1 0 41492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1666464484
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666464484
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_457
timestamp 1666464484
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_470
timestamp 1666464484
transform 1 0 44344 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1666464484
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_487
timestamp 1666464484
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_497
timestamp 1666464484
transform 1 0 46828 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1666464484
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1666464484
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_513
timestamp 1666464484
transform 1 0 48300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_523
timestamp 1666464484
transform 1 0 49220 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1666464484
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1666464484
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_541
timestamp 1666464484
transform 1 0 50876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_551
timestamp 1666464484
transform 1 0 51796 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1666464484
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_561
timestamp 1666464484
transform 1 0 52716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_567
timestamp 1666464484
transform 1 0 53268 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1666464484
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_589
timestamp 1666464484
transform 1 0 55292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_595
timestamp 1666464484
transform 1 0 55844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_603
timestamp 1666464484
transform 1 0 56580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_607
timestamp 1666464484
transform 1 0 56948 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1666464484
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_617
timestamp 1666464484
transform 1 0 57868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_623
timestamp 1666464484
transform 1 0 58420 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1666464484
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_39
timestamp 1666464484
transform 1 0 4692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1666464484
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_65
timestamp 1666464484
transform 1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1666464484
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1666464484
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_100
timestamp 1666464484
transform 1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666464484
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_120
timestamp 1666464484
transform 1 0 12144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_128
timestamp 1666464484
transform 1 0 12880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1666464484
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_146
timestamp 1666464484
transform 1 0 14536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1666464484
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1666464484
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1666464484
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_191
timestamp 1666464484
transform 1 0 18676 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_211
timestamp 1666464484
transform 1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_215
timestamp 1666464484
transform 1 0 20884 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1666464484
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1666464484
transform 1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_259
timestamp 1666464484
transform 1 0 24932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_268
timestamp 1666464484
transform 1 0 25760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1666464484
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_289
timestamp 1666464484
transform 1 0 27692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_297
timestamp 1666464484
transform 1 0 28428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_314
timestamp 1666464484
transform 1 0 29992 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_322
timestamp 1666464484
transform 1 0 30728 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1666464484
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1666464484
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_345
timestamp 1666464484
transform 1 0 32844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_355
timestamp 1666464484
transform 1 0 33764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_365
timestamp 1666464484
transform 1 0 34684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_375
timestamp 1666464484
transform 1 0 35604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1666464484
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1666464484
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1666464484
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_401
timestamp 1666464484
transform 1 0 37996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_411
timestamp 1666464484
transform 1 0 38916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_421
timestamp 1666464484
transform 1 0 39836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1666464484
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1666464484
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1666464484
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1666464484
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_457
timestamp 1666464484
transform 1 0 43148 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_465
timestamp 1666464484
transform 1 0 43884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_484
timestamp 1666464484
transform 1 0 45632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_492
timestamp 1666464484
transform 1 0 46368 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1666464484
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1666464484
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_511
timestamp 1666464484
transform 1 0 48116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_521
timestamp 1666464484
transform 1 0 49036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_531
timestamp 1666464484
transform 1 0 49956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_539
timestamp 1666464484
transform 1 0 50692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_547
timestamp 1666464484
transform 1 0 51428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_555
timestamp 1666464484
transform 1 0 52164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1666464484
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1666464484
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_567
timestamp 1666464484
transform 1 0 53268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_575
timestamp 1666464484
transform 1 0 54004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_583
timestamp 1666464484
transform 1 0 54740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_591
timestamp 1666464484
transform 1 0 55476 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_599
timestamp 1666464484
transform 1 0 56212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_604
timestamp 1666464484
transform 1 0 56672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1666464484
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_617
timestamp 1666464484
transform 1 0 57868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_623
timestamp 1666464484
transform 1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_11
timestamp 1666464484
transform 1 0 2116 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1666464484
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1666464484
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1666464484
transform 1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_61
timestamp 1666464484
transform 1 0 6716 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1666464484
transform 1 0 7176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1666464484
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1666464484
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_100
timestamp 1666464484
transform 1 0 10304 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_108
timestamp 1666464484
transform 1 0 11040 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1666464484
transform 1 0 11684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_125
timestamp 1666464484
transform 1 0 12604 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_131
timestamp 1666464484
transform 1 0 13156 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1666464484
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_147
timestamp 1666464484
transform 1 0 14628 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154
timestamp 1666464484
transform 1 0 15272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_164
timestamp 1666464484
transform 1 0 16192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_174
timestamp 1666464484
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1666464484
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1666464484
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1666464484
transform 1 0 20884 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_223
timestamp 1666464484
transform 1 0 21620 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1666464484
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1666464484
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1666464484
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_264
timestamp 1666464484
transform 1 0 25392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_284
timestamp 1666464484
transform 1 0 27232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_288
timestamp 1666464484
transform 1 0 27600 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_292
timestamp 1666464484
transform 1 0 27968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1666464484
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1666464484
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_323
timestamp 1666464484
transform 1 0 30820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_327
timestamp 1666464484
transform 1 0 31188 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_332
timestamp 1666464484
transform 1 0 31648 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_353
timestamp 1666464484
transform 1 0 33580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_361
timestamp 1666464484
transform 1 0 34316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1666464484
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_373
timestamp 1666464484
transform 1 0 35420 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_383
timestamp 1666464484
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_393
timestamp 1666464484
transform 1 0 37260 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_401
timestamp 1666464484
transform 1 0 37996 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_410
timestamp 1666464484
transform 1 0 38824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1666464484
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1666464484
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_427
timestamp 1666464484
transform 1 0 40388 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_439
timestamp 1666464484
transform 1 0 41492 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_457
timestamp 1666464484
transform 1 0 43148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_470
timestamp 1666464484
transform 1 0 44344 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1666464484
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_496
timestamp 1666464484
transform 1 0 46736 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_504
timestamp 1666464484
transform 1 0 47472 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1666464484
transform 1 0 48208 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_520
timestamp 1666464484
transform 1 0 48944 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_530
timestamp 1666464484
transform 1 0 49864 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_533
timestamp 1666464484
transform 1 0 50140 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_539
timestamp 1666464484
transform 1 0 50692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_547
timestamp 1666464484
transform 1 0 51428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_555
timestamp 1666464484
transform 1 0 52164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_563
timestamp 1666464484
transform 1 0 52900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_571
timestamp 1666464484
transform 1 0 53636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_579
timestamp 1666464484
transform 1 0 54372 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1666464484
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_589
timestamp 1666464484
transform 1 0 55292 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_602
timestamp 1666464484
transform 1 0 56488 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_622
timestamp 1666464484
transform 1 0 58328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_11
timestamp 1666464484
transform 1 0 2116 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_23
timestamp 1666464484
transform 1 0 3220 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_35
timestamp 1666464484
transform 1 0 4324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1666464484
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_65
timestamp 1666464484
transform 1 0 7084 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_70
timestamp 1666464484
transform 1 0 7544 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_78
timestamp 1666464484
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1666464484
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 1666464484
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1666464484
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1666464484
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 1666464484
transform 1 0 12788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_131
timestamp 1666464484
transform 1 0 13156 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1666464484
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_146
timestamp 1666464484
transform 1 0 14536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_156
timestamp 1666464484
transform 1 0 15456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1666464484
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_177
timestamp 1666464484
transform 1 0 17388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1666464484
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_198
timestamp 1666464484
transform 1 0 19320 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_211
timestamp 1666464484
transform 1 0 20516 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_215
timestamp 1666464484
transform 1 0 20884 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666464484
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_243
timestamp 1666464484
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_247
timestamp 1666464484
transform 1 0 23828 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_264
timestamp 1666464484
transform 1 0 25392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp 1666464484
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_292
timestamp 1666464484
transform 1 0 27968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_296
timestamp 1666464484
transform 1 0 28336 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_302
timestamp 1666464484
transform 1 0 28888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_315
timestamp 1666464484
transform 1 0 30084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_323
timestamp 1666464484
transform 1 0 30820 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1666464484
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_343
timestamp 1666464484
transform 1 0 32660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_351
timestamp 1666464484
transform 1 0 33396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_360
timestamp 1666464484
transform 1 0 34224 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_373
timestamp 1666464484
transform 1 0 35420 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_383
timestamp 1666464484
transform 1 0 36340 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1666464484
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1666464484
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_401
timestamp 1666464484
transform 1 0 37996 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_409
timestamp 1666464484
transform 1 0 38732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_417
timestamp 1666464484
transform 1 0 39468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_425
timestamp 1666464484
transform 1 0 40204 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_433
timestamp 1666464484
transform 1 0 40940 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_439
timestamp 1666464484
transform 1 0 41492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_446
timestamp 1666464484
transform 1 0 42136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_449
timestamp 1666464484
transform 1 0 42412 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_465
timestamp 1666464484
transform 1 0 43884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_473
timestamp 1666464484
transform 1 0 44620 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_492
timestamp 1666464484
transform 1 0 46368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_500
timestamp 1666464484
transform 1 0 47104 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_505
timestamp 1666464484
transform 1 0 47564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_511
timestamp 1666464484
transform 1 0 48116 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_519
timestamp 1666464484
transform 1 0 48852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_531
timestamp 1666464484
transform 1 0 49956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_543
timestamp 1666464484
transform 1 0 51060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_555
timestamp 1666464484
transform 1 0 52164 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1666464484
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1666464484
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1666464484
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_585
timestamp 1666464484
transform 1 0 54924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_589
timestamp 1666464484
transform 1 0 55292 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_593
timestamp 1666464484
transform 1 0 55660 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_613
timestamp 1666464484
transform 1 0 57500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_617
timestamp 1666464484
transform 1 0 57868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_623
timestamp 1666464484
transform 1 0 58420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_11
timestamp 1666464484
transform 1 0 2116 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1666464484
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1666464484
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_65
timestamp 1666464484
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_72
timestamp 1666464484
transform 1 0 7728 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1666464484
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp 1666464484
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_96
timestamp 1666464484
transform 1 0 9936 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_102
timestamp 1666464484
transform 1 0 10488 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_110
timestamp 1666464484
transform 1 0 11224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_121
timestamp 1666464484
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_131
timestamp 1666464484
transform 1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1666464484
transform 1 0 14444 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_152
timestamp 1666464484
transform 1 0 15088 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_160
timestamp 1666464484
transform 1 0 15824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_179
timestamp 1666464484
transform 1 0 17572 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1666464484
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_209
timestamp 1666464484
transform 1 0 20332 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_218
timestamp 1666464484
transform 1 0 21160 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_228
timestamp 1666464484
transform 1 0 22080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_241
timestamp 1666464484
transform 1 0 23276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 1666464484
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_264
timestamp 1666464484
transform 1 0 25392 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_272
timestamp 1666464484
transform 1 0 26128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_278
timestamp 1666464484
transform 1 0 26680 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_285
timestamp 1666464484
transform 1 0 27324 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_292
timestamp 1666464484
transform 1 0 27968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_299
timestamp 1666464484
transform 1 0 28612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1666464484
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_333
timestamp 1666464484
transform 1 0 31740 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_342
timestamp 1666464484
transform 1 0 32568 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_350
timestamp 1666464484
transform 1 0 33304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_356
timestamp 1666464484
transform 1 0 33856 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1666464484
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_373
timestamp 1666464484
transform 1 0 35420 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_379
timestamp 1666464484
transform 1 0 35972 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_386
timestamp 1666464484
transform 1 0 36616 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_398
timestamp 1666464484
transform 1 0 37720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_406
timestamp 1666464484
transform 1 0 38456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_414
timestamp 1666464484
transform 1 0 39192 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_421
timestamp 1666464484
transform 1 0 39836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_427
timestamp 1666464484
transform 1 0 40388 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_435
timestamp 1666464484
transform 1 0 41124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_443
timestamp 1666464484
transform 1 0 41860 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_451
timestamp 1666464484
transform 1 0 42596 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_461
timestamp 1666464484
transform 1 0 43516 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_471
timestamp 1666464484
transform 1 0 44436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1666464484
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_477
timestamp 1666464484
transform 1 0 44988 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_483
timestamp 1666464484
transform 1 0 45540 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_491
timestamp 1666464484
transform 1 0 46276 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_499
timestamp 1666464484
transform 1 0 47012 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_507
timestamp 1666464484
transform 1 0 47748 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_515
timestamp 1666464484
transform 1 0 48484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_527
timestamp 1666464484
transform 1 0 49588 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1666464484
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1666464484
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1666464484
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1666464484
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1666464484
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1666464484
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1666464484
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1666464484
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_601
timestamp 1666464484
transform 1 0 56396 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_614
timestamp 1666464484
transform 1 0 57592 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_623
timestamp 1666464484
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_11
timestamp 1666464484
transform 1 0 2116 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_23
timestamp 1666464484
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_35
timestamp 1666464484
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1666464484
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1666464484
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_93
timestamp 1666464484
transform 1 0 9660 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_97
timestamp 1666464484
transform 1 0 10028 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_102
timestamp 1666464484
transform 1 0 10488 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1666464484
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_119
timestamp 1666464484
transform 1 0 12052 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_124
timestamp 1666464484
transform 1 0 12512 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_132
timestamp 1666464484
transform 1 0 13248 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1666464484
transform 1 0 13892 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1666464484
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1666464484
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1666464484
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_182
timestamp 1666464484
transform 1 0 17848 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_186
timestamp 1666464484
transform 1 0 18216 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1666464484
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_207
timestamp 1666464484
transform 1 0 20148 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_215
timestamp 1666464484
transform 1 0 20884 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp 1666464484
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_231
timestamp 1666464484
transform 1 0 22356 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_238
timestamp 1666464484
transform 1 0 23000 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_259
timestamp 1666464484
transform 1 0 24932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_265
timestamp 1666464484
transform 1 0 25484 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_271
timestamp 1666464484
transform 1 0 26036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1666464484
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_287
timestamp 1666464484
transform 1 0 27508 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_312
timestamp 1666464484
transform 1 0 29808 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_327
timestamp 1666464484
transform 1 0 31188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1666464484
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_348
timestamp 1666464484
transform 1 0 33120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_356
timestamp 1666464484
transform 1 0 33856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_362
timestamp 1666464484
transform 1 0 34408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_367
timestamp 1666464484
transform 1 0 34868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_375
timestamp 1666464484
transform 1 0 35604 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1666464484
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1666464484
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_399
timestamp 1666464484
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_407
timestamp 1666464484
transform 1 0 38548 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_415
timestamp 1666464484
transform 1 0 39284 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_423
timestamp 1666464484
transform 1 0 40020 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_431
timestamp 1666464484
transform 1 0 40756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_443
timestamp 1666464484
transform 1 0 41860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1666464484
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_449
timestamp 1666464484
transform 1 0 42412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_455
timestamp 1666464484
transform 1 0 42964 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_463
timestamp 1666464484
transform 1 0 43700 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_468
timestamp 1666464484
transform 1 0 44160 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_476
timestamp 1666464484
transform 1 0 44896 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_488
timestamp 1666464484
transform 1 0 46000 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1666464484
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1666464484
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1666464484
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1666464484
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1666464484
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1666464484
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1666464484
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1666464484
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1666464484
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1666464484
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_597
timestamp 1666464484
transform 1 0 56028 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_610
timestamp 1666464484
transform 1 0 57224 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_617
timestamp 1666464484
transform 1 0 57868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_623
timestamp 1666464484
transform 1 0 58420 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1666464484
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1666464484
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1666464484
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1666464484
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_115
timestamp 1666464484
transform 1 0 11684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_120
timestamp 1666464484
transform 1 0 12144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_124
timestamp 1666464484
transform 1 0 12512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_129
timestamp 1666464484
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1666464484
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_147
timestamp 1666464484
transform 1 0 14628 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_159
timestamp 1666464484
transform 1 0 15732 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_171
timestamp 1666464484
transform 1 0 16836 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_177
timestamp 1666464484
transform 1 0 17388 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_181
timestamp 1666464484
transform 1 0 17756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1666464484
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_215
timestamp 1666464484
transform 1 0 20884 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_227
timestamp 1666464484
transform 1 0 21988 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_231
timestamp 1666464484
transform 1 0 22356 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_239
timestamp 1666464484
transform 1 0 23092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1666464484
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_262
timestamp 1666464484
transform 1 0 25208 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_273
timestamp 1666464484
transform 1 0 26220 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_285
timestamp 1666464484
transform 1 0 27324 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_299
timestamp 1666464484
transform 1 0 28612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1666464484
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_322
timestamp 1666464484
transform 1 0 30728 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_334
timestamp 1666464484
transform 1 0 31832 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_342
timestamp 1666464484
transform 1 0 32568 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_354
timestamp 1666464484
transform 1 0 33672 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1666464484
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1666464484
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_371
timestamp 1666464484
transform 1 0 35236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_379
timestamp 1666464484
transform 1 0 35972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_383
timestamp 1666464484
transform 1 0 36340 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1666464484
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1666464484
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1666464484
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1666464484
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1666464484
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1666464484
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1666464484
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1666464484
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1666464484
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1666464484
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1666464484
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1666464484
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1666464484
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1666464484
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1666464484
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1666464484
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1666464484
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1666464484
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1666464484
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1666464484
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1666464484
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_601
timestamp 1666464484
transform 1 0 56396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_613
timestamp 1666464484
transform 1 0 57500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_623
timestamp 1666464484
transform 1 0 58420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_11
timestamp 1666464484
transform 1 0 2116 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_23
timestamp 1666464484
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_35
timestamp 1666464484
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_47
timestamp 1666464484
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1666464484
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1666464484
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_101
timestamp 1666464484
transform 1 0 10396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1666464484
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_121
timestamp 1666464484
transform 1 0 12236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_133
timestamp 1666464484
transform 1 0 13340 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_142
timestamp 1666464484
transform 1 0 14168 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_154
timestamp 1666464484
transform 1 0 15272 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1666464484
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_181
timestamp 1666464484
transform 1 0 17756 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1666464484
transform 1 0 18676 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_211
timestamp 1666464484
transform 1 0 20516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_239
timestamp 1666464484
transform 1 0 23092 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_250
timestamp 1666464484
transform 1 0 24104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_263
timestamp 1666464484
transform 1 0 25300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_267
timestamp 1666464484
transform 1 0 25668 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1666464484
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_292
timestamp 1666464484
transform 1 0 27968 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_298
timestamp 1666464484
transform 1 0 28520 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_318
timestamp 1666464484
transform 1 0 30360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_322
timestamp 1666464484
transform 1 0 30728 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_328
timestamp 1666464484
transform 1 0 31280 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_343
timestamp 1666464484
transform 1 0 32660 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1666464484
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_373
timestamp 1666464484
transform 1 0 35420 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp 1666464484
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1666464484
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_401
timestamp 1666464484
transform 1 0 37996 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_413
timestamp 1666464484
transform 1 0 39100 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_425
timestamp 1666464484
transform 1 0 40204 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_437
timestamp 1666464484
transform 1 0 41308 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_445
timestamp 1666464484
transform 1 0 42044 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1666464484
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1666464484
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1666464484
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1666464484
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1666464484
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666464484
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1666464484
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1666464484
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1666464484
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1666464484
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1666464484
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1666464484
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1666464484
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1666464484
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1666464484
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1666464484
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_609
timestamp 1666464484
transform 1 0 57132 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_614
timestamp 1666464484
transform 1 0 57592 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1666464484
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_11
timestamp 1666464484
transform 1 0 2116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1666464484
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1666464484
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1666464484
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_99
timestamp 1666464484
transform 1 0 10212 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_107
timestamp 1666464484
transform 1 0 10948 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_115
timestamp 1666464484
transform 1 0 11684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_127
timestamp 1666464484
transform 1 0 12788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_131
timestamp 1666464484
transform 1 0 13156 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1666464484
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_149
timestamp 1666464484
transform 1 0 14812 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_156
timestamp 1666464484
transform 1 0 15456 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_168
timestamp 1666464484
transform 1 0 16560 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_180
timestamp 1666464484
transform 1 0 17664 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1666464484
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_210
timestamp 1666464484
transform 1 0 20424 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_222
timestamp 1666464484
transform 1 0 21528 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_230
timestamp 1666464484
transform 1 0 22264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_238
timestamp 1666464484
transform 1 0 23000 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1666464484
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_262
timestamp 1666464484
transform 1 0 25208 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1666464484
transform 1 0 26312 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_291
timestamp 1666464484
transform 1 0 27876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_295
timestamp 1666464484
transform 1 0 28244 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1666464484
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_321
timestamp 1666464484
transform 1 0 30636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_332
timestamp 1666464484
transform 1 0 31648 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_340
timestamp 1666464484
transform 1 0 32384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_348
timestamp 1666464484
transform 1 0 33120 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_356
timestamp 1666464484
transform 1 0 33856 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1666464484
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_365
timestamp 1666464484
transform 1 0 34684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_380
timestamp 1666464484
transform 1 0 36064 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_384
timestamp 1666464484
transform 1 0 36432 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_394
timestamp 1666464484
transform 1 0 37352 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_398
timestamp 1666464484
transform 1 0 37720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_407
timestamp 1666464484
transform 1 0 38548 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_414
timestamp 1666464484
transform 1 0 39192 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1666464484
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1666464484
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1666464484
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1666464484
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1666464484
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1666464484
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1666464484
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1666464484
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1666464484
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1666464484
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1666464484
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1666464484
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1666464484
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1666464484
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1666464484
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1666464484
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1666464484
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1666464484
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1666464484
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_601
timestamp 1666464484
transform 1 0 56396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_605
timestamp 1666464484
transform 1 0 56764 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_622
timestamp 1666464484
transform 1 0 58328 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_11
timestamp 1666464484
transform 1 0 2116 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_23
timestamp 1666464484
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1666464484
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1666464484
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1666464484
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1666464484
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1666464484
transform 1 0 12420 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_133
timestamp 1666464484
transform 1 0 13340 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_145
timestamp 1666464484
transform 1 0 14444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_157
timestamp 1666464484
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1666464484
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_181
timestamp 1666464484
transform 1 0 17756 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_191
timestamp 1666464484
transform 1 0 18676 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_203
timestamp 1666464484
transform 1 0 19780 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_214
timestamp 1666464484
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1666464484
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_237
timestamp 1666464484
transform 1 0 22908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_241
timestamp 1666464484
transform 1 0 23276 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_262
timestamp 1666464484
transform 1 0 25208 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_274
timestamp 1666464484
transform 1 0 26312 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_309
timestamp 1666464484
transform 1 0 29532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1666464484
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_342
timestamp 1666464484
transform 1 0 32568 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_351
timestamp 1666464484
transform 1 0 33396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_362
timestamp 1666464484
transform 1 0 34408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_366
timestamp 1666464484
transform 1 0 34776 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_376
timestamp 1666464484
transform 1 0 35696 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp 1666464484
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_393
timestamp 1666464484
transform 1 0 37260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_403
timestamp 1666464484
transform 1 0 38180 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_407
timestamp 1666464484
transform 1 0 38548 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_415
timestamp 1666464484
transform 1 0 39284 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_422
timestamp 1666464484
transform 1 0 39928 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_434
timestamp 1666464484
transform 1 0 41032 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1666464484
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1666464484
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1666464484
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1666464484
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1666464484
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1666464484
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1666464484
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1666464484
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1666464484
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1666464484
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1666464484
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1666464484
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1666464484
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1666464484
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1666464484
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1666464484
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_597
timestamp 1666464484
transform 1 0 56028 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_604
timestamp 1666464484
transform 1 0 56672 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_614
timestamp 1666464484
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_617
timestamp 1666464484
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_623
timestamp 1666464484
transform 1 0 58420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_11
timestamp 1666464484
transform 1 0 2116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1666464484
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1666464484
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1666464484
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1666464484
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_113
timestamp 1666464484
transform 1 0 11500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_120
timestamp 1666464484
transform 1 0 12144 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_132
timestamp 1666464484
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1666464484
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_169
timestamp 1666464484
transform 1 0 16652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_178
timestamp 1666464484
transform 1 0 17480 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_186
timestamp 1666464484
transform 1 0 18216 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1666464484
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_216
timestamp 1666464484
transform 1 0 20976 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_228
timestamp 1666464484
transform 1 0 22080 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_240
timestamp 1666464484
transform 1 0 23184 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1666464484
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_277
timestamp 1666464484
transform 1 0 26588 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_290
timestamp 1666464484
transform 1 0 27784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_300
timestamp 1666464484
transform 1 0 28704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_318
timestamp 1666464484
transform 1 0 30360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_329
timestamp 1666464484
transform 1 0 31372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_342
timestamp 1666464484
transform 1 0 32568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_355
timestamp 1666464484
transform 1 0 33764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666464484
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1666464484
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_386
timestamp 1666464484
transform 1 0 36616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_397
timestamp 1666464484
transform 1 0 37628 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_412
timestamp 1666464484
transform 1 0 39008 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_421
timestamp 1666464484
transform 1 0 39836 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_428
timestamp 1666464484
transform 1 0 40480 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_440
timestamp 1666464484
transform 1 0 41584 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_452
timestamp 1666464484
transform 1 0 42688 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_464
timestamp 1666464484
transform 1 0 43792 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1666464484
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1666464484
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1666464484
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1666464484
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1666464484
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1666464484
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1666464484
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1666464484
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1666464484
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1666464484
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1666464484
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1666464484
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_589
timestamp 1666464484
transform 1 0 55292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_594
timestamp 1666464484
transform 1 0 55752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_602
timestamp 1666464484
transform 1 0 56488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_622
timestamp 1666464484
transform 1 0 58328 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1666464484
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1666464484
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1666464484
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1666464484
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1666464484
transform 1 0 12420 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_134
timestamp 1666464484
transform 1 0 13432 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_146
timestamp 1666464484
transform 1 0 14536 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_158
timestamp 1666464484
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1666464484
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_181
timestamp 1666464484
transform 1 0 17756 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_191
timestamp 1666464484
transform 1 0 18676 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_211
timestamp 1666464484
transform 1 0 20516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_237
timestamp 1666464484
transform 1 0 22908 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_265
timestamp 1666464484
transform 1 0 25484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_278
timestamp 1666464484
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_289
timestamp 1666464484
transform 1 0 27692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_297
timestamp 1666464484
transform 1 0 28428 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_306
timestamp 1666464484
transform 1 0 29256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_313
timestamp 1666464484
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_323
timestamp 1666464484
transform 1 0 30820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1666464484
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_341
timestamp 1666464484
transform 1 0 32476 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_345
timestamp 1666464484
transform 1 0 32844 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_357
timestamp 1666464484
transform 1 0 33948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_369
timestamp 1666464484
transform 1 0 35052 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_379
timestamp 1666464484
transform 1 0 35972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1666464484
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_393
timestamp 1666464484
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_399
timestamp 1666464484
transform 1 0 37812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_412
timestamp 1666464484
transform 1 0 39008 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_426
timestamp 1666464484
transform 1 0 40296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_438
timestamp 1666464484
transform 1 0 41400 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_446
timestamp 1666464484
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1666464484
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1666464484
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1666464484
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1666464484
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1666464484
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1666464484
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1666464484
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1666464484
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1666464484
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1666464484
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1666464484
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1666464484
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1666464484
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1666464484
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1666464484
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_597
timestamp 1666464484
transform 1 0 56028 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_604
timestamp 1666464484
transform 1 0 56672 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_614
timestamp 1666464484
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_617
timestamp 1666464484
transform 1 0 57868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_623
timestamp 1666464484
transform 1 0 58420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_11
timestamp 1666464484
transform 1 0 2116 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1666464484
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1666464484
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1666464484
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1666464484
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1666464484
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1666464484
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1666464484
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_215
timestamp 1666464484
transform 1 0 20884 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_227
timestamp 1666464484
transform 1 0 21988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_239
timestamp 1666464484
transform 1 0 23092 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_243
timestamp 1666464484
transform 1 0 23460 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1666464484
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_271
timestamp 1666464484
transform 1 0 26036 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_283
timestamp 1666464484
transform 1 0 27140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_295
timestamp 1666464484
transform 1 0 28244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1666464484
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_317
timestamp 1666464484
transform 1 0 30268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_328
timestamp 1666464484
transform 1 0 31280 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_338
timestamp 1666464484
transform 1 0 32200 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1666464484
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1666464484
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666464484
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_365
timestamp 1666464484
transform 1 0 34684 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_375
timestamp 1666464484
transform 1 0 35604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_387
timestamp 1666464484
transform 1 0 36708 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_391
timestamp 1666464484
transform 1 0 37076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_396
timestamp 1666464484
transform 1 0 37536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_404
timestamp 1666464484
transform 1 0 38272 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_408
timestamp 1666464484
transform 1 0 38640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_415
timestamp 1666464484
transform 1 0 39284 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1666464484
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_421
timestamp 1666464484
transform 1 0 39836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_430
timestamp 1666464484
transform 1 0 40664 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_439
timestamp 1666464484
transform 1 0 41492 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_451
timestamp 1666464484
transform 1 0 42596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_463
timestamp 1666464484
transform 1 0 43700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1666464484
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1666464484
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1666464484
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1666464484
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1666464484
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1666464484
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1666464484
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1666464484
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1666464484
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1666464484
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1666464484
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1666464484
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1666464484
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1666464484
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_601
timestamp 1666464484
transform 1 0 56396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_605
timestamp 1666464484
transform 1 0 56764 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_622
timestamp 1666464484
transform 1 0 58328 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_11
timestamp 1666464484
transform 1 0 2116 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_23
timestamp 1666464484
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_35
timestamp 1666464484
transform 1 0 4324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1666464484
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666464484
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1666464484
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1666464484
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_121
timestamp 1666464484
transform 1 0 12236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_129
timestamp 1666464484
transform 1 0 12972 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_146
timestamp 1666464484
transform 1 0 14536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1666464484
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1666464484
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1666464484
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_208
timestamp 1666464484
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1666464484
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1666464484
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1666464484
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666464484
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_291
timestamp 1666464484
transform 1 0 27876 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_298
timestamp 1666464484
transform 1 0 28520 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_310
timestamp 1666464484
transform 1 0 29624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_318
timestamp 1666464484
transform 1 0 30360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_330
timestamp 1666464484
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1666464484
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_361
timestamp 1666464484
transform 1 0 34316 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_367
timestamp 1666464484
transform 1 0 34868 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_377
timestamp 1666464484
transform 1 0 35788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_389
timestamp 1666464484
transform 1 0 36892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_393
timestamp 1666464484
transform 1 0 37260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_399
timestamp 1666464484
transform 1 0 37812 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_403
timestamp 1666464484
transform 1 0 38180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_415
timestamp 1666464484
transform 1 0 39284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_424
timestamp 1666464484
transform 1 0 40112 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_444
timestamp 1666464484
transform 1 0 41952 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1666464484
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1666464484
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1666464484
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1666464484
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1666464484
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1666464484
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1666464484
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1666464484
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1666464484
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1666464484
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1666464484
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1666464484
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1666464484
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1666464484
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1666464484
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1666464484
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_609
timestamp 1666464484
transform 1 0 57132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_614
timestamp 1666464484
transform 1 0 57592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1666464484
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_11
timestamp 1666464484
transform 1 0 2116 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1666464484
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1666464484
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1666464484
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1666464484
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_121
timestamp 1666464484
transform 1 0 12236 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_149
timestamp 1666464484
transform 1 0 14812 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_161
timestamp 1666464484
transform 1 0 15916 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_173
timestamp 1666464484
transform 1 0 17020 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_185
timestamp 1666464484
transform 1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1666464484
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_209
timestamp 1666464484
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_227
timestamp 1666464484
transform 1 0 21988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_239
timestamp 1666464484
transform 1 0 23092 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_243
timestamp 1666464484
transform 1 0 23460 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1666464484
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_281
timestamp 1666464484
transform 1 0 26956 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_305
timestamp 1666464484
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_320
timestamp 1666464484
transform 1 0 30544 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_343
timestamp 1666464484
transform 1 0 32660 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_355
timestamp 1666464484
transform 1 0 33764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666464484
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1666464484
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1666464484
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_389
timestamp 1666464484
transform 1 0 36892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_397
timestamp 1666464484
transform 1 0 37628 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_408
timestamp 1666464484
transform 1 0 38640 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_421
timestamp 1666464484
transform 1 0 39836 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_431
timestamp 1666464484
transform 1 0 40756 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_443
timestamp 1666464484
transform 1 0 41860 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_455
timestamp 1666464484
transform 1 0 42964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_467
timestamp 1666464484
transform 1 0 44068 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1666464484
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1666464484
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1666464484
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1666464484
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1666464484
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1666464484
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1666464484
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1666464484
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1666464484
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1666464484
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1666464484
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1666464484
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1666464484
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1666464484
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_601
timestamp 1666464484
transform 1 0 56396 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_613
timestamp 1666464484
transform 1 0 57500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_623
timestamp 1666464484
transform 1 0 58420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp 1666464484
transform 1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1666464484
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1666464484
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1666464484
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1666464484
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1666464484
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_125
timestamp 1666464484
transform 1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_135
timestamp 1666464484
transform 1 0 13524 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_147
timestamp 1666464484
transform 1 0 14628 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_155
timestamp 1666464484
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_175
timestamp 1666464484
transform 1 0 17204 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_185
timestamp 1666464484
transform 1 0 18124 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_197
timestamp 1666464484
transform 1 0 19228 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_205
timestamp 1666464484
transform 1 0 19964 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1666464484
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_236
timestamp 1666464484
transform 1 0 22816 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_244
timestamp 1666464484
transform 1 0 23552 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1666464484
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1666464484
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_302
timestamp 1666464484
transform 1 0 28888 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_309
timestamp 1666464484
transform 1 0 29532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_321
timestamp 1666464484
transform 1 0 30636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1666464484
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_349
timestamp 1666464484
transform 1 0 33212 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_355
timestamp 1666464484
transform 1 0 33764 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_372
timestamp 1666464484
transform 1 0 35328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_383
timestamp 1666464484
transform 1 0 36340 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1666464484
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_393
timestamp 1666464484
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_411
timestamp 1666464484
transform 1 0 38916 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_423
timestamp 1666464484
transform 1 0 40020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_435
timestamp 1666464484
transform 1 0 41124 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1666464484
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1666464484
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1666464484
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1666464484
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1666464484
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1666464484
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666464484
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1666464484
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1666464484
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1666464484
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1666464484
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1666464484
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1666464484
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1666464484
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1666464484
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1666464484
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_597
timestamp 1666464484
transform 1 0 56028 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1666464484
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1666464484
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_617
timestamp 1666464484
transform 1 0 57868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_622
timestamp 1666464484
transform 1 0 58328 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1666464484
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1666464484
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1666464484
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1666464484
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_121
timestamp 1666464484
transform 1 0 12236 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1666464484
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1666464484
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_177
timestamp 1666464484
transform 1 0 17388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 1666464484
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1666464484
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_228
timestamp 1666464484
transform 1 0 22080 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_239
timestamp 1666464484
transform 1 0 23092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_258
timestamp 1666464484
transform 1 0 24840 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_292
timestamp 1666464484
transform 1 0 27968 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_305
timestamp 1666464484
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1666464484
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_333
timestamp 1666464484
transform 1 0 31740 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_339
timestamp 1666464484
transform 1 0 32292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_347
timestamp 1666464484
transform 1 0 33028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1666464484
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1666464484
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_383
timestamp 1666464484
transform 1 0 36340 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_398
timestamp 1666464484
transform 1 0 37720 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1666464484
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1666464484
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1666464484
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1666464484
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1666464484
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1666464484
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1666464484
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1666464484
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1666464484
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1666464484
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1666464484
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1666464484
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1666464484
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1666464484
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1666464484
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1666464484
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1666464484
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1666464484
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1666464484
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1666464484
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1666464484
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_601
timestamp 1666464484
transform 1 0 56396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_605
timestamp 1666464484
transform 1 0 56764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_622
timestamp 1666464484
transform 1 0 58328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1666464484
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1666464484
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1666464484
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1666464484
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666464484
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1666464484
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1666464484
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp 1666464484
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_136
timestamp 1666464484
transform 1 0 13616 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_148
timestamp 1666464484
transform 1 0 14720 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_156
timestamp 1666464484
transform 1 0 15456 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 1666464484
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_175
timestamp 1666464484
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_186
timestamp 1666464484
transform 1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_197
timestamp 1666464484
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_207
timestamp 1666464484
transform 1 0 20148 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1666464484
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_233
timestamp 1666464484
transform 1 0 22540 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_241
timestamp 1666464484
transform 1 0 23276 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_248
timestamp 1666464484
transform 1 0 23920 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1666464484
transform 1 0 26680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_285
timestamp 1666464484
transform 1 0 27324 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_302
timestamp 1666464484
transform 1 0 28888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1666464484
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_349
timestamp 1666464484
transform 1 0 33212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_353
timestamp 1666464484
transform 1 0 33580 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_362
timestamp 1666464484
transform 1 0 34408 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_375
timestamp 1666464484
transform 1 0 35604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_387
timestamp 1666464484
transform 1 0 36708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1666464484
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_393
timestamp 1666464484
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_401
timestamp 1666464484
transform 1 0 37996 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_409
timestamp 1666464484
transform 1 0 38732 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_421
timestamp 1666464484
transform 1 0 39836 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_433
timestamp 1666464484
transform 1 0 40940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_445
timestamp 1666464484
transform 1 0 42044 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1666464484
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1666464484
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1666464484
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1666464484
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1666464484
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1666464484
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1666464484
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1666464484
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1666464484
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1666464484
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1666464484
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1666464484
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1666464484
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1666464484
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1666464484
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_597
timestamp 1666464484
transform 1 0 56028 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_605
timestamp 1666464484
transform 1 0 56764 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_614
timestamp 1666464484
transform 1 0 57592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1666464484
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_11
timestamp 1666464484
transform 1 0 2116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1666464484
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1666464484
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1666464484
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1666464484
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_121
timestamp 1666464484
transform 1 0 12236 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_129
timestamp 1666464484
transform 1 0 12972 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1666464484
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_153
timestamp 1666464484
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_164
timestamp 1666464484
transform 1 0 16192 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1666464484
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_203
timestamp 1666464484
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_213
timestamp 1666464484
transform 1 0 20700 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1666464484
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_264
timestamp 1666464484
transform 1 0 25392 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_270
timestamp 1666464484
transform 1 0 25944 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_297
timestamp 1666464484
transform 1 0 28428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp 1666464484
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_320
timestamp 1666464484
transform 1 0 30544 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_327
timestamp 1666464484
transform 1 0 31188 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_339
timestamp 1666464484
transform 1 0 32292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_351
timestamp 1666464484
transform 1 0 33396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666464484
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1666464484
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1666464484
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1666464484
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1666464484
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1666464484
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1666464484
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1666464484
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1666464484
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1666464484
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1666464484
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1666464484
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1666464484
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1666464484
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1666464484
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1666464484
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1666464484
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1666464484
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1666464484
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1666464484
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1666464484
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1666464484
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1666464484
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1666464484
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1666464484
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1666464484
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_601
timestamp 1666464484
transform 1 0 56396 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_613
timestamp 1666464484
transform 1 0 57500 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_623
timestamp 1666464484
transform 1 0 58420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_11
timestamp 1666464484
transform 1 0 2116 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_23
timestamp 1666464484
transform 1 0 3220 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_35
timestamp 1666464484
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1666464484
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1666464484
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1666464484
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1666464484
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_145
timestamp 1666464484
transform 1 0 14444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1666464484
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_177
timestamp 1666464484
transform 1 0 17388 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_204
timestamp 1666464484
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_208
timestamp 1666464484
transform 1 0 20240 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1666464484
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_235
timestamp 1666464484
transform 1 0 22724 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_241
timestamp 1666464484
transform 1 0 23276 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_268
timestamp 1666464484
transform 1 0 25760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1666464484
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_286
timestamp 1666464484
transform 1 0 27416 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_292
timestamp 1666464484
transform 1 0 27968 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_319
timestamp 1666464484
transform 1 0 30452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1666464484
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_349
timestamp 1666464484
transform 1 0 33212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_353
timestamp 1666464484
transform 1 0 33580 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_362
timestamp 1666464484
transform 1 0 34408 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_374
timestamp 1666464484
transform 1 0 35512 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_386
timestamp 1666464484
transform 1 0 36616 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1666464484
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1666464484
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1666464484
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1666464484
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1666464484
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1666464484
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1666464484
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1666464484
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1666464484
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1666464484
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1666464484
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1666464484
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1666464484
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1666464484
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_545
timestamp 1666464484
transform 1 0 51244 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_557
timestamp 1666464484
transform 1 0 52348 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1666464484
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1666464484
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1666464484
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_597
timestamp 1666464484
transform 1 0 56028 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1666464484
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1666464484
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_617
timestamp 1666464484
transform 1 0 57868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_622
timestamp 1666464484
transform 1 0 58328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_11
timestamp 1666464484
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1666464484
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1666464484
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1666464484
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1666464484
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1666464484
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_164
timestamp 1666464484
transform 1 0 16192 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1666464484
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_209
timestamp 1666464484
transform 1 0 20332 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_243
timestamp 1666464484
transform 1 0 23460 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1666464484
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_281
timestamp 1666464484
transform 1 0 26956 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1666464484
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666464484
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_327
timestamp 1666464484
transform 1 0 31188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_339
timestamp 1666464484
transform 1 0 32292 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1666464484
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1666464484
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1666464484
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1666464484
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1666464484
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1666464484
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1666464484
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1666464484
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1666464484
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1666464484
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1666464484
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1666464484
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1666464484
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1666464484
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1666464484
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1666464484
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1666464484
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1666464484
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1666464484
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1666464484
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1666464484
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1666464484
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1666464484
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1666464484
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1666464484
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1666464484
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_601
timestamp 1666464484
transform 1 0 56396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_605
timestamp 1666464484
transform 1 0 56764 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_622
timestamp 1666464484
transform 1 0 58328 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1666464484
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1666464484
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1666464484
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1666464484
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1666464484
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1666464484
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_190
timestamp 1666464484
transform 1 0 18584 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1666464484
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_244
timestamp 1666464484
transform 1 0 23552 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_248
timestamp 1666464484
transform 1 0 23920 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_275
timestamp 1666464484
transform 1 0 26404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_299
timestamp 1666464484
transform 1 0 28612 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_312
timestamp 1666464484
transform 1 0 29808 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_318
timestamp 1666464484
transform 1 0 30360 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_331
timestamp 1666464484
transform 1 0 31556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1666464484
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_344
timestamp 1666464484
transform 1 0 32752 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_352
timestamp 1666464484
transform 1 0 33488 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_360
timestamp 1666464484
transform 1 0 34224 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_372
timestamp 1666464484
transform 1 0 35328 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_384
timestamp 1666464484
transform 1 0 36432 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1666464484
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_405
timestamp 1666464484
transform 1 0 38364 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1666464484
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1666464484
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1666464484
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1666464484
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1666464484
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1666464484
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1666464484
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1666464484
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1666464484
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1666464484
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1666464484
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1666464484
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1666464484
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1666464484
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1666464484
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1666464484
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1666464484
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1666464484
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_597
timestamp 1666464484
transform 1 0 56028 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_605
timestamp 1666464484
transform 1 0 56764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_614
timestamp 1666464484
transform 1 0 57592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1666464484
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_11
timestamp 1666464484
transform 1 0 2116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1666464484
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1666464484
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1666464484
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1666464484
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1666464484
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1666464484
transform 1 0 14812 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_158
timestamp 1666464484
transform 1 0 15640 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1666464484
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_220
timestamp 1666464484
transform 1 0 21344 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1666464484
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_262
timestamp 1666464484
transform 1 0 25208 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_270
timestamp 1666464484
transform 1 0 25944 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_298
timestamp 1666464484
transform 1 0 28520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1666464484
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_323
timestamp 1666464484
transform 1 0 30820 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_335
timestamp 1666464484
transform 1 0 31924 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_344
timestamp 1666464484
transform 1 0 32752 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_356
timestamp 1666464484
transform 1 0 33856 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1666464484
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1666464484
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1666464484
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1666464484
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1666464484
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1666464484
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1666464484
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1666464484
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1666464484
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1666464484
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1666464484
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1666464484
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1666464484
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1666464484
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1666464484
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1666464484
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1666464484
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1666464484
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1666464484
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1666464484
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1666464484
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1666464484
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1666464484
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1666464484
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1666464484
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1666464484
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_613
timestamp 1666464484
transform 1 0 57500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_623
timestamp 1666464484
transform 1 0 58420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_11
timestamp 1666464484
transform 1 0 2116 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_23
timestamp 1666464484
transform 1 0 3220 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_35
timestamp 1666464484
transform 1 0 4324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1666464484
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1666464484
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1666464484
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1666464484
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_143
timestamp 1666464484
transform 1 0 14260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1666464484
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1666464484
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_180
timestamp 1666464484
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_190
timestamp 1666464484
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_201
timestamp 1666464484
transform 1 0 19596 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1666464484
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_231
timestamp 1666464484
transform 1 0 22356 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_248
timestamp 1666464484
transform 1 0 23920 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1666464484
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_309
timestamp 1666464484
transform 1 0 29532 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1666464484
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_361
timestamp 1666464484
transform 1 0 34316 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_381
timestamp 1666464484
transform 1 0 36156 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_389
timestamp 1666464484
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1666464484
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1666464484
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1666464484
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1666464484
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1666464484
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1666464484
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1666464484
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1666464484
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1666464484
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1666464484
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1666464484
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1666464484
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1666464484
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1666464484
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1666464484
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1666464484
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1666464484
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1666464484
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1666464484
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1666464484
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1666464484
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1666464484
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1666464484
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1666464484
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1666464484
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_11
timestamp 1666464484
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1666464484
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1666464484
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1666464484
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1666464484
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1666464484
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_149
timestamp 1666464484
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_178
timestamp 1666464484
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_185
timestamp 1666464484
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1666464484
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_204
timestamp 1666464484
transform 1 0 19872 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_234
timestamp 1666464484
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1666464484
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_271
timestamp 1666464484
transform 1 0 26036 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_279
timestamp 1666464484
transform 1 0 26772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1666464484
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_337
timestamp 1666464484
transform 1 0 32108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_361
timestamp 1666464484
transform 1 0 34316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1666464484
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_376
timestamp 1666464484
transform 1 0 35696 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_388
timestamp 1666464484
transform 1 0 36800 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_400
timestamp 1666464484
transform 1 0 37904 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_412
timestamp 1666464484
transform 1 0 39008 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1666464484
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1666464484
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1666464484
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1666464484
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1666464484
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1666464484
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1666464484
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_489
timestamp 1666464484
transform 1 0 46092 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_517
timestamp 1666464484
transform 1 0 48668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_529
timestamp 1666464484
transform 1 0 49772 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1666464484
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1666464484
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1666464484
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1666464484
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1666464484
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1666464484
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1666464484
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_601
timestamp 1666464484
transform 1 0 56396 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_613
timestamp 1666464484
transform 1 0 57500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_623
timestamp 1666464484
transform 1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_11
timestamp 1666464484
transform 1 0 2116 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_23
timestamp 1666464484
transform 1 0 3220 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_35
timestamp 1666464484
transform 1 0 4324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1666464484
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1666464484
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1666464484
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1666464484
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1666464484
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1666464484
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1666464484
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_188
timestamp 1666464484
transform 1 0 18400 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_201
timestamp 1666464484
transform 1 0 19596 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_214
timestamp 1666464484
transform 1 0 20792 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1666464484
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_231
timestamp 1666464484
transform 1 0 22356 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_248
timestamp 1666464484
transform 1 0 23920 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1666464484
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_309
timestamp 1666464484
transform 1 0 29532 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1666464484
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1666464484
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_351
timestamp 1666464484
transform 1 0 33396 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_364
timestamp 1666464484
transform 1 0 34592 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_372
timestamp 1666464484
transform 1 0 35328 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1666464484
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1666464484
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1666464484
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_433
timestamp 1666464484
transform 1 0 40940 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_445
timestamp 1666464484
transform 1 0 42044 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1666464484
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1666464484
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1666464484
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1666464484
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1666464484
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1666464484
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1666464484
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1666464484
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1666464484
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1666464484
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1666464484
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1666464484
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1666464484
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1666464484
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1666464484
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_597
timestamp 1666464484
transform 1 0 56028 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_603
timestamp 1666464484
transform 1 0 56580 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_611
timestamp 1666464484
transform 1 0 57316 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1666464484
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_617
timestamp 1666464484
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1666464484
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1666464484
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1666464484
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_97
timestamp 1666464484
transform 1 0 10028 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_117
timestamp 1666464484
transform 1 0 11868 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_129
timestamp 1666464484
transform 1 0 12972 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1666464484
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1666464484
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_153
timestamp 1666464484
transform 1 0 15180 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_161
timestamp 1666464484
transform 1 0 15916 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1666464484
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_183
timestamp 1666464484
transform 1 0 17940 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1666464484
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_208
timestamp 1666464484
transform 1 0 20240 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_218
timestamp 1666464484
transform 1 0 21160 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1666464484
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_262
timestamp 1666464484
transform 1 0 25208 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_266
timestamp 1666464484
transform 1 0 25576 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_276
timestamp 1666464484
transform 1 0 26496 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1666464484
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_328
timestamp 1666464484
transform 1 0 31280 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_339
timestamp 1666464484
transform 1 0 32292 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_348
timestamp 1666464484
transform 1 0 33120 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1666464484
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1666464484
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_377
timestamp 1666464484
transform 1 0 35788 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_381
timestamp 1666464484
transform 1 0 36156 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_391
timestamp 1666464484
transform 1 0 37076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_403
timestamp 1666464484
transform 1 0 38180 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_411
timestamp 1666464484
transform 1 0 38916 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_418
timestamp 1666464484
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_421
timestamp 1666464484
transform 1 0 39836 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_431
timestamp 1666464484
transform 1 0 40756 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_443
timestamp 1666464484
transform 1 0 41860 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_455
timestamp 1666464484
transform 1 0 42964 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_467
timestamp 1666464484
transform 1 0 44068 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1666464484
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1666464484
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1666464484
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1666464484
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1666464484
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1666464484
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1666464484
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1666464484
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1666464484
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1666464484
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1666464484
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1666464484
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1666464484
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_589
timestamp 1666464484
transform 1 0 55292 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_602
timestamp 1666464484
transform 1 0 56488 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_622
timestamp 1666464484
transform 1 0 58328 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_11
timestamp 1666464484
transform 1 0 2116 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_23
timestamp 1666464484
transform 1 0 3220 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_35
timestamp 1666464484
transform 1 0 4324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1666464484
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1666464484
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1666464484
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1666464484
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_149
timestamp 1666464484
transform 1 0 14812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_157
timestamp 1666464484
transform 1 0 15548 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_184
timestamp 1666464484
transform 1 0 18032 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_190
timestamp 1666464484
transform 1 0 18584 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_200
timestamp 1666464484
transform 1 0 19504 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_212
timestamp 1666464484
transform 1 0 20608 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1666464484
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_232
timestamp 1666464484
transform 1 0 22448 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_262
timestamp 1666464484
transform 1 0 25208 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1666464484
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_303
timestamp 1666464484
transform 1 0 28980 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_319
timestamp 1666464484
transform 1 0 30452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1666464484
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1666464484
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_344
timestamp 1666464484
transform 1 0 32752 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_358
timestamp 1666464484
transform 1 0 34040 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_371
timestamp 1666464484
transform 1 0 35236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_383
timestamp 1666464484
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1666464484
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1666464484
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_405
timestamp 1666464484
transform 1 0 38364 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_411
timestamp 1666464484
transform 1 0 38916 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_417
timestamp 1666464484
transform 1 0 39468 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_427
timestamp 1666464484
transform 1 0 40388 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_439
timestamp 1666464484
transform 1 0 41492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1666464484
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1666464484
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1666464484
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1666464484
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1666464484
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1666464484
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1666464484
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1666464484
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1666464484
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1666464484
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1666464484
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1666464484
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1666464484
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1666464484
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1666464484
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1666464484
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_597
timestamp 1666464484
transform 1 0 56028 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_605
timestamp 1666464484
transform 1 0 56764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_614
timestamp 1666464484
transform 1 0 57592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_617
timestamp 1666464484
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_11
timestamp 1666464484
transform 1 0 2116 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1666464484
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1666464484
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1666464484
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1666464484
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1666464484
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_153
timestamp 1666464484
transform 1 0 15180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_157
timestamp 1666464484
transform 1 0 15548 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_161
timestamp 1666464484
transform 1 0 15916 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_172
timestamp 1666464484
transform 1 0 16928 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_185
timestamp 1666464484
transform 1 0 18124 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1666464484
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_229
timestamp 1666464484
transform 1 0 22172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1666464484
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_258
timestamp 1666464484
transform 1 0 24840 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_269
timestamp 1666464484
transform 1 0 25852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_299
timestamp 1666464484
transform 1 0 28612 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1666464484
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_319
timestamp 1666464484
transform 1 0 30452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_328
timestamp 1666464484
transform 1 0 31280 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_332
timestamp 1666464484
transform 1 0 31648 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_340
timestamp 1666464484
transform 1 0 32384 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_352
timestamp 1666464484
transform 1 0 33488 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_365
timestamp 1666464484
transform 1 0 34684 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_373
timestamp 1666464484
transform 1 0 35420 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_393
timestamp 1666464484
transform 1 0 37260 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_406
timestamp 1666464484
transform 1 0 38456 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 1666464484
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1666464484
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_433
timestamp 1666464484
transform 1 0 40940 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_441
timestamp 1666464484
transform 1 0 41676 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_450
timestamp 1666464484
transform 1 0 42504 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_462
timestamp 1666464484
transform 1 0 43608 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_474
timestamp 1666464484
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1666464484
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1666464484
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1666464484
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1666464484
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1666464484
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1666464484
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1666464484
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1666464484
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1666464484
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1666464484
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1666464484
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1666464484
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1666464484
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_601
timestamp 1666464484
transform 1 0 56396 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_613
timestamp 1666464484
transform 1 0 57500 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_623
timestamp 1666464484
transform 1 0 58420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_11
timestamp 1666464484
transform 1 0 2116 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_23
timestamp 1666464484
transform 1 0 3220 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_35
timestamp 1666464484
transform 1 0 4324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1666464484
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666464484
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1666464484
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_93
timestamp 1666464484
transform 1 0 9660 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_103
timestamp 1666464484
transform 1 0 10580 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1666464484
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_156
timestamp 1666464484
transform 1 0 15456 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1666464484
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1666464484
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_183
timestamp 1666464484
transform 1 0 17940 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_192
timestamp 1666464484
transform 1 0 18768 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1666464484
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_248
timestamp 1666464484
transform 1 0 23920 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_278
timestamp 1666464484
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_286
timestamp 1666464484
transform 1 0 27416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_306
timestamp 1666464484
transform 1 0 29256 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_314
timestamp 1666464484
transform 1 0 29992 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1666464484
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_345
timestamp 1666464484
transform 1 0 32844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_357
timestamp 1666464484
transform 1 0 33948 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_369
timestamp 1666464484
transform 1 0 35052 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_381
timestamp 1666464484
transform 1 0 36156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_389
timestamp 1666464484
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_393
timestamp 1666464484
transform 1 0 37260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_397
timestamp 1666464484
transform 1 0 37628 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_406
timestamp 1666464484
transform 1 0 38456 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_415
timestamp 1666464484
transform 1 0 39284 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_419
timestamp 1666464484
transform 1 0 39652 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1666464484
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_441
timestamp 1666464484
transform 1 0 41676 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_445
timestamp 1666464484
transform 1 0 42044 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_449
timestamp 1666464484
transform 1 0 42412 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_467
timestamp 1666464484
transform 1 0 44068 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_479
timestamp 1666464484
transform 1 0 45172 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_491
timestamp 1666464484
transform 1 0 46276 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1666464484
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1666464484
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1666464484
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1666464484
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1666464484
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1666464484
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1666464484
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1666464484
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1666464484
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1666464484
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_597
timestamp 1666464484
transform 1 0 56028 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_611
timestamp 1666464484
transform 1 0 57316 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1666464484
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_617
timestamp 1666464484
transform 1 0 57868 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_622
timestamp 1666464484
transform 1 0 58328 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_11
timestamp 1666464484
transform 1 0 2116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1666464484
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1666464484
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1666464484
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_97
timestamp 1666464484
transform 1 0 10028 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_112
timestamp 1666464484
transform 1 0 11408 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_124
timestamp 1666464484
transform 1 0 12512 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1666464484
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_153
timestamp 1666464484
transform 1 0 15180 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_161
timestamp 1666464484
transform 1 0 15916 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_167
timestamp 1666464484
transform 1 0 16468 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_179
timestamp 1666464484
transform 1 0 17572 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1666464484
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_220
timestamp 1666464484
transform 1 0 21344 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1666464484
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_258
timestamp 1666464484
transform 1 0 24840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_288
timestamp 1666464484
transform 1 0 27600 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_300
timestamp 1666464484
transform 1 0 28704 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_334
timestamp 1666464484
transform 1 0 31832 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_346
timestamp 1666464484
transform 1 0 32936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1666464484
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_365
timestamp 1666464484
transform 1 0 34684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_381
timestamp 1666464484
transform 1 0 36156 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_401
timestamp 1666464484
transform 1 0 37996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1666464484
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1666464484
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1666464484
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1666464484
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_445
timestamp 1666464484
transform 1 0 42044 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_453
timestamp 1666464484
transform 1 0 42780 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_458
timestamp 1666464484
transform 1 0 43240 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_462
timestamp 1666464484
transform 1 0 43608 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_472
timestamp 1666464484
transform 1 0 44528 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1666464484
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1666464484
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1666464484
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1666464484
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1666464484
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1666464484
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1666464484
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1666464484
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1666464484
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1666464484
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1666464484
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1666464484
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1666464484
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_601
timestamp 1666464484
transform 1 0 56396 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_605
timestamp 1666464484
transform 1 0 56764 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_623
timestamp 1666464484
transform 1 0 58420 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1666464484
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1666464484
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1666464484
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1666464484
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1666464484
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_149
timestamp 1666464484
transform 1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1666464484
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1666464484
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_192
timestamp 1666464484
transform 1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1666464484
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_248
timestamp 1666464484
transform 1 0 23920 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1666464484
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_290
timestamp 1666464484
transform 1 0 27784 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_304
timestamp 1666464484
transform 1 0 29072 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1666464484
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_365
timestamp 1666464484
transform 1 0 34684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_386
timestamp 1666464484
transform 1 0 36616 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1666464484
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_403
timestamp 1666464484
transform 1 0 38180 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_426
timestamp 1666464484
transform 1 0 40296 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_438
timestamp 1666464484
transform 1 0 41400 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1666464484
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1666464484
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_461
timestamp 1666464484
transform 1 0 43516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_465
timestamp 1666464484
transform 1 0 43884 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_482
timestamp 1666464484
transform 1 0 45448 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_494
timestamp 1666464484
transform 1 0 46552 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_502
timestamp 1666464484
transform 1 0 47288 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1666464484
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1666464484
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1666464484
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1666464484
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_558
timestamp 1666464484
transform 1 0 52440 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1666464484
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1666464484
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1666464484
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_597
timestamp 1666464484
transform 1 0 56028 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1666464484
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1666464484
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1666464484
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_11
timestamp 1666464484
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1666464484
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1666464484
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1666464484
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1666464484
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1666464484
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_153
timestamp 1666464484
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1666464484
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1666464484
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_229
timestamp 1666464484
transform 1 0 22172 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_233
timestamp 1666464484
transform 1 0 22540 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1666464484
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_259
timestamp 1666464484
transform 1 0 24932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_289
timestamp 1666464484
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_297
timestamp 1666464484
transform 1 0 28428 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1666464484
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_325
timestamp 1666464484
transform 1 0 31004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_329
timestamp 1666464484
transform 1 0 31372 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_356
timestamp 1666464484
transform 1 0 33856 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1666464484
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_393
timestamp 1666464484
transform 1 0 37260 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1666464484
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1666464484
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_429
timestamp 1666464484
transform 1 0 40572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_433
timestamp 1666464484
transform 1 0 40940 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_441
timestamp 1666464484
transform 1 0 41676 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_453
timestamp 1666464484
transform 1 0 42780 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_465
timestamp 1666464484
transform 1 0 43884 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_473
timestamp 1666464484
transform 1 0 44620 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_477
timestamp 1666464484
transform 1 0 44988 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_493
timestamp 1666464484
transform 1 0 46460 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_505
timestamp 1666464484
transform 1 0 47564 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_517
timestamp 1666464484
transform 1 0 48668 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_529
timestamp 1666464484
transform 1 0 49772 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1666464484
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_545
timestamp 1666464484
transform 1 0 51244 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_561
timestamp 1666464484
transform 1 0 52716 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_573
timestamp 1666464484
transform 1 0 53820 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_585
timestamp 1666464484
transform 1 0 54924 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1666464484
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_601
timestamp 1666464484
transform 1 0 56396 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_613
timestamp 1666464484
transform 1 0 57500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_623
timestamp 1666464484
transform 1 0 58420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_11
timestamp 1666464484
transform 1 0 2116 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_23
timestamp 1666464484
transform 1 0 3220 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_35
timestamp 1666464484
transform 1 0 4324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_47
timestamp 1666464484
transform 1 0 5428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1666464484
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1666464484
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1666464484
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_149
timestamp 1666464484
transform 1 0 14812 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_157
timestamp 1666464484
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1666464484
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_178
timestamp 1666464484
transform 1 0 17480 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_184
timestamp 1666464484
transform 1 0 18032 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1666464484
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1666464484
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_248
timestamp 1666464484
transform 1 0 23920 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1666464484
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_290
timestamp 1666464484
transform 1 0 27784 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_298
timestamp 1666464484
transform 1 0 28520 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_325
timestamp 1666464484
transform 1 0 31004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1666464484
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_365
timestamp 1666464484
transform 1 0 34684 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_373
timestamp 1666464484
transform 1 0 35420 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_384
timestamp 1666464484
transform 1 0 36432 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1666464484
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_401
timestamp 1666464484
transform 1 0 37996 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_409
timestamp 1666464484
transform 1 0 38732 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_416
timestamp 1666464484
transform 1 0 39376 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_424
timestamp 1666464484
transform 1 0 40112 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1666464484
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1666464484
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1666464484
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1666464484
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1666464484
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_473
timestamp 1666464484
transform 1 0 44620 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_488
timestamp 1666464484
transform 1 0 46000 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1666464484
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1666464484
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1666464484
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_536
timestamp 1666464484
transform 1 0 50416 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_548
timestamp 1666464484
transform 1 0 51520 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_561
timestamp 1666464484
transform 1 0 52716 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_580
timestamp 1666464484
transform 1 0 54464 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_592
timestamp 1666464484
transform 1 0 55568 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_604
timestamp 1666464484
transform 1 0 56672 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1666464484
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_11
timestamp 1666464484
transform 1 0 2116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 1666464484
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1666464484
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1666464484
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1666464484
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1666464484
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_164
timestamp 1666464484
transform 1 0 16192 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1666464484
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_216
timestamp 1666464484
transform 1 0 20976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1666464484
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_262
timestamp 1666464484
transform 1 0 25208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_292
timestamp 1666464484
transform 1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_302
timestamp 1666464484
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_314
timestamp 1666464484
transform 1 0 29992 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_344
timestamp 1666464484
transform 1 0 32752 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_359
timestamp 1666464484
transform 1 0 34132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1666464484
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1666464484
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_374
timestamp 1666464484
transform 1 0 35512 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_390
timestamp 1666464484
transform 1 0 36984 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_399
timestamp 1666464484
transform 1 0 37812 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_407
timestamp 1666464484
transform 1 0 38548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1666464484
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_421
timestamp 1666464484
transform 1 0 39836 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_435
timestamp 1666464484
transform 1 0 41124 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_439
timestamp 1666464484
transform 1 0 41492 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_460
timestamp 1666464484
transform 1 0 43424 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_472
timestamp 1666464484
transform 1 0 44528 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1666464484
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_489
timestamp 1666464484
transform 1 0 46092 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_517
timestamp 1666464484
transform 1 0 48668 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_529
timestamp 1666464484
transform 1 0 49772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_533
timestamp 1666464484
transform 1 0 50140 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_551
timestamp 1666464484
transform 1 0 51796 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_563
timestamp 1666464484
transform 1 0 52900 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_575
timestamp 1666464484
transform 1 0 54004 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1666464484
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_589
timestamp 1666464484
transform 1 0 55292 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_595
timestamp 1666464484
transform 1 0 55844 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_602
timestamp 1666464484
transform 1 0 56488 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_622
timestamp 1666464484
transform 1 0 58328 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_9
timestamp 1666464484
transform 1 0 1932 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_21
timestamp 1666464484
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_33
timestamp 1666464484
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1666464484
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1666464484
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1666464484
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1666464484
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1666464484
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_144
timestamp 1666464484
transform 1 0 14352 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_159
timestamp 1666464484
transform 1 0 15732 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1666464484
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_192
timestamp 1666464484
transform 1 0 18768 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1666464484
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_248
timestamp 1666464484
transform 1 0 23920 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1666464484
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_291
timestamp 1666464484
transform 1 0 27876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_325
timestamp 1666464484
transform 1 0 31004 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_334
timestamp 1666464484
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_356
timestamp 1666464484
transform 1 0 33856 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_369
timestamp 1666464484
transform 1 0 35052 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_381
timestamp 1666464484
transform 1 0 36156 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_390
timestamp 1666464484
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1666464484
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_404
timestamp 1666464484
transform 1 0 38272 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_416
timestamp 1666464484
transform 1 0 39376 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_424
timestamp 1666464484
transform 1 0 40112 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_444
timestamp 1666464484
transform 1 0 41952 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1666464484
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_461
timestamp 1666464484
transform 1 0 43516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_465
timestamp 1666464484
transform 1 0 43884 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_482
timestamp 1666464484
transform 1 0 45448 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_494
timestamp 1666464484
transform 1 0 46552 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_502
timestamp 1666464484
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1666464484
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1666464484
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_529
timestamp 1666464484
transform 1 0 49772 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_537
timestamp 1666464484
transform 1 0 50508 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_549
timestamp 1666464484
transform 1 0 51612 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_557
timestamp 1666464484
transform 1 0 52348 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1666464484
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1666464484
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1666464484
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_597
timestamp 1666464484
transform 1 0 56028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_604
timestamp 1666464484
transform 1 0 56672 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_614
timestamp 1666464484
transform 1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_617
timestamp 1666464484
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1666464484
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1666464484
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1666464484
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1666464484
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1666464484
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1666464484
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_152
timestamp 1666464484
transform 1 0 15088 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_164
timestamp 1666464484
transform 1 0 16192 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1666464484
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_215
timestamp 1666464484
transform 1 0 20884 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_223
timestamp 1666464484
transform 1 0 21620 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1666464484
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_271
timestamp 1666464484
transform 1 0 26036 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_279
timestamp 1666464484
transform 1 0 26772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1666464484
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_320
timestamp 1666464484
transform 1 0 30544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_324
timestamp 1666464484
transform 1 0 30912 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_351
timestamp 1666464484
transform 1 0 33396 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1666464484
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1666464484
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_386
timestamp 1666464484
transform 1 0 36616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_394
timestamp 1666464484
transform 1 0 37352 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_405
timestamp 1666464484
transform 1 0 38364 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_414
timestamp 1666464484
transform 1 0 39192 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1666464484
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_429
timestamp 1666464484
transform 1 0 40572 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_441
timestamp 1666464484
transform 1 0 41676 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_453
timestamp 1666464484
transform 1 0 42780 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_460
timestamp 1666464484
transform 1 0 43424 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_472
timestamp 1666464484
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_477
timestamp 1666464484
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_487
timestamp 1666464484
transform 1 0 45908 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_491
timestamp 1666464484
transform 1 0 46276 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_503
timestamp 1666464484
transform 1 0 47380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_511
timestamp 1666464484
transform 1 0 48116 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_520
timestamp 1666464484
transform 1 0 48944 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1666464484
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1666464484
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1666464484
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1666464484
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1666464484
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1666464484
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1666464484
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1666464484
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_613
timestamp 1666464484
transform 1 0 57500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_623
timestamp 1666464484
transform 1 0 58420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_11
timestamp 1666464484
transform 1 0 2116 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_23
timestamp 1666464484
transform 1 0 3220 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_35
timestamp 1666464484
transform 1 0 4324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_47
timestamp 1666464484
transform 1 0 5428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666464484
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1666464484
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1666464484
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1666464484
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1666464484
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_182
timestamp 1666464484
transform 1 0 17848 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_214
timestamp 1666464484
transform 1 0 20792 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1666464484
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_231
timestamp 1666464484
transform 1 0 22356 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_248
timestamp 1666464484
transform 1 0 23920 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1666464484
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_300
timestamp 1666464484
transform 1 0 28704 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1666464484
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_365
timestamp 1666464484
transform 1 0 34684 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_377
timestamp 1666464484
transform 1 0 35788 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_381
timestamp 1666464484
transform 1 0 36156 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1666464484
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1666464484
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_400
timestamp 1666464484
transform 1 0 37904 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_408
timestamp 1666464484
transform 1 0 38640 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_427
timestamp 1666464484
transform 1 0 40388 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_439
timestamp 1666464484
transform 1 0 41492 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1666464484
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1666464484
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_461
timestamp 1666464484
transform 1 0 43516 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_467
timestamp 1666464484
transform 1 0 44068 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_488
timestamp 1666464484
transform 1 0 46000 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_500
timestamp 1666464484
transform 1 0 47104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_505
timestamp 1666464484
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_524
timestamp 1666464484
transform 1 0 49312 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_536
timestamp 1666464484
transform 1 0 50416 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_548
timestamp 1666464484
transform 1 0 51520 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1666464484
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1666464484
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1666464484
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_597
timestamp 1666464484
transform 1 0 56028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_601
timestamp 1666464484
transform 1 0 56396 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_605
timestamp 1666464484
transform 1 0 56764 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_613
timestamp 1666464484
transform 1 0 57500 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_617
timestamp 1666464484
transform 1 0 57868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1666464484
transform 1 0 58420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_11
timestamp 1666464484
transform 1 0 2116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 1666464484
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1666464484
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1666464484
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1666464484
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1666464484
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_153
timestamp 1666464484
transform 1 0 15180 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_178
timestamp 1666464484
transform 1 0 17480 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_186
timestamp 1666464484
transform 1 0 18216 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1666464484
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_206
timestamp 1666464484
transform 1 0 20056 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_218
timestamp 1666464484
transform 1 0 21160 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1666464484
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_260
timestamp 1666464484
transform 1 0 25024 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1666464484
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_274
timestamp 1666464484
transform 1 0 26312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1666464484
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_319
timestamp 1666464484
transform 1 0 30452 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_351
timestamp 1666464484
transform 1 0 33396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1666464484
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_365
timestamp 1666464484
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_380
timestamp 1666464484
transform 1 0 36064 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_384
timestamp 1666464484
transform 1 0 36432 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_402
timestamp 1666464484
transform 1 0 38088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_414
timestamp 1666464484
transform 1 0 39192 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1666464484
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_431
timestamp 1666464484
transform 1 0 40756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_443
timestamp 1666464484
transform 1 0 41860 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_452
timestamp 1666464484
transform 1 0 42688 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_466
timestamp 1666464484
transform 1 0 43976 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_474
timestamp 1666464484
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1666464484
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1666464484
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_501
timestamp 1666464484
transform 1 0 47196 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_515
timestamp 1666464484
transform 1 0 48484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_527
timestamp 1666464484
transform 1 0 49588 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1666464484
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_533
timestamp 1666464484
transform 1 0 50140 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_542
timestamp 1666464484
transform 1 0 50968 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_554
timestamp 1666464484
transform 1 0 52072 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_566
timestamp 1666464484
transform 1 0 53176 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_570
timestamp 1666464484
transform 1 0 53544 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_580
timestamp 1666464484
transform 1 0 54464 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_589
timestamp 1666464484
transform 1 0 55292 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_595
timestamp 1666464484
transform 1 0 55844 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_602
timestamp 1666464484
transform 1 0 56488 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_622
timestamp 1666464484
transform 1 0 58328 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_11
timestamp 1666464484
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_23
timestamp 1666464484
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_35
timestamp 1666464484
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1666464484
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666464484
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1666464484
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1666464484
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_125
timestamp 1666464484
transform 1 0 12604 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_133
timestamp 1666464484
transform 1 0 13340 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_140
timestamp 1666464484
transform 1 0 13984 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_152
timestamp 1666464484
transform 1 0 15088 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_156
timestamp 1666464484
transform 1 0 15456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_162
timestamp 1666464484
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_181
timestamp 1666464484
transform 1 0 17756 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_199
timestamp 1666464484
transform 1 0 19412 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_216
timestamp 1666464484
transform 1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_236
timestamp 1666464484
transform 1 0 22816 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_240
timestamp 1666464484
transform 1 0 23184 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_244
timestamp 1666464484
transform 1 0 23552 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_274
timestamp 1666464484
transform 1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_292
timestamp 1666464484
transform 1 0 27968 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_322
timestamp 1666464484
transform 1 0 30728 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1666464484
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_348
timestamp 1666464484
transform 1 0 33120 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_371
timestamp 1666464484
transform 1 0 35236 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_383
timestamp 1666464484
transform 1 0 36340 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1666464484
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_393
timestamp 1666464484
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_401
timestamp 1666464484
transform 1 0 37996 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_408
timestamp 1666464484
transform 1 0 38640 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1666464484
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_441
timestamp 1666464484
transform 1 0 41676 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_446
timestamp 1666464484
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1666464484
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_467
timestamp 1666464484
transform 1 0 44068 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_474
timestamp 1666464484
transform 1 0 44712 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_486
timestamp 1666464484
transform 1 0 45816 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_498
timestamp 1666464484
transform 1 0 46920 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1666464484
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1666464484
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_529
timestamp 1666464484
transform 1 0 49772 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_551
timestamp 1666464484
transform 1 0 51796 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1666464484
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_561
timestamp 1666464484
transform 1 0 52716 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_568
timestamp 1666464484
transform 1 0 53360 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_589
timestamp 1666464484
transform 1 0 55292 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_597
timestamp 1666464484
transform 1 0 56028 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_614
timestamp 1666464484
transform 1 0 57592 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1666464484
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_11
timestamp 1666464484
transform 1 0 2116 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_23
timestamp 1666464484
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1666464484
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1666464484
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1666464484
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1666464484
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1666464484
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_165
timestamp 1666464484
transform 1 0 16284 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_185
timestamp 1666464484
transform 1 0 18124 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_193
timestamp 1666464484
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_216
timestamp 1666464484
transform 1 0 20976 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_226
timestamp 1666464484
transform 1 0 21896 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1666464484
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666464484
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1666464484
transform 1 0 26036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1666464484
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1666464484
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_313
timestamp 1666464484
transform 1 0 29900 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_331
timestamp 1666464484
transform 1 0 31556 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_352
timestamp 1666464484
transform 1 0 33488 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1666464484
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1666464484
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1666464484
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1666464484
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1666464484
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1666464484
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1666464484
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1666464484
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1666464484
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_457
timestamp 1666464484
transform 1 0 43148 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_474
timestamp 1666464484
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1666464484
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1666464484
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1666464484
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1666464484
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1666464484
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_533
timestamp 1666464484
transform 1 0 50140 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_540
timestamp 1666464484
transform 1 0 50784 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_546
timestamp 1666464484
transform 1 0 51336 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_555
timestamp 1666464484
transform 1 0 52164 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_576
timestamp 1666464484
transform 1 0 54096 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_585
timestamp 1666464484
transform 1 0 54924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_589
timestamp 1666464484
transform 1 0 55292 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_613
timestamp 1666464484
transform 1 0 57500 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_623
timestamp 1666464484
transform 1 0 58420 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1666464484
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1666464484
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1666464484
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1666464484
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1666464484
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1666464484
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_149
timestamp 1666464484
transform 1 0 14812 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_157
timestamp 1666464484
transform 1 0 15548 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_165
timestamp 1666464484
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1666464484
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_193
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_197
timestamp 1666464484
transform 1 0 19228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_202
timestamp 1666464484
transform 1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1666464484
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_229
timestamp 1666464484
transform 1 0 22172 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_235
timestamp 1666464484
transform 1 0 22724 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1666464484
transform 1 0 23460 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_270
timestamp 1666464484
transform 1 0 25944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_274
timestamp 1666464484
transform 1 0 26312 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1666464484
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_305
timestamp 1666464484
transform 1 0 29164 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_325
timestamp 1666464484
transform 1 0 31004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_334
timestamp 1666464484
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_347
timestamp 1666464484
transform 1 0 33028 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_351
timestamp 1666464484
transform 1 0 33396 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_363
timestamp 1666464484
transform 1 0 34500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_375
timestamp 1666464484
transform 1 0 35604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_387
timestamp 1666464484
transform 1 0 36708 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1666464484
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1666464484
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1666464484
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1666464484
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1666464484
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1666464484
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1666464484
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1666464484
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1666464484
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_473
timestamp 1666464484
transform 1 0 44620 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_489
timestamp 1666464484
transform 1 0 46092 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_501
timestamp 1666464484
transform 1 0 47196 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1666464484
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1666464484
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1666464484
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1666464484
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1666464484
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1666464484
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1666464484
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_573
timestamp 1666464484
transform 1 0 53820 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_586
timestamp 1666464484
transform 1 0 55016 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_590
timestamp 1666464484
transform 1 0 55384 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_598
timestamp 1666464484
transform 1 0 56120 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1666464484
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1666464484
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_617
timestamp 1666464484
transform 1 0 57868 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_623
timestamp 1666464484
transform 1 0 58420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_11
timestamp 1666464484
transform 1 0 2116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_20
timestamp 1666464484
transform 1 0 2944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1666464484
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1666464484
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666464484
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1666464484
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1666464484
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1666464484
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_153
timestamp 1666464484
transform 1 0 15180 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_161
timestamp 1666464484
transform 1 0 15916 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_171
timestamp 1666464484
transform 1 0 16836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_183
timestamp 1666464484
transform 1 0 17940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666464484
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_214
timestamp 1666464484
transform 1 0 20792 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_218
timestamp 1666464484
transform 1 0 21160 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_229
timestamp 1666464484
transform 1 0 22172 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_241
timestamp 1666464484
transform 1 0 23276 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1666464484
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_275
timestamp 1666464484
transform 1 0 26404 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_299
timestamp 1666464484
transform 1 0 28612 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1666464484
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_316
timestamp 1666464484
transform 1 0 30176 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_328
timestamp 1666464484
transform 1 0 31280 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_340
timestamp 1666464484
transform 1 0 32384 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_352
timestamp 1666464484
transform 1 0 33488 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1666464484
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1666464484
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1666464484
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1666464484
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1666464484
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1666464484
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1666464484
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1666464484
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1666464484
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1666464484
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1666464484
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1666464484
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1666464484
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1666464484
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1666464484
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1666464484
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1666464484
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1666464484
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1666464484
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1666464484
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1666464484
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1666464484
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1666464484
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1666464484
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_589
timestamp 1666464484
transform 1 0 55292 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_600
timestamp 1666464484
transform 1 0 56304 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_609
timestamp 1666464484
transform 1 0 57132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_623
timestamp 1666464484
transform 1 0 58420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_11
timestamp 1666464484
transform 1 0 2116 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_23
timestamp 1666464484
transform 1 0 3220 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_35
timestamp 1666464484
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1666464484
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666464484
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1666464484
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1666464484
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1666464484
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1666464484
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1666464484
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666464484
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1666464484
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_193
timestamp 1666464484
transform 1 0 18860 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_201
timestamp 1666464484
transform 1 0 19596 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_205
timestamp 1666464484
transform 1 0 19964 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_216
timestamp 1666464484
transform 1 0 20976 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1666464484
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_261
timestamp 1666464484
transform 1 0 25116 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_264
timestamp 1666464484
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1666464484
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666464484
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_298
timestamp 1666464484
transform 1 0 28520 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_311
timestamp 1666464484
transform 1 0 29716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_323
timestamp 1666464484
transform 1 0 30820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666464484
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1666464484
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1666464484
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1666464484
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1666464484
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666464484
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1666464484
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1666464484
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1666464484
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1666464484
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1666464484
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1666464484
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1666464484
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1666464484
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1666464484
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1666464484
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1666464484
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1666464484
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1666464484
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1666464484
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1666464484
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1666464484
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1666464484
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1666464484
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1666464484
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1666464484
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1666464484
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1666464484
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1666464484
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1666464484
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_617
timestamp 1666464484
transform 1 0 57868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_623
timestamp 1666464484
transform 1 0 58420 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_11
timestamp 1666464484
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_20
timestamp 1666464484
transform 1 0 2944 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1666464484
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1666464484
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1666464484
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1666464484
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1666464484
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666464484
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1666464484
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_177
timestamp 1666464484
transform 1 0 17388 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1666464484
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_210
timestamp 1666464484
transform 1 0 20424 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_222
timestamp 1666464484
transform 1 0 21528 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_234
timestamp 1666464484
transform 1 0 22632 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_246
timestamp 1666464484
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_261
timestamp 1666464484
transform 1 0 25116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_265
timestamp 1666464484
transform 1 0 25484 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_276
timestamp 1666464484
transform 1 0 26496 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_44_287
timestamp 1666464484
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1666464484
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1666464484
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1666464484
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1666464484
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1666464484
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1666464484
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1666464484
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1666464484
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1666464484
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1666464484
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1666464484
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1666464484
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1666464484
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1666464484
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1666464484
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1666464484
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1666464484
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1666464484
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1666464484
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1666464484
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1666464484
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1666464484
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1666464484
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1666464484
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1666464484
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1666464484
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1666464484
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1666464484
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1666464484
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1666464484
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1666464484
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1666464484
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1666464484
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_613
timestamp 1666464484
transform 1 0 57500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_623
timestamp 1666464484
transform 1 0 58420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_11
timestamp 1666464484
transform 1 0 2116 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_20
timestamp 1666464484
transform 1 0 2944 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_32
timestamp 1666464484
transform 1 0 4048 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_44
timestamp 1666464484
transform 1 0 5152 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1666464484
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1666464484
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1666464484
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666464484
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1666464484
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1666464484
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1666464484
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_181
timestamp 1666464484
transform 1 0 17756 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_195
timestamp 1666464484
transform 1 0 19044 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_212
timestamp 1666464484
transform 1 0 20608 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1666464484
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1666464484
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1666464484
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1666464484
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666464484
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1666464484
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1666464484
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1666464484
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1666464484
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1666464484
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1666464484
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1666464484
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1666464484
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1666464484
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1666464484
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1666464484
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1666464484
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1666464484
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1666464484
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1666464484
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1666464484
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1666464484
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1666464484
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1666464484
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1666464484
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1666464484
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666464484
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1666464484
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1666464484
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1666464484
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1666464484
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1666464484
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1666464484
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1666464484
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1666464484
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1666464484
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1666464484
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1666464484
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1666464484
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1666464484
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_9
timestamp 1666464484
transform 1 0 1932 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1666464484
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1666464484
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1666464484
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1666464484
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666464484
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1666464484
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1666464484
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1666464484
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1666464484
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1666464484
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_177
timestamp 1666464484
transform 1 0 17388 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1666464484
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1666464484
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1666464484
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1666464484
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1666464484
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666464484
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1666464484
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1666464484
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1666464484
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1666464484
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1666464484
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1666464484
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1666464484
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1666464484
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1666464484
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1666464484
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1666464484
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1666464484
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1666464484
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1666464484
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1666464484
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1666464484
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1666464484
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1666464484
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1666464484
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1666464484
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1666464484
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1666464484
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1666464484
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1666464484
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1666464484
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1666464484
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1666464484
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1666464484
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1666464484
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1666464484
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1666464484
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1666464484
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1666464484
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1666464484
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1666464484
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1666464484
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_613
timestamp 1666464484
transform 1 0 57500 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_623
timestamp 1666464484
transform 1 0 58420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_9
timestamp 1666464484
transform 1 0 1932 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_13
timestamp 1666464484
transform 1 0 2300 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_20
timestamp 1666464484
transform 1 0 2944 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1666464484
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1666464484
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1666464484
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1666464484
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1666464484
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1666464484
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666464484
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1666464484
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1666464484
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1666464484
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1666464484
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1666464484
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1666464484
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1666464484
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1666464484
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1666464484
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1666464484
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1666464484
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1666464484
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1666464484
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1666464484
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1666464484
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1666464484
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1666464484
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1666464484
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1666464484
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1666464484
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1666464484
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1666464484
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1666464484
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1666464484
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1666464484
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1666464484
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1666464484
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1666464484
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1666464484
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1666464484
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1666464484
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1666464484
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1666464484
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1666464484
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1666464484
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1666464484
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1666464484
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1666464484
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1666464484
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1666464484
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1666464484
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1666464484
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1666464484
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1666464484
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1666464484
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1666464484
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1666464484
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1666464484
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1666464484
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1666464484
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_11
timestamp 1666464484
transform 1 0 2116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_20
timestamp 1666464484
transform 1 0 2944 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1666464484
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1666464484
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1666464484
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1666464484
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1666464484
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1666464484
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1666464484
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1666464484
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1666464484
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666464484
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1666464484
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1666464484
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1666464484
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1666464484
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666464484
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1666464484
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1666464484
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1666464484
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1666464484
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666464484
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1666464484
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1666464484
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1666464484
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1666464484
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666464484
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1666464484
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1666464484
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1666464484
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1666464484
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1666464484
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1666464484
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1666464484
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1666464484
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1666464484
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1666464484
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1666464484
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1666464484
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1666464484
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1666464484
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1666464484
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1666464484
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1666464484
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1666464484
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1666464484
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1666464484
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1666464484
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1666464484
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1666464484
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1666464484
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1666464484
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1666464484
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_613
timestamp 1666464484
transform 1 0 57500 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_623
timestamp 1666464484
transform 1 0 58420 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_11
timestamp 1666464484
transform 1 0 2116 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_23
timestamp 1666464484
transform 1 0 3220 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_35
timestamp 1666464484
transform 1 0 4324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp 1666464484
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1666464484
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1666464484
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1666464484
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666464484
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1666464484
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1666464484
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1666464484
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1666464484
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_181
timestamp 1666464484
transform 1 0 17756 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_194
timestamp 1666464484
transform 1 0 18952 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_198
timestamp 1666464484
transform 1 0 19320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_203
timestamp 1666464484
transform 1 0 19780 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1666464484
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1666464484
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_237
timestamp 1666464484
transform 1 0 22908 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_247
timestamp 1666464484
transform 1 0 23828 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_254
timestamp 1666464484
transform 1 0 24472 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_266
timestamp 1666464484
transform 1 0 25576 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1666464484
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1666464484
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1666464484
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1666464484
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1666464484
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1666464484
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1666464484
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1666464484
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1666464484
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1666464484
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1666464484
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1666464484
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1666464484
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1666464484
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1666464484
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1666464484
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666464484
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1666464484
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1666464484
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1666464484
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1666464484
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1666464484
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1666464484
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1666464484
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1666464484
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1666464484
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1666464484
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1666464484
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1666464484
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1666464484
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1666464484
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1666464484
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1666464484
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1666464484
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1666464484
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1666464484
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_11
timestamp 1666464484
transform 1 0 2116 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_23
timestamp 1666464484
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1666464484
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1666464484
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1666464484
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1666464484
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1666464484
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1666464484
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666464484
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_158
timestamp 1666464484
transform 1 0 15640 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_170
timestamp 1666464484
transform 1 0 16744 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_182
timestamp 1666464484
transform 1 0 17848 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1666464484
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_218
timestamp 1666464484
transform 1 0 21160 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_228
timestamp 1666464484
transform 1 0 22080 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_240
timestamp 1666464484
transform 1 0 23184 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1666464484
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1666464484
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1666464484
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1666464484
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666464484
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1666464484
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1666464484
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1666464484
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1666464484
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666464484
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1666464484
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_374
timestamp 1666464484
transform 1 0 35512 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_386
timestamp 1666464484
transform 1 0 36616 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_398
timestamp 1666464484
transform 1 0 37720 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_410
timestamp 1666464484
transform 1 0 38824 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_418
timestamp 1666464484
transform 1 0 39560 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1666464484
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1666464484
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1666464484
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_466
timestamp 1666464484
transform 1 0 43976 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_474
timestamp 1666464484
transform 1 0 44712 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1666464484
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1666464484
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1666464484
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1666464484
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1666464484
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1666464484
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1666464484
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1666464484
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1666464484
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1666464484
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1666464484
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1666464484
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1666464484
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_601
timestamp 1666464484
transform 1 0 56396 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 1666464484
transform 1 0 57500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_623
timestamp 1666464484
transform 1 0 58420 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1666464484
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1666464484
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1666464484
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1666464484
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1666464484
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1666464484
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1666464484
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1666464484
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666464484
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_177
timestamp 1666464484
transform 1 0 17388 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_193
timestamp 1666464484
transform 1 0 18860 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_203
timestamp 1666464484
transform 1 0 19780 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1666464484
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_234
timestamp 1666464484
transform 1 0 22632 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_246
timestamp 1666464484
transform 1 0 23736 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_258
timestamp 1666464484
transform 1 0 24840 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_270
timestamp 1666464484
transform 1 0 25944 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1666464484
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1666464484
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1666464484
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1666464484
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1666464484
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666464484
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1666464484
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1666464484
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1666464484
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1666464484
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1666464484
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1666464484
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_402
timestamp 1666464484
transform 1 0 38088 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_414
timestamp 1666464484
transform 1 0 39192 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_426
timestamp 1666464484
transform 1 0 40296 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_438
timestamp 1666464484
transform 1 0 41400 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_446
timestamp 1666464484
transform 1 0 42136 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1666464484
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1666464484
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1666464484
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1666464484
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1666464484
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1666464484
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1666464484
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1666464484
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1666464484
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1666464484
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1666464484
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1666464484
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1666464484
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1666464484
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1666464484
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1666464484
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1666464484
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1666464484
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1666464484
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1666464484
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1666464484
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1666464484
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1666464484
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1666464484
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1666464484
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1666464484
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1666464484
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666464484
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1666464484
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1666464484
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_190
timestamp 1666464484
transform 1 0 18584 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_216
timestamp 1666464484
transform 1 0 20976 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_234
timestamp 1666464484
transform 1 0 22632 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1666464484
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666464484
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_262
timestamp 1666464484
transform 1 0 25208 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_274
timestamp 1666464484
transform 1 0 26312 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_286
timestamp 1666464484
transform 1 0 27416 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_298
timestamp 1666464484
transform 1 0 28520 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1666464484
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_325
timestamp 1666464484
transform 1 0 31004 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_337
timestamp 1666464484
transform 1 0 32108 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_349
timestamp 1666464484
transform 1 0 33212 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1666464484
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1666464484
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_385
timestamp 1666464484
transform 1 0 36524 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_397
timestamp 1666464484
transform 1 0 37628 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_408
timestamp 1666464484
transform 1 0 38640 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1666464484
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1666464484
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1666464484
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1666464484
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1666464484
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1666464484
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1666464484
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1666464484
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1666464484
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1666464484
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1666464484
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1666464484
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1666464484
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1666464484
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1666464484
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1666464484
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1666464484
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1666464484
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1666464484
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1666464484
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_613
timestamp 1666464484
transform 1 0 57500 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_623
timestamp 1666464484
transform 1 0 58420 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_9
timestamp 1666464484
transform 1 0 1932 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_21
timestamp 1666464484
transform 1 0 3036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1666464484
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1666464484
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1666464484
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1666464484
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1666464484
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1666464484
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666464484
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1666464484
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1666464484
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1666464484
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1666464484
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666464484
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_181
timestamp 1666464484
transform 1 0 17756 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_203
timestamp 1666464484
transform 1 0 19780 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1666464484
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_244
timestamp 1666464484
transform 1 0 23552 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_256
timestamp 1666464484
transform 1 0 24656 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_265
timestamp 1666464484
transform 1 0 25484 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1666464484
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1666464484
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1666464484
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1666464484
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1666464484
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1666464484
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_349
timestamp 1666464484
transform 1 0 33212 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_364
timestamp 1666464484
transform 1 0 34592 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_376
timestamp 1666464484
transform 1 0 35696 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_382
timestamp 1666464484
transform 1 0 36248 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1666464484
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1666464484
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1666464484
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1666464484
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1666464484
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1666464484
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1666464484
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1666464484
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1666464484
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1666464484
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1666464484
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1666464484
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1666464484
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1666464484
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1666464484
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1666464484
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1666464484
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1666464484
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1666464484
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1666464484
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1666464484
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1666464484
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1666464484
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1666464484
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1666464484
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1666464484
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_9
timestamp 1666464484
transform 1 0 1932 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1666464484
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1666464484
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1666464484
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666464484
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1666464484
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1666464484
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1666464484
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1666464484
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1666464484
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_165
timestamp 1666464484
transform 1 0 16284 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_173
timestamp 1666464484
transform 1 0 17020 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1666464484
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_212
timestamp 1666464484
transform 1 0 20608 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_216
timestamp 1666464484
transform 1 0 20976 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_229
timestamp 1666464484
transform 1 0 22172 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_237
timestamp 1666464484
transform 1 0 22908 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1666464484
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666464484
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_259
timestamp 1666464484
transform 1 0 24932 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_269
timestamp 1666464484
transform 1 0 25852 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_281
timestamp 1666464484
transform 1 0 26956 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_293
timestamp 1666464484
transform 1 0 28060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_305
timestamp 1666464484
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1666464484
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1666464484
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1666464484
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666464484
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1666464484
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1666464484
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1666464484
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1666464484
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1666464484
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1666464484
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1666464484
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1666464484
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_445
timestamp 1666464484
transform 1 0 42044 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_455
timestamp 1666464484
transform 1 0 42964 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_463
timestamp 1666464484
transform 1 0 43700 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_474
timestamp 1666464484
transform 1 0 44712 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1666464484
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1666464484
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1666464484
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1666464484
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1666464484
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1666464484
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1666464484
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1666464484
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1666464484
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1666464484
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1666464484
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1666464484
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1666464484
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1666464484
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_613
timestamp 1666464484
transform 1 0 57500 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_623
timestamp 1666464484
transform 1 0 58420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_9
timestamp 1666464484
transform 1 0 1932 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_21
timestamp 1666464484
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_33
timestamp 1666464484
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1666464484
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1666464484
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1666464484
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1666464484
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1666464484
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1666464484
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_181
timestamp 1666464484
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_198
timestamp 1666464484
transform 1 0 19320 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_213
timestamp 1666464484
transform 1 0 20700 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_221
timestamp 1666464484
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_235
timestamp 1666464484
transform 1 0 22724 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_247
timestamp 1666464484
transform 1 0 23828 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_259
timestamp 1666464484
transform 1 0 24932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_263
timestamp 1666464484
transform 1 0 25300 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_271
timestamp 1666464484
transform 1 0 26036 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1666464484
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1666464484
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1666464484
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1666464484
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1666464484
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1666464484
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_357
timestamp 1666464484
transform 1 0 33948 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_369
timestamp 1666464484
transform 1 0 35052 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_381
timestamp 1666464484
transform 1 0 36156 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_389
timestamp 1666464484
transform 1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1666464484
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1666464484
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1666464484
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1666464484
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1666464484
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1666464484
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1666464484
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1666464484
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_473
timestamp 1666464484
transform 1 0 44620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_482
timestamp 1666464484
transform 1 0 45448 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_494
timestamp 1666464484
transform 1 0 46552 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_502
timestamp 1666464484
transform 1 0 47288 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1666464484
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1666464484
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1666464484
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1666464484
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1666464484
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1666464484
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1666464484
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1666464484
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1666464484
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1666464484
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1666464484
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1666464484
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1666464484
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1666464484
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666464484
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1666464484
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1666464484
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1666464484
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1666464484
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1666464484
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1666464484
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666464484
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1666464484
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_165
timestamp 1666464484
transform 1 0 16284 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_173
timestamp 1666464484
transform 1 0 17020 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1666464484
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666464484
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_209
timestamp 1666464484
transform 1 0 20332 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_215
timestamp 1666464484
transform 1 0 20884 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1666464484
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1666464484
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666464484
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_274
timestamp 1666464484
transform 1 0 26312 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_287
timestamp 1666464484
transform 1 0 27508 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_299
timestamp 1666464484
transform 1 0 28612 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1666464484
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1666464484
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1666464484
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_352
timestamp 1666464484
transform 1 0 33488 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1666464484
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1666464484
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1666464484
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1666464484
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1666464484
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1666464484
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1666464484
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1666464484
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1666464484
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_445
timestamp 1666464484
transform 1 0 42044 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_453
timestamp 1666464484
transform 1 0 42780 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_463
timestamp 1666464484
transform 1 0 43700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1666464484
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1666464484
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1666464484
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1666464484
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1666464484
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1666464484
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1666464484
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1666464484
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1666464484
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1666464484
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1666464484
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1666464484
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1666464484
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1666464484
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_601
timestamp 1666464484
transform 1 0 56396 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_613
timestamp 1666464484
transform 1 0 57500 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_623
timestamp 1666464484
transform 1 0 58420 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_9
timestamp 1666464484
transform 1 0 1932 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1666464484
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1666464484
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1666464484
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1666464484
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1666464484
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1666464484
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1666464484
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1666464484
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666464484
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1666464484
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1666464484
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1666464484
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_177
timestamp 1666464484
transform 1 0 17388 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_191
timestamp 1666464484
transform 1 0 18676 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_203
timestamp 1666464484
transform 1 0 19780 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_212
timestamp 1666464484
transform 1 0 20608 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_237
timestamp 1666464484
transform 1 0 22908 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_243
timestamp 1666464484
transform 1 0 23460 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_256
timestamp 1666464484
transform 1 0 24656 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_269
timestamp 1666464484
transform 1 0 25852 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 1666464484
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_300
timestamp 1666464484
transform 1 0 28704 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_313
timestamp 1666464484
transform 1 0 29900 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_325
timestamp 1666464484
transform 1 0 31004 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1666464484
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_343
timestamp 1666464484
transform 1 0 32660 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_351
timestamp 1666464484
transform 1 0 33396 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_363
timestamp 1666464484
transform 1 0 34500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_375
timestamp 1666464484
transform 1 0 35604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_387
timestamp 1666464484
transform 1 0 36708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1666464484
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1666464484
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1666464484
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1666464484
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1666464484
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1666464484
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1666464484
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1666464484
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1666464484
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1666464484
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1666464484
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1666464484
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666464484
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1666464484
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1666464484
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1666464484
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1666464484
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1666464484
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1666464484
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1666464484
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1666464484
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1666464484
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1666464484
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1666464484
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1666464484
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_617
timestamp 1666464484
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_9
timestamp 1666464484
transform 1 0 1932 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_21
timestamp 1666464484
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666464484
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1666464484
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1666464484
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1666464484
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1666464484
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1666464484
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666464484
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1666464484
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1666464484
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1666464484
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1666464484
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1666464484
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666464484
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1666464484
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1666464484
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_165
timestamp 1666464484
transform 1 0 16284 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_181
timestamp 1666464484
transform 1 0 17756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 1666464484
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_197
timestamp 1666464484
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_212
timestamp 1666464484
transform 1 0 20608 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_224
timestamp 1666464484
transform 1 0 21712 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_228
timestamp 1666464484
transform 1 0 22080 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_234
timestamp 1666464484
transform 1 0 22632 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_247
timestamp 1666464484
transform 1 0 23828 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1666464484
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1666464484
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_263
timestamp 1666464484
transform 1 0 25300 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_275
timestamp 1666464484
transform 1 0 26404 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_287
timestamp 1666464484
transform 1 0 27508 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_299
timestamp 1666464484
transform 1 0 28612 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1666464484
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1666464484
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1666464484
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1666464484
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1666464484
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1666464484
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1666464484
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1666464484
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1666464484
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1666464484
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1666464484
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1666464484
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1666464484
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_421
timestamp 1666464484
transform 1 0 39836 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_433
timestamp 1666464484
transform 1 0 40940 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_441
timestamp 1666464484
transform 1 0 41676 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_453
timestamp 1666464484
transform 1 0 42780 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_465
timestamp 1666464484
transform 1 0 43884 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_473
timestamp 1666464484
transform 1 0 44620 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1666464484
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1666464484
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1666464484
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1666464484
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1666464484
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1666464484
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1666464484
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1666464484
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1666464484
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1666464484
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1666464484
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1666464484
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1666464484
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1666464484
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_613
timestamp 1666464484
transform 1 0 57500 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_623
timestamp 1666464484
transform 1 0 58420 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_9
timestamp 1666464484
transform 1 0 1932 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_21
timestamp 1666464484
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_33
timestamp 1666464484
transform 1 0 4140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_45
timestamp 1666464484
transform 1 0 5244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1666464484
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1666464484
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1666464484
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1666464484
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1666464484
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1666464484
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666464484
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1666464484
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1666464484
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1666464484
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1666464484
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1666464484
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666464484
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1666464484
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1666464484
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1666464484
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1666464484
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1666464484
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1666464484
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_225
timestamp 1666464484
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_236
timestamp 1666464484
transform 1 0 22816 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1666464484
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1666464484
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1666464484
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1666464484
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1666464484
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1666464484
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1666464484
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1666464484
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1666464484
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1666464484
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1666464484
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1666464484
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1666464484
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1666464484
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1666464484
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1666464484
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1666464484
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1666464484
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1666464484
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1666464484
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1666464484
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1666464484
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1666464484
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1666464484
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1666464484
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1666464484
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1666464484
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1666464484
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1666464484
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1666464484
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1666464484
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1666464484
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1666464484
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1666464484
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1666464484
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1666464484
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1666464484
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1666464484
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1666464484
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1666464484
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_9
timestamp 1666464484
transform 1 0 1932 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_18
timestamp 1666464484
transform 1 0 2760 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1666464484
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1666464484
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1666464484
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1666464484
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1666464484
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1666464484
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666464484
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1666464484
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1666464484
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1666464484
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1666464484
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1666464484
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666464484
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1666464484
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_153
timestamp 1666464484
transform 1 0 15180 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_176
timestamp 1666464484
transform 1 0 17296 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_188
timestamp 1666464484
transform 1 0 18400 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1666464484
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_209
timestamp 1666464484
transform 1 0 20332 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_213
timestamp 1666464484
transform 1 0 20700 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_216
timestamp 1666464484
transform 1 0 20976 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_224
timestamp 1666464484
transform 1 0 21712 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_237
timestamp 1666464484
transform 1 0 22908 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_241
timestamp 1666464484
transform 1 0 23276 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_244
timestamp 1666464484
transform 1 0 23552 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1666464484
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1666464484
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_257
timestamp 1666464484
transform 1 0 24748 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1666464484
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1666464484
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1666464484
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1666464484
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1666464484
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1666464484
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1666464484
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1666464484
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1666464484
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1666464484
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1666464484
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1666464484
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1666464484
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1666464484
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1666464484
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1666464484
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1666464484
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1666464484
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1666464484
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1666464484
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1666464484
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1666464484
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1666464484
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1666464484
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1666464484
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1666464484
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1666464484
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1666464484
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1666464484
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1666464484
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1666464484
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1666464484
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1666464484
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1666464484
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1666464484
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1666464484
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1666464484
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1666464484
transform 1 0 57500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_623
timestamp 1666464484
transform 1 0 58420 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_9
timestamp 1666464484
transform 1 0 1932 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_18
timestamp 1666464484
transform 1 0 2760 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_30
timestamp 1666464484
transform 1 0 3864 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_42
timestamp 1666464484
transform 1 0 4968 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1666464484
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1666464484
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1666464484
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1666464484
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1666464484
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1666464484
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666464484
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1666464484
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1666464484
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1666464484
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1666464484
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1666464484
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666464484
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1666464484
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_181
timestamp 1666464484
transform 1 0 17756 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_185
timestamp 1666464484
transform 1 0 18124 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1666464484
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_205
timestamp 1666464484
transform 1 0 19964 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_209
timestamp 1666464484
transform 1 0 20332 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_212
timestamp 1666464484
transform 1 0 20608 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1666464484
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1666464484
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_243
timestamp 1666464484
transform 1 0 23460 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_251
timestamp 1666464484
transform 1 0 24196 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_266
timestamp 1666464484
transform 1 0 25576 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1666464484
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1666464484
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1666464484
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1666464484
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1666464484
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1666464484
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1666464484
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1666464484
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1666464484
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1666464484
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1666464484
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1666464484
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1666464484
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1666464484
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1666464484
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1666464484
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1666464484
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1666464484
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1666464484
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1666464484
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1666464484
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1666464484
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1666464484
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1666464484
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1666464484
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1666464484
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1666464484
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1666464484
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1666464484
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1666464484
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1666464484
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1666464484
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1666464484
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1666464484
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1666464484
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1666464484
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1666464484
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1666464484
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_9
timestamp 1666464484
transform 1 0 1932 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1666464484
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666464484
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1666464484
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1666464484
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1666464484
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1666464484
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1666464484
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666464484
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1666464484
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1666464484
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1666464484
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1666464484
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1666464484
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666464484
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1666464484
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1666464484
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1666464484
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_177
timestamp 1666464484
transform 1 0 17388 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1666464484
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1666464484
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_209
timestamp 1666464484
transform 1 0 20332 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_217
timestamp 1666464484
transform 1 0 21068 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_227
timestamp 1666464484
transform 1 0 21988 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_240
timestamp 1666464484
transform 1 0 23184 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1666464484
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_262
timestamp 1666464484
transform 1 0 25208 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_274
timestamp 1666464484
transform 1 0 26312 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_286
timestamp 1666464484
transform 1 0 27416 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_298
timestamp 1666464484
transform 1 0 28520 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1666464484
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1666464484
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1666464484
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1666464484
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1666464484
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1666464484
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1666464484
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1666464484
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1666464484
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1666464484
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1666464484
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1666464484
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1666464484
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1666464484
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1666464484
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1666464484
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1666464484
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1666464484
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1666464484
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1666464484
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1666464484
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1666464484
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1666464484
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1666464484
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1666464484
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1666464484
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1666464484
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1666464484
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1666464484
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1666464484
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1666464484
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1666464484
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1666464484
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 1666464484
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_623
timestamp 1666464484
transform 1 0 58420 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_9
timestamp 1666464484
transform 1 0 1932 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_21
timestamp 1666464484
transform 1 0 3036 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_33
timestamp 1666464484
transform 1 0 4140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_45
timestamp 1666464484
transform 1 0 5244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_53
timestamp 1666464484
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1666464484
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1666464484
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1666464484
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1666464484
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1666464484
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666464484
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1666464484
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1666464484
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1666464484
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1666464484
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1666464484
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1666464484
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1666464484
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1666464484
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1666464484
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_205
timestamp 1666464484
transform 1 0 19964 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_211
timestamp 1666464484
transform 1 0 20516 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_221
timestamp 1666464484
transform 1 0 21436 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1666464484
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_244
timestamp 1666464484
transform 1 0 23552 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_256
timestamp 1666464484
transform 1 0 24656 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_268
timestamp 1666464484
transform 1 0 25760 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1666464484
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1666464484
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1666464484
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1666464484
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1666464484
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1666464484
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1666464484
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1666464484
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1666464484
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1666464484
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1666464484
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1666464484
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1666464484
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1666464484
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1666464484
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1666464484
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1666464484
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1666464484
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1666464484
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1666464484
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_473
timestamp 1666464484
transform 1 0 44620 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_487
timestamp 1666464484
transform 1 0 45908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_499
timestamp 1666464484
transform 1 0 47012 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1666464484
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1666464484
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1666464484
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1666464484
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1666464484
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1666464484
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1666464484
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1666464484
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1666464484
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1666464484
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1666464484
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1666464484
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1666464484
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1666464484
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_9
timestamp 1666464484
transform 1 0 1932 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_17
timestamp 1666464484
transform 1 0 2668 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_25
timestamp 1666464484
transform 1 0 3404 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1666464484
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1666464484
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1666464484
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1666464484
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1666464484
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1666464484
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1666464484
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1666464484
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1666464484
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1666464484
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1666464484
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1666464484
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1666464484
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1666464484
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1666464484
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1666464484
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1666464484
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1666464484
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_197
timestamp 1666464484
transform 1 0 19228 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_206
timestamp 1666464484
transform 1 0 20056 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_222
timestamp 1666464484
transform 1 0 21528 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1666464484
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1666464484
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1666464484
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1666464484
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1666464484
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1666464484
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1666464484
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1666464484
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1666464484
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1666464484
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1666464484
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1666464484
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1666464484
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1666464484
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1666464484
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1666464484
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1666464484
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1666464484
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1666464484
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1666464484
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1666464484
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1666464484
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1666464484
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1666464484
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1666464484
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1666464484
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1666464484
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_477
timestamp 1666464484
transform 1 0 44988 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_486
timestamp 1666464484
transform 1 0 45816 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_497
timestamp 1666464484
transform 1 0 46828 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_509
timestamp 1666464484
transform 1 0 47932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_521
timestamp 1666464484
transform 1 0 49036 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_529
timestamp 1666464484
transform 1 0 49772 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1666464484
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1666464484
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1666464484
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1666464484
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1666464484
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1666464484
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1666464484
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1666464484
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_613
timestamp 1666464484
transform 1 0 57500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_623
timestamp 1666464484
transform 1 0 58420 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_3
timestamp 1666464484
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_9
timestamp 1666464484
transform 1 0 1932 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_18
timestamp 1666464484
transform 1 0 2760 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_30
timestamp 1666464484
transform 1 0 3864 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_42
timestamp 1666464484
transform 1 0 4968 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1666464484
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1666464484
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1666464484
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1666464484
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1666464484
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1666464484
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1666464484
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1666464484
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_122
timestamp 1666464484
transform 1 0 12328 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_134
timestamp 1666464484
transform 1 0 13432 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_146
timestamp 1666464484
transform 1 0 14536 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_158
timestamp 1666464484
transform 1 0 15640 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1666464484
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1666464484
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_181
timestamp 1666464484
transform 1 0 17756 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_189
timestamp 1666464484
transform 1 0 18492 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_198
timestamp 1666464484
transform 1 0 19320 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1666464484
transform 1 0 21528 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_225
timestamp 1666464484
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_244
timestamp 1666464484
transform 1 0 23552 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_256
timestamp 1666464484
transform 1 0 24656 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_268
timestamp 1666464484
transform 1 0 25760 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1666464484
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1666464484
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1666464484
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1666464484
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1666464484
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1666464484
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1666464484
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1666464484
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1666464484
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1666464484
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1666464484
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1666464484
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1666464484
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1666464484
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1666464484
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1666464484
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1666464484
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1666464484
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1666464484
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1666464484
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1666464484
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1666464484
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1666464484
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1666464484
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1666464484
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1666464484
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1666464484
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1666464484
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1666464484
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1666464484
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1666464484
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1666464484
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1666464484
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1666464484
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1666464484
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1666464484
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_617
timestamp 1666464484
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_66_3
timestamp 1666464484
transform 1 0 1380 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_26
timestamp 1666464484
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1666464484
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1666464484
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1666464484
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1666464484
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1666464484
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1666464484
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1666464484
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1666464484
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1666464484
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1666464484
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1666464484
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1666464484
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1666464484
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1666464484
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1666464484
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1666464484
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1666464484
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1666464484
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_197
timestamp 1666464484
transform 1 0 19228 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_203
timestamp 1666464484
transform 1 0 19780 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_216
timestamp 1666464484
transform 1 0 20976 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_229
timestamp 1666464484
transform 1 0 22172 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_241
timestamp 1666464484
transform 1 0 23276 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_249
timestamp 1666464484
transform 1 0 24012 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1666464484
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1666464484
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1666464484
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1666464484
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1666464484
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1666464484
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1666464484
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1666464484
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1666464484
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1666464484
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1666464484
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1666464484
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1666464484
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1666464484
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1666464484
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1666464484
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1666464484
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1666464484
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1666464484
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1666464484
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1666464484
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1666464484
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1666464484
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1666464484
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1666464484
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1666464484
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1666464484
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1666464484
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1666464484
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1666464484
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1666464484
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1666464484
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1666464484
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1666464484
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1666464484
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1666464484
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1666464484
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_601
timestamp 1666464484
transform 1 0 56396 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_613
timestamp 1666464484
transform 1 0 57500 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_623
timestamp 1666464484
transform 1 0 58420 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1666464484
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_9
timestamp 1666464484
transform 1 0 1932 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_21
timestamp 1666464484
transform 1 0 3036 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_33
timestamp 1666464484
transform 1 0 4140 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_45
timestamp 1666464484
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1666464484
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1666464484
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1666464484
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1666464484
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1666464484
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1666464484
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666464484
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1666464484
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1666464484
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1666464484
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1666464484
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1666464484
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1666464484
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1666464484
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1666464484
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1666464484
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_205
timestamp 1666464484
transform 1 0 19964 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_209
timestamp 1666464484
transform 1 0 20332 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_218
timestamp 1666464484
transform 1 0 21160 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_225
timestamp 1666464484
transform 1 0 21804 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_233
timestamp 1666464484
transform 1 0 22540 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_242
timestamp 1666464484
transform 1 0 23368 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_254
timestamp 1666464484
transform 1 0 24472 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_266
timestamp 1666464484
transform 1 0 25576 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_278
timestamp 1666464484
transform 1 0 26680 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1666464484
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1666464484
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1666464484
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1666464484
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1666464484
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1666464484
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1666464484
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1666464484
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1666464484
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1666464484
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1666464484
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1666464484
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1666464484
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1666464484
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1666464484
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1666464484
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1666464484
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1666464484
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1666464484
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1666464484
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1666464484
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1666464484
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1666464484
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1666464484
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1666464484
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1666464484
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1666464484
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1666464484
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1666464484
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1666464484
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1666464484
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1666464484
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1666464484
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1666464484
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1666464484
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1666464484
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_617
timestamp 1666464484
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1666464484
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_9
timestamp 1666464484
transform 1 0 1932 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_21
timestamp 1666464484
transform 1 0 3036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1666464484
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1666464484
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1666464484
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1666464484
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1666464484
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1666464484
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1666464484
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1666464484
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1666464484
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1666464484
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1666464484
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1666464484
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1666464484
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1666464484
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1666464484
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1666464484
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1666464484
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1666464484
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1666464484
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1666464484
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1666464484
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1666464484
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_233
timestamp 1666464484
transform 1 0 22540 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_237
timestamp 1666464484
transform 1 0 22908 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_247
timestamp 1666464484
transform 1 0 23828 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1666464484
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1666464484
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1666464484
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1666464484
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1666464484
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1666464484
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1666464484
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1666464484
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1666464484
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1666464484
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1666464484
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1666464484
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1666464484
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1666464484
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1666464484
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1666464484
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1666464484
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1666464484
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1666464484
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1666464484
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1666464484
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1666464484
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1666464484
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1666464484
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1666464484
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1666464484
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1666464484
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1666464484
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1666464484
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1666464484
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1666464484
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1666464484
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1666464484
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1666464484
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1666464484
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1666464484
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1666464484
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1666464484
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_601
timestamp 1666464484
transform 1 0 56396 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_613
timestamp 1666464484
transform 1 0 57500 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_623
timestamp 1666464484
transform 1 0 58420 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_3
timestamp 1666464484
transform 1 0 1380 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_9
timestamp 1666464484
transform 1 0 1932 0 -1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_23
timestamp 1666464484
transform 1 0 3220 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_35
timestamp 1666464484
transform 1 0 4324 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_47
timestamp 1666464484
transform 1 0 5428 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1666464484
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1666464484
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1666464484
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1666464484
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1666464484
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1666464484
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1666464484
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1666464484
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1666464484
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1666464484
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1666464484
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1666464484
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1666464484
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1666464484
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1666464484
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1666464484
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1666464484
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1666464484
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1666464484
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1666464484
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1666464484
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1666464484
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1666464484
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1666464484
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1666464484
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1666464484
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1666464484
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1666464484
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1666464484
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1666464484
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1666464484
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1666464484
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1666464484
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1666464484
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1666464484
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1666464484
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1666464484
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1666464484
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1666464484
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1666464484
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1666464484
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1666464484
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1666464484
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1666464484
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1666464484
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1666464484
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1666464484
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1666464484
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1666464484
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1666464484
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1666464484
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1666464484
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1666464484
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1666464484
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1666464484
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1666464484
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1666464484
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1666464484
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1666464484
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1666464484
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1666464484
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_617
timestamp 1666464484
transform 1 0 57868 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_623
timestamp 1666464484
transform 1 0 58420 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1666464484
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_9
timestamp 1666464484
transform 1 0 1932 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_21
timestamp 1666464484
transform 1 0 3036 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1666464484
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1666464484
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1666464484
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1666464484
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1666464484
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1666464484
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1666464484
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1666464484
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1666464484
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1666464484
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1666464484
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1666464484
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1666464484
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1666464484
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1666464484
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1666464484
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1666464484
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1666464484
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1666464484
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1666464484
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1666464484
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1666464484
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_233
timestamp 1666464484
transform 1 0 22540 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_241
timestamp 1666464484
transform 1 0 23276 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_249
timestamp 1666464484
transform 1 0 24012 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1666464484
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1666464484
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1666464484
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1666464484
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1666464484
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1666464484
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1666464484
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1666464484
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1666464484
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1666464484
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1666464484
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1666464484
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1666464484
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1666464484
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1666464484
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1666464484
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1666464484
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1666464484
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1666464484
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1666464484
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1666464484
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1666464484
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1666464484
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1666464484
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1666464484
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1666464484
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1666464484
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1666464484
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1666464484
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1666464484
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1666464484
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1666464484
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1666464484
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1666464484
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1666464484
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1666464484
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1666464484
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1666464484
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_613
timestamp 1666464484
transform 1 0 57500 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_623
timestamp 1666464484
transform 1 0 58420 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1666464484
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_9
timestamp 1666464484
transform 1 0 1932 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_21
timestamp 1666464484
transform 1 0 3036 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_27
timestamp 1666464484
transform 1 0 3588 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_36
timestamp 1666464484
transform 1 0 4416 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_48
timestamp 1666464484
transform 1 0 5520 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1666464484
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1666464484
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1666464484
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1666464484
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1666464484
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1666464484
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1666464484
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1666464484
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1666464484
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1666464484
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1666464484
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1666464484
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1666464484
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1666464484
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1666464484
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1666464484
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1666464484
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1666464484
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1666464484
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1666464484
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1666464484
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1666464484
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1666464484
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1666464484
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1666464484
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1666464484
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1666464484
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1666464484
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1666464484
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1666464484
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1666464484
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1666464484
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1666464484
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1666464484
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1666464484
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1666464484
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1666464484
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1666464484
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1666464484
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1666464484
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1666464484
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1666464484
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1666464484
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1666464484
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1666464484
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1666464484
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1666464484
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1666464484
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1666464484
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1666464484
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1666464484
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1666464484
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1666464484
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1666464484
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1666464484
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1666464484
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1666464484
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1666464484
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1666464484
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1666464484
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1666464484
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1666464484
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_9
timestamp 1666464484
transform 1 0 1932 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_21
timestamp 1666464484
transform 1 0 3036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1666464484
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1666464484
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1666464484
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1666464484
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1666464484
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1666464484
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1666464484
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1666464484
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1666464484
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1666464484
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1666464484
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1666464484
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1666464484
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1666464484
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1666464484
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1666464484
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1666464484
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1666464484
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1666464484
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1666464484
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1666464484
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1666464484
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_233
timestamp 1666464484
transform 1 0 22540 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_241
timestamp 1666464484
transform 1 0 23276 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_249
timestamp 1666464484
transform 1 0 24012 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1666464484
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1666464484
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1666464484
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1666464484
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1666464484
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1666464484
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1666464484
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1666464484
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1666464484
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1666464484
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1666464484
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1666464484
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1666464484
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1666464484
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1666464484
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1666464484
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1666464484
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1666464484
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1666464484
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1666464484
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1666464484
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1666464484
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1666464484
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1666464484
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1666464484
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1666464484
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1666464484
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1666464484
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1666464484
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1666464484
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1666464484
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1666464484
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1666464484
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1666464484
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1666464484
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1666464484
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1666464484
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_601
timestamp 1666464484
transform 1 0 56396 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_613
timestamp 1666464484
transform 1 0 57500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_623
timestamp 1666464484
transform 1 0 58420 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_3
timestamp 1666464484
transform 1 0 1380 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_9
timestamp 1666464484
transform 1 0 1932 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_21
timestamp 1666464484
transform 1 0 3036 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_33
timestamp 1666464484
transform 1 0 4140 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_43
timestamp 1666464484
transform 1 0 5060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1666464484
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1666464484
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1666464484
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1666464484
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1666464484
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1666464484
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1666464484
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1666464484
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1666464484
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1666464484
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1666464484
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1666464484
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1666464484
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1666464484
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1666464484
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1666464484
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1666464484
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1666464484
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1666464484
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1666464484
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_244
timestamp 1666464484
transform 1 0 23552 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_256
timestamp 1666464484
transform 1 0 24656 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_268
timestamp 1666464484
transform 1 0 25760 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1666464484
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1666464484
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1666464484
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1666464484
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1666464484
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1666464484
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1666464484
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1666464484
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1666464484
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1666464484
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1666464484
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1666464484
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1666464484
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1666464484
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1666464484
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1666464484
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1666464484
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1666464484
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1666464484
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1666464484
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1666464484
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1666464484
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1666464484
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1666464484
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1666464484
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1666464484
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1666464484
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1666464484
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1666464484
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1666464484
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1666464484
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1666464484
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1666464484
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1666464484
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1666464484
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1666464484
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1666464484
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1666464484
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_11
timestamp 1666464484
transform 1 0 2116 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_23
timestamp 1666464484
transform 1 0 3220 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1666464484
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1666464484
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1666464484
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1666464484
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1666464484
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1666464484
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1666464484
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1666464484
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1666464484
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1666464484
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1666464484
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1666464484
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1666464484
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1666464484
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1666464484
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1666464484
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1666464484
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1666464484
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1666464484
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1666464484
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1666464484
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1666464484
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_233
timestamp 1666464484
transform 1 0 22540 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_246
timestamp 1666464484
transform 1 0 23736 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1666464484
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1666464484
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1666464484
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1666464484
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1666464484
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1666464484
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1666464484
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1666464484
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1666464484
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1666464484
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1666464484
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1666464484
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1666464484
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1666464484
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1666464484
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1666464484
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1666464484
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1666464484
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1666464484
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1666464484
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1666464484
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1666464484
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1666464484
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1666464484
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1666464484
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1666464484
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1666464484
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1666464484
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1666464484
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1666464484
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1666464484
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1666464484
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1666464484
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1666464484
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1666464484
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1666464484
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1666464484
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_601
timestamp 1666464484
transform 1 0 56396 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_613
timestamp 1666464484
transform 1 0 57500 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_623
timestamp 1666464484
transform 1 0 58420 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1666464484
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_9
timestamp 1666464484
transform 1 0 1932 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_21
timestamp 1666464484
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_33
timestamp 1666464484
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1666464484
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1666464484
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1666464484
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1666464484
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1666464484
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1666464484
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1666464484
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1666464484
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1666464484
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1666464484
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1666464484
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1666464484
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1666464484
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1666464484
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1666464484
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1666464484
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1666464484
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1666464484
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1666464484
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1666464484
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1666464484
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1666464484
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1666464484
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1666464484
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1666464484
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1666464484
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1666464484
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1666464484
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1666464484
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1666464484
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1666464484
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1666464484
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1666464484
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1666464484
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1666464484
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1666464484
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1666464484
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1666464484
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1666464484
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1666464484
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1666464484
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1666464484
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1666464484
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1666464484
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1666464484
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1666464484
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1666464484
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1666464484
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1666464484
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1666464484
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1666464484
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1666464484
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1666464484
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1666464484
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1666464484
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1666464484
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1666464484
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1666464484
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1666464484
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1666464484
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1666464484
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1666464484
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_617
timestamp 1666464484
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1666464484
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1666464484
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1666464484
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1666464484
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1666464484
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1666464484
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1666464484
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1666464484
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1666464484
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1666464484
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1666464484
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1666464484
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1666464484
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1666464484
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1666464484
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_141
timestamp 1666464484
transform 1 0 14076 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_149
timestamp 1666464484
transform 1 0 14812 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1666464484
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1666464484
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1666464484
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1666464484
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1666464484
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1666464484
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1666464484
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1666464484
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1666464484
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1666464484
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1666464484
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1666464484
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1666464484
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1666464484
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1666464484
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1666464484
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1666464484
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1666464484
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1666464484
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1666464484
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1666464484
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1666464484
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1666464484
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1666464484
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1666464484
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1666464484
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1666464484
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1666464484
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1666464484
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1666464484
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1666464484
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1666464484
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1666464484
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1666464484
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1666464484
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1666464484
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1666464484
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1666464484
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1666464484
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1666464484
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1666464484
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1666464484
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1666464484
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1666464484
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1666464484
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1666464484
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1666464484
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1666464484
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_613
timestamp 1666464484
transform 1 0 57500 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_623
timestamp 1666464484
transform 1 0 58420 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1666464484
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_9
timestamp 1666464484
transform 1 0 1932 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_21
timestamp 1666464484
transform 1 0 3036 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_33
timestamp 1666464484
transform 1 0 4140 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_45
timestamp 1666464484
transform 1 0 5244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_53
timestamp 1666464484
transform 1 0 5980 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1666464484
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1666464484
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1666464484
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1666464484
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1666464484
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1666464484
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1666464484
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1666464484
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1666464484
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1666464484
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1666464484
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1666464484
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1666464484
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1666464484
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1666464484
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1666464484
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1666464484
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1666464484
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1666464484
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1666464484
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1666464484
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1666464484
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1666464484
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1666464484
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1666464484
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1666464484
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1666464484
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1666464484
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1666464484
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1666464484
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1666464484
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1666464484
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1666464484
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1666464484
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1666464484
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1666464484
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1666464484
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1666464484
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1666464484
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1666464484
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1666464484
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1666464484
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1666464484
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1666464484
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1666464484
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1666464484
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1666464484
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1666464484
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1666464484
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1666464484
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1666464484
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1666464484
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1666464484
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1666464484
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1666464484
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1666464484
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1666464484
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1666464484
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1666464484
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1666464484
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_617
timestamp 1666464484
transform 1 0 57868 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1666464484
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_9
timestamp 1666464484
transform 1 0 1932 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_21
timestamp 1666464484
transform 1 0 3036 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1666464484
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1666464484
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1666464484
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1666464484
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1666464484
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1666464484
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1666464484
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1666464484
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1666464484
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1666464484
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1666464484
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1666464484
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1666464484
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1666464484
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1666464484
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1666464484
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1666464484
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1666464484
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1666464484
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1666464484
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1666464484
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1666464484
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1666464484
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1666464484
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1666464484
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1666464484
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1666464484
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1666464484
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1666464484
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1666464484
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1666464484
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1666464484
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1666464484
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1666464484
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1666464484
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1666464484
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1666464484
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1666464484
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1666464484
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1666464484
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1666464484
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1666464484
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1666464484
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1666464484
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1666464484
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1666464484
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1666464484
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1666464484
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1666464484
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1666464484
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1666464484
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1666464484
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1666464484
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1666464484
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1666464484
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1666464484
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1666464484
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1666464484
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1666464484
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1666464484
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1666464484
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1666464484
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_601
timestamp 1666464484
transform 1 0 56396 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_613
timestamp 1666464484
transform 1 0 57500 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_623
timestamp 1666464484
transform 1 0 58420 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_3
timestamp 1666464484
transform 1 0 1380 0 -1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_9
timestamp 1666464484
transform 1 0 1932 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_21
timestamp 1666464484
transform 1 0 3036 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_33
timestamp 1666464484
transform 1 0 4140 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_45
timestamp 1666464484
transform 1 0 5244 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_53
timestamp 1666464484
transform 1 0 5980 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1666464484
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1666464484
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1666464484
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1666464484
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1666464484
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1666464484
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1666464484
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1666464484
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1666464484
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1666464484
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1666464484
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1666464484
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1666464484
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1666464484
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1666464484
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1666464484
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1666464484
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1666464484
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1666464484
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1666464484
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1666464484
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1666464484
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1666464484
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1666464484
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1666464484
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1666464484
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1666464484
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1666464484
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1666464484
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1666464484
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1666464484
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1666464484
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1666464484
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1666464484
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1666464484
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1666464484
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1666464484
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1666464484
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1666464484
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1666464484
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1666464484
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1666464484
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1666464484
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1666464484
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1666464484
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1666464484
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1666464484
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1666464484
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1666464484
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1666464484
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1666464484
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1666464484
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1666464484
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1666464484
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1666464484
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1666464484
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1666464484
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1666464484
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1666464484
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1666464484
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1666464484
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1666464484
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_9
timestamp 1666464484
transform 1 0 1932 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1666464484
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1666464484
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1666464484
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1666464484
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1666464484
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1666464484
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1666464484
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1666464484
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1666464484
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1666464484
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1666464484
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1666464484
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1666464484
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1666464484
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1666464484
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1666464484
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1666464484
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1666464484
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1666464484
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1666464484
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1666464484
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1666464484
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_221
timestamp 1666464484
transform 1 0 21436 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_229
timestamp 1666464484
transform 1 0 22172 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_80_234
timestamp 1666464484
transform 1 0 22632 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_243
timestamp 1666464484
transform 1 0 23460 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1666464484
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1666464484
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1666464484
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1666464484
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1666464484
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1666464484
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1666464484
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1666464484
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1666464484
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1666464484
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1666464484
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1666464484
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1666464484
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1666464484
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1666464484
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1666464484
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1666464484
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1666464484
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1666464484
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1666464484
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1666464484
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1666464484
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1666464484
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1666464484
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1666464484
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1666464484
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1666464484
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1666464484
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1666464484
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1666464484
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1666464484
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1666464484
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1666464484
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1666464484
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1666464484
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1666464484
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1666464484
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1666464484
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1666464484
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_613
timestamp 1666464484
transform 1 0 57500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_623
timestamp 1666464484
transform 1 0 58420 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1666464484
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1666464484
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1666464484
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1666464484
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1666464484
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1666464484
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1666464484
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1666464484
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1666464484
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1666464484
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1666464484
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1666464484
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1666464484
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1666464484
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1666464484
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1666464484
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1666464484
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1666464484
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1666464484
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1666464484
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1666464484
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1666464484
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1666464484
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1666464484
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1666464484
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1666464484
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1666464484
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1666464484
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1666464484
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1666464484
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1666464484
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1666464484
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1666464484
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1666464484
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1666464484
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1666464484
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1666464484
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1666464484
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1666464484
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1666464484
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1666464484
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1666464484
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1666464484
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1666464484
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1666464484
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1666464484
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1666464484
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1666464484
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1666464484
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1666464484
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1666464484
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1666464484
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1666464484
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1666464484
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1666464484
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1666464484
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1666464484
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1666464484
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1666464484
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1666464484
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1666464484
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1666464484
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1666464484
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1666464484
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1666464484
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1666464484
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1666464484
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1666464484
transform 1 0 1380 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_9
timestamp 1666464484
transform 1 0 1932 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1666464484
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1666464484
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1666464484
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1666464484
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1666464484
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1666464484
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1666464484
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1666464484
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1666464484
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1666464484
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1666464484
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1666464484
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1666464484
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1666464484
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1666464484
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1666464484
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1666464484
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1666464484
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1666464484
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1666464484
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1666464484
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1666464484
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1666464484
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1666464484
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1666464484
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1666464484
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1666464484
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1666464484
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1666464484
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1666464484
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1666464484
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1666464484
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1666464484
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1666464484
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1666464484
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1666464484
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1666464484
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1666464484
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1666464484
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1666464484
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1666464484
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1666464484
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1666464484
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1666464484
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1666464484
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1666464484
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1666464484
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1666464484
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1666464484
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1666464484
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1666464484
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1666464484
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1666464484
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1666464484
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1666464484
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1666464484
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1666464484
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1666464484
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1666464484
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1666464484
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1666464484
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1666464484
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1666464484
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1666464484
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_613
timestamp 1666464484
transform 1 0 57500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_623
timestamp 1666464484
transform 1 0 58420 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_3
timestamp 1666464484
transform 1 0 1380 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_9
timestamp 1666464484
transform 1 0 1932 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_21
timestamp 1666464484
transform 1 0 3036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_33
timestamp 1666464484
transform 1 0 4140 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_45
timestamp 1666464484
transform 1 0 5244 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_53
timestamp 1666464484
transform 1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1666464484
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1666464484
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1666464484
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1666464484
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1666464484
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1666464484
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1666464484
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1666464484
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1666464484
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1666464484
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1666464484
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1666464484
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1666464484
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1666464484
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1666464484
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1666464484
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1666464484
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1666464484
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1666464484
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1666464484
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1666464484
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1666464484
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1666464484
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1666464484
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1666464484
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1666464484
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1666464484
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1666464484
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1666464484
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1666464484
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1666464484
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1666464484
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1666464484
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1666464484
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1666464484
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1666464484
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1666464484
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1666464484
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1666464484
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1666464484
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1666464484
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1666464484
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1666464484
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1666464484
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1666464484
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1666464484
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1666464484
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1666464484
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1666464484
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1666464484
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1666464484
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1666464484
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1666464484
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1666464484
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1666464484
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1666464484
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1666464484
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1666464484
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1666464484
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1666464484
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1666464484
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1666464484
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_9
timestamp 1666464484
transform 1 0 1932 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_21
timestamp 1666464484
transform 1 0 3036 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1666464484
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1666464484
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1666464484
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1666464484
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1666464484
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1666464484
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1666464484
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1666464484
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1666464484
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1666464484
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1666464484
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1666464484
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1666464484
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1666464484
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1666464484
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1666464484
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1666464484
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1666464484
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1666464484
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1666464484
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1666464484
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1666464484
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1666464484
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1666464484
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1666464484
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1666464484
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1666464484
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1666464484
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1666464484
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1666464484
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1666464484
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1666464484
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1666464484
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1666464484
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1666464484
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1666464484
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1666464484
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1666464484
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1666464484
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1666464484
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1666464484
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1666464484
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1666464484
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1666464484
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1666464484
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1666464484
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1666464484
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1666464484
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1666464484
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1666464484
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1666464484
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1666464484
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1666464484
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1666464484
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1666464484
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1666464484
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1666464484
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1666464484
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1666464484
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1666464484
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1666464484
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1666464484
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_601
timestamp 1666464484
transform 1 0 56396 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_613
timestamp 1666464484
transform 1 0 57500 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_623
timestamp 1666464484
transform 1 0 58420 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_3
timestamp 1666464484
transform 1 0 1380 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_9
timestamp 1666464484
transform 1 0 1932 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_21
timestamp 1666464484
transform 1 0 3036 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_33
timestamp 1666464484
transform 1 0 4140 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_45
timestamp 1666464484
transform 1 0 5244 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_53
timestamp 1666464484
transform 1 0 5980 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1666464484
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1666464484
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1666464484
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1666464484
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1666464484
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1666464484
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1666464484
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1666464484
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1666464484
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1666464484
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1666464484
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1666464484
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1666464484
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1666464484
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_193
timestamp 1666464484
transform 1 0 18860 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_201
timestamp 1666464484
transform 1 0 19596 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_209
timestamp 1666464484
transform 1 0 20332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_221
timestamp 1666464484
transform 1 0 21436 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_225
timestamp 1666464484
transform 1 0 21804 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_235
timestamp 1666464484
transform 1 0 22724 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_239
timestamp 1666464484
transform 1 0 23092 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_251
timestamp 1666464484
transform 1 0 24196 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_263
timestamp 1666464484
transform 1 0 25300 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_275
timestamp 1666464484
transform 1 0 26404 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1666464484
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1666464484
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1666464484
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1666464484
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1666464484
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1666464484
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1666464484
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1666464484
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1666464484
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1666464484
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1666464484
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1666464484
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1666464484
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1666464484
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1666464484
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1666464484
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1666464484
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1666464484
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1666464484
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1666464484
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1666464484
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1666464484
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1666464484
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1666464484
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1666464484
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1666464484
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1666464484
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1666464484
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1666464484
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1666464484
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1666464484
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1666464484
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1666464484
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1666464484
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1666464484
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1666464484
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1666464484
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_617
timestamp 1666464484
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1666464484
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1666464484
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1666464484
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1666464484
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1666464484
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1666464484
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1666464484
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1666464484
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1666464484
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1666464484
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1666464484
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1666464484
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1666464484
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1666464484
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1666464484
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1666464484
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1666464484
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1666464484
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1666464484
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1666464484
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1666464484
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1666464484
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_209
timestamp 1666464484
transform 1 0 20332 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_217
timestamp 1666464484
transform 1 0 21068 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_225
timestamp 1666464484
transform 1 0 21804 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_237
timestamp 1666464484
transform 1 0 22908 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_249
timestamp 1666464484
transform 1 0 24012 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1666464484
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1666464484
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1666464484
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1666464484
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1666464484
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1666464484
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1666464484
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1666464484
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1666464484
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1666464484
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1666464484
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1666464484
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1666464484
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1666464484
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1666464484
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1666464484
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1666464484
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1666464484
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1666464484
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1666464484
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1666464484
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1666464484
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1666464484
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1666464484
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1666464484
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1666464484
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1666464484
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1666464484
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1666464484
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1666464484
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1666464484
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1666464484
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1666464484
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1666464484
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1666464484
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1666464484
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1666464484
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1666464484
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_613
timestamp 1666464484
transform 1 0 57500 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_623
timestamp 1666464484
transform 1 0 58420 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_3
timestamp 1666464484
transform 1 0 1380 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_9
timestamp 1666464484
transform 1 0 1932 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_21
timestamp 1666464484
transform 1 0 3036 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_33
timestamp 1666464484
transform 1 0 4140 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_45
timestamp 1666464484
transform 1 0 5244 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_53
timestamp 1666464484
transform 1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1666464484
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1666464484
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1666464484
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1666464484
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1666464484
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1666464484
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1666464484
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1666464484
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1666464484
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1666464484
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1666464484
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1666464484
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1666464484
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1666464484
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1666464484
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_205
timestamp 1666464484
transform 1 0 19964 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_87_218
timestamp 1666464484
transform 1 0 21160 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1666464484
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1666464484
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1666464484
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1666464484
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1666464484
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1666464484
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1666464484
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1666464484
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1666464484
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1666464484
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1666464484
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1666464484
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1666464484
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1666464484
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1666464484
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1666464484
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1666464484
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1666464484
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1666464484
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1666464484
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1666464484
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1666464484
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1666464484
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1666464484
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1666464484
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1666464484
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1666464484
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1666464484
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1666464484
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1666464484
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1666464484
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1666464484
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1666464484
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1666464484
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1666464484
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1666464484
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1666464484
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1666464484
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1666464484
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1666464484
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1666464484
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1666464484
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1666464484
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_3
timestamp 1666464484
transform 1 0 1380 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_9
timestamp 1666464484
transform 1 0 1932 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_21
timestamp 1666464484
transform 1 0 3036 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1666464484
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1666464484
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1666464484
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1666464484
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1666464484
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1666464484
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1666464484
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1666464484
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1666464484
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1666464484
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1666464484
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1666464484
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1666464484
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1666464484
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1666464484
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1666464484
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1666464484
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1666464484
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1666464484
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1666464484
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1666464484
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1666464484
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1666464484
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1666464484
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1666464484
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1666464484
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1666464484
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1666464484
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1666464484
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1666464484
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1666464484
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1666464484
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1666464484
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1666464484
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1666464484
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1666464484
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1666464484
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1666464484
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1666464484
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1666464484
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1666464484
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1666464484
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1666464484
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1666464484
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1666464484
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1666464484
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1666464484
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1666464484
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1666464484
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1666464484
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1666464484
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1666464484
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1666464484
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1666464484
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1666464484
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1666464484
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1666464484
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1666464484
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1666464484
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1666464484
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1666464484
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1666464484
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1666464484
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_613
timestamp 1666464484
transform 1 0 57500 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_623
timestamp 1666464484
transform 1 0 58420 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1666464484
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_9
timestamp 1666464484
transform 1 0 1932 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_21
timestamp 1666464484
transform 1 0 3036 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_33
timestamp 1666464484
transform 1 0 4140 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_45
timestamp 1666464484
transform 1 0 5244 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_53
timestamp 1666464484
transform 1 0 5980 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1666464484
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1666464484
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1666464484
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1666464484
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1666464484
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1666464484
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1666464484
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1666464484
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1666464484
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1666464484
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1666464484
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1666464484
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1666464484
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1666464484
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1666464484
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1666464484
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1666464484
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1666464484
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1666464484
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1666464484
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1666464484
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1666464484
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1666464484
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1666464484
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1666464484
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1666464484
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1666464484
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1666464484
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1666464484
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1666464484
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1666464484
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1666464484
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1666464484
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1666464484
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1666464484
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1666464484
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1666464484
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1666464484
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1666464484
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1666464484
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1666464484
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1666464484
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1666464484
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1666464484
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1666464484
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1666464484
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1666464484
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1666464484
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1666464484
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1666464484
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1666464484
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1666464484
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1666464484
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1666464484
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1666464484
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1666464484
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1666464484
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1666464484
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1666464484
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1666464484
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1666464484
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_3
timestamp 1666464484
transform 1 0 1380 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_9
timestamp 1666464484
transform 1 0 1932 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_21
timestamp 1666464484
transform 1 0 3036 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1666464484
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1666464484
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1666464484
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1666464484
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1666464484
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1666464484
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1666464484
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1666464484
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1666464484
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1666464484
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1666464484
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1666464484
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1666464484
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1666464484
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1666464484
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1666464484
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1666464484
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1666464484
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1666464484
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1666464484
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1666464484
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_221
timestamp 1666464484
transform 1 0 21436 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_90_229
timestamp 1666464484
transform 1 0 22172 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_240
timestamp 1666464484
transform 1 0 23184 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1666464484
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1666464484
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1666464484
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1666464484
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1666464484
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1666464484
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1666464484
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1666464484
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1666464484
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1666464484
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1666464484
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1666464484
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1666464484
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1666464484
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1666464484
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1666464484
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1666464484
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1666464484
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1666464484
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1666464484
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1666464484
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1666464484
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1666464484
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1666464484
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1666464484
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1666464484
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1666464484
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1666464484
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1666464484
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1666464484
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1666464484
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1666464484
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1666464484
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1666464484
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1666464484
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1666464484
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1666464484
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1666464484
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_613
timestamp 1666464484
transform 1 0 57500 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_619
timestamp 1666464484
transform 1 0 58052 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_623
timestamp 1666464484
transform 1 0 58420 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1666464484
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1666464484
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1666464484
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_39
timestamp 1666464484
transform 1 0 4692 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_43
timestamp 1666464484
transform 1 0 5060 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_52
timestamp 1666464484
transform 1 0 5888 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1666464484
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1666464484
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1666464484
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1666464484
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1666464484
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1666464484
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1666464484
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1666464484
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1666464484
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1666464484
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1666464484
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1666464484
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1666464484
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1666464484
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1666464484
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1666464484
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1666464484
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1666464484
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1666464484
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1666464484
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1666464484
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1666464484
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1666464484
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1666464484
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1666464484
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1666464484
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1666464484
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1666464484
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1666464484
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1666464484
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1666464484
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1666464484
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1666464484
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1666464484
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1666464484
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1666464484
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1666464484
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1666464484
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1666464484
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1666464484
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1666464484
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1666464484
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1666464484
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1666464484
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1666464484
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1666464484
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1666464484
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1666464484
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1666464484
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1666464484
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1666464484
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1666464484
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1666464484
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1666464484
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1666464484
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1666464484
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1666464484
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1666464484
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1666464484
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1666464484
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1666464484
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1666464484
transform 1 0 1380 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_9
timestamp 1666464484
transform 1 0 1932 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_21
timestamp 1666464484
transform 1 0 3036 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1666464484
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1666464484
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1666464484
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1666464484
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1666464484
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1666464484
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1666464484
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1666464484
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1666464484
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1666464484
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1666464484
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1666464484
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1666464484
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1666464484
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1666464484
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1666464484
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1666464484
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1666464484
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1666464484
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1666464484
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1666464484
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1666464484
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1666464484
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1666464484
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1666464484
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1666464484
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1666464484
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1666464484
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1666464484
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1666464484
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1666464484
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1666464484
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1666464484
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1666464484
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1666464484
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1666464484
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1666464484
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1666464484
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1666464484
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1666464484
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1666464484
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1666464484
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1666464484
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1666464484
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1666464484
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1666464484
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1666464484
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1666464484
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1666464484
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1666464484
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1666464484
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1666464484
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1666464484
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1666464484
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1666464484
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1666464484
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1666464484
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1666464484
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1666464484
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1666464484
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1666464484
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1666464484
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1666464484
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1666464484
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1666464484
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_9
timestamp 1666464484
transform 1 0 1932 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_21
timestamp 1666464484
transform 1 0 3036 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_33
timestamp 1666464484
transform 1 0 4140 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_45
timestamp 1666464484
transform 1 0 5244 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_53
timestamp 1666464484
transform 1 0 5980 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1666464484
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1666464484
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1666464484
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1666464484
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1666464484
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1666464484
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1666464484
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1666464484
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1666464484
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1666464484
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1666464484
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1666464484
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1666464484
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1666464484
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1666464484
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1666464484
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1666464484
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1666464484
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1666464484
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1666464484
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1666464484
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1666464484
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1666464484
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1666464484
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1666464484
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1666464484
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1666464484
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1666464484
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1666464484
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1666464484
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1666464484
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1666464484
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1666464484
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1666464484
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1666464484
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1666464484
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1666464484
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1666464484
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1666464484
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1666464484
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1666464484
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1666464484
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1666464484
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1666464484
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1666464484
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1666464484
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1666464484
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1666464484
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1666464484
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1666464484
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1666464484
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1666464484
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1666464484
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1666464484
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1666464484
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1666464484
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1666464484
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1666464484
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1666464484
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1666464484
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_93_617
timestamp 1666464484
transform 1 0 57868 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_623
timestamp 1666464484
transform 1 0 58420 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1666464484
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_9
timestamp 1666464484
transform 1 0 1932 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_21
timestamp 1666464484
transform 1 0 3036 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1666464484
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1666464484
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1666464484
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1666464484
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1666464484
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1666464484
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1666464484
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1666464484
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1666464484
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1666464484
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1666464484
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1666464484
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1666464484
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1666464484
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1666464484
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1666464484
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1666464484
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1666464484
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1666464484
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1666464484
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1666464484
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1666464484
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1666464484
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1666464484
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1666464484
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1666464484
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1666464484
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1666464484
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1666464484
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1666464484
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1666464484
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1666464484
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1666464484
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1666464484
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1666464484
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1666464484
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1666464484
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1666464484
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1666464484
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1666464484
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1666464484
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1666464484
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1666464484
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1666464484
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1666464484
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1666464484
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1666464484
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1666464484
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1666464484
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1666464484
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1666464484
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1666464484
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1666464484
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1666464484
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1666464484
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1666464484
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1666464484
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1666464484
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1666464484
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1666464484
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1666464484
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1666464484
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1666464484
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1666464484
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_3
timestamp 1666464484
transform 1 0 1380 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_11
timestamp 1666464484
transform 1 0 2116 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_23
timestamp 1666464484
transform 1 0 3220 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_35
timestamp 1666464484
transform 1 0 4324 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_47
timestamp 1666464484
transform 1 0 5428 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1666464484
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1666464484
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1666464484
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1666464484
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1666464484
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1666464484
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1666464484
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1666464484
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1666464484
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1666464484
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1666464484
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1666464484
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1666464484
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1666464484
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1666464484
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1666464484
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1666464484
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1666464484
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1666464484
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1666464484
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1666464484
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1666464484
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1666464484
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1666464484
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1666464484
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1666464484
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1666464484
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1666464484
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1666464484
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1666464484
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1666464484
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1666464484
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1666464484
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1666464484
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1666464484
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1666464484
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1666464484
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1666464484
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1666464484
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1666464484
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1666464484
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1666464484
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1666464484
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_449
timestamp 1666464484
transform 1 0 42412 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_465
timestamp 1666464484
transform 1 0 43884 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_477
timestamp 1666464484
transform 1 0 44988 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_489
timestamp 1666464484
transform 1 0 46092 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_501
timestamp 1666464484
transform 1 0 47196 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1666464484
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1666464484
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1666464484
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1666464484
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1666464484
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1666464484
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1666464484
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1666464484
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1666464484
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1666464484
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1666464484
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1666464484
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_617
timestamp 1666464484
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1666464484
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1666464484
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1666464484
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1666464484
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1666464484
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1666464484
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1666464484
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1666464484
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1666464484
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1666464484
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1666464484
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1666464484
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1666464484
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1666464484
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1666464484
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1666464484
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1666464484
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1666464484
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1666464484
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1666464484
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1666464484
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1666464484
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1666464484
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1666464484
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1666464484
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1666464484
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1666464484
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1666464484
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1666464484
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1666464484
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1666464484
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1666464484
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1666464484
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1666464484
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1666464484
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1666464484
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1666464484
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1666464484
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1666464484
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1666464484
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1666464484
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1666464484
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1666464484
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1666464484
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1666464484
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1666464484
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1666464484
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1666464484
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1666464484
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1666464484
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1666464484
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1666464484
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1666464484
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1666464484
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1666464484
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1666464484
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1666464484
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1666464484
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1666464484
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1666464484
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1666464484
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1666464484
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1666464484
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1666464484
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1666464484
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_613
timestamp 1666464484
transform 1 0 57500 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_619
timestamp 1666464484
transform 1 0 58052 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_623
timestamp 1666464484
transform 1 0 58420 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_3
timestamp 1666464484
transform 1 0 1380 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_9
timestamp 1666464484
transform 1 0 1932 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_21
timestamp 1666464484
transform 1 0 3036 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_33
timestamp 1666464484
transform 1 0 4140 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_45
timestamp 1666464484
transform 1 0 5244 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_53
timestamp 1666464484
transform 1 0 5980 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1666464484
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1666464484
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1666464484
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1666464484
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1666464484
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1666464484
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1666464484
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1666464484
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1666464484
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1666464484
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1666464484
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1666464484
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1666464484
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1666464484
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1666464484
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1666464484
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1666464484
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1666464484
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1666464484
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1666464484
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1666464484
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1666464484
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1666464484
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1666464484
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1666464484
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1666464484
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1666464484
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1666464484
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1666464484
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1666464484
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1666464484
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1666464484
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1666464484
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1666464484
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1666464484
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1666464484
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1666464484
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1666464484
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1666464484
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1666464484
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1666464484
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1666464484
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_97_449
timestamp 1666464484
transform 1 0 42412 0 -1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_97_469
timestamp 1666464484
transform 1 0 44252 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_481
timestamp 1666464484
transform 1 0 45356 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_493
timestamp 1666464484
transform 1 0 46460 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_97_501
timestamp 1666464484
transform 1 0 47196 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1666464484
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1666464484
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1666464484
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1666464484
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1666464484
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1666464484
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1666464484
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1666464484
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1666464484
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1666464484
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1666464484
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1666464484
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_617
timestamp 1666464484
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_3
timestamp 1666464484
transform 1 0 1380 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_11
timestamp 1666464484
transform 1 0 2116 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_23
timestamp 1666464484
transform 1 0 3220 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1666464484
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1666464484
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1666464484
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1666464484
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1666464484
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1666464484
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1666464484
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1666464484
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1666464484
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1666464484
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1666464484
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1666464484
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1666464484
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1666464484
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1666464484
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1666464484
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1666464484
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1666464484
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1666464484
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1666464484
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1666464484
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1666464484
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1666464484
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1666464484
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1666464484
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1666464484
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1666464484
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1666464484
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1666464484
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1666464484
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1666464484
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1666464484
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1666464484
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1666464484
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1666464484
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1666464484
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1666464484
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1666464484
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1666464484
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1666464484
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1666464484
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1666464484
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1666464484
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1666464484
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1666464484
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1666464484
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1666464484
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1666464484
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1666464484
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1666464484
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1666464484
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1666464484
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1666464484
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1666464484
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1666464484
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1666464484
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1666464484
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1666464484
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1666464484
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1666464484
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1666464484
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1666464484
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1666464484
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1666464484
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_3
timestamp 1666464484
transform 1 0 1380 0 -1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_99_9
timestamp 1666464484
transform 1 0 1932 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_21
timestamp 1666464484
transform 1 0 3036 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_33
timestamp 1666464484
transform 1 0 4140 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_45
timestamp 1666464484
transform 1 0 5244 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_53
timestamp 1666464484
transform 1 0 5980 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1666464484
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1666464484
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1666464484
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1666464484
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1666464484
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1666464484
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1666464484
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1666464484
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1666464484
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_149
timestamp 1666464484
transform 1 0 14812 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_99_162
timestamp 1666464484
transform 1 0 16008 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1666464484
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1666464484
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1666464484
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1666464484
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1666464484
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1666464484
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1666464484
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1666464484
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1666464484
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1666464484
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1666464484
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1666464484
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1666464484
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1666464484
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_305
timestamp 1666464484
transform 1 0 29164 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_99_316
timestamp 1666464484
transform 1 0 30176 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_328
timestamp 1666464484
transform 1 0 31280 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1666464484
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_349
timestamp 1666464484
transform 1 0 33212 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_360
timestamp 1666464484
transform 1 0 34224 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1666464484
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1666464484
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1666464484
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1666464484
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1666464484
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1666464484
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1666464484
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1666464484
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1666464484
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1666464484
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1666464484
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1666464484
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1666464484
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1666464484
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1666464484
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1666464484
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1666464484
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1666464484
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1666464484
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1666464484
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1666464484
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1666464484
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1666464484
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1666464484
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1666464484
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1666464484
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1666464484
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_99_617
timestamp 1666464484
transform 1 0 57868 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1666464484
transform 1 0 58420 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_3
timestamp 1666464484
transform 1 0 1380 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_11
timestamp 1666464484
transform 1 0 2116 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_23
timestamp 1666464484
transform 1 0 3220 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1666464484
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1666464484
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1666464484
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1666464484
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1666464484
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1666464484
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1666464484
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1666464484
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1666464484
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1666464484
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1666464484
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1666464484
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1666464484
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1666464484
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1666464484
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1666464484
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1666464484
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1666464484
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1666464484
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1666464484
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1666464484
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_221
timestamp 1666464484
transform 1 0 21436 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_232
timestamp 1666464484
transform 1 0 22448 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_244
timestamp 1666464484
transform 1 0 23552 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1666464484
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1666464484
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1666464484
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1666464484
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1666464484
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1666464484
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1666464484
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1666464484
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1666464484
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1666464484
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1666464484
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1666464484
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1666464484
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1666464484
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1666464484
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1666464484
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1666464484
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1666464484
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1666464484
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1666464484
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1666464484
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_457
timestamp 1666464484
transform 1 0 43148 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_474
timestamp 1666464484
transform 1 0 44712 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1666464484
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1666464484
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1666464484
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1666464484
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1666464484
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1666464484
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1666464484
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1666464484
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_557
timestamp 1666464484
transform 1 0 52348 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_565
timestamp 1666464484
transform 1 0 53084 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_100_582
timestamp 1666464484
transform 1 0 54648 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1666464484
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1666464484
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_613
timestamp 1666464484
transform 1 0 57500 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_100_623
timestamp 1666464484
transform 1 0 58420 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1666464484
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1666464484
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_27
timestamp 1666464484
transform 1 0 3588 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_39
timestamp 1666464484
transform 1 0 4692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_51
timestamp 1666464484
transform 1 0 5796 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1666464484
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1666464484
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1666464484
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_81
timestamp 1666464484
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_93
timestamp 1666464484
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1666464484
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1666464484
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1666464484
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1666464484
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_137
timestamp 1666464484
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_149
timestamp 1666464484
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_161
timestamp 1666464484
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_167
timestamp 1666464484
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1666464484
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1666464484
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_193
timestamp 1666464484
transform 1 0 18860 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_201
timestamp 1666464484
transform 1 0 19596 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_205
timestamp 1666464484
transform 1 0 19964 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_214
timestamp 1666464484
transform 1 0 20792 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_222
timestamp 1666464484
transform 1 0 21528 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1666464484
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1666464484
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_249
timestamp 1666464484
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_261
timestamp 1666464484
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_273
timestamp 1666464484
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1666464484
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1666464484
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1666464484
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_305
timestamp 1666464484
transform 1 0 29164 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_334
timestamp 1666464484
transform 1 0 31832 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1666464484
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1666464484
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_361
timestamp 1666464484
transform 1 0 34316 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_369
timestamp 1666464484
transform 1 0 35052 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_388
timestamp 1666464484
transform 1 0 36800 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_393
timestamp 1666464484
transform 1 0 37260 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_401
timestamp 1666464484
transform 1 0 37996 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_409
timestamp 1666464484
transform 1 0 38732 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_421
timestamp 1666464484
transform 1 0 39836 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_433
timestamp 1666464484
transform 1 0 40940 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1666464484
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1666464484
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1666464484
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_473
timestamp 1666464484
transform 1 0 44620 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_485
timestamp 1666464484
transform 1 0 45724 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1666464484
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1666464484
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1666464484
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1666464484
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_529
timestamp 1666464484
transform 1 0 49772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_541
timestamp 1666464484
transform 1 0 50876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_553
timestamp 1666464484
transform 1 0 51980 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1666464484
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1666464484
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_587
timestamp 1666464484
transform 1 0 55108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_599
timestamp 1666464484
transform 1 0 56212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_611
timestamp 1666464484
transform 1 0 57316 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1666464484
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_617
timestamp 1666464484
transform 1 0 57868 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_623
timestamp 1666464484
transform 1 0 58420 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_102_3
timestamp 1666464484
transform 1 0 1380 0 1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_9
timestamp 1666464484
transform 1 0 1932 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_21
timestamp 1666464484
transform 1 0 3036 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1666464484
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1666464484
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1666464484
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1666464484
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_65
timestamp 1666464484
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1666464484
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1666464484
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_85
timestamp 1666464484
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_97
timestamp 1666464484
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_109
timestamp 1666464484
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_121
timestamp 1666464484
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1666464484
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1666464484
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_141
timestamp 1666464484
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_153
timestamp 1666464484
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_165
timestamp 1666464484
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_177
timestamp 1666464484
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_189
timestamp 1666464484
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_195
timestamp 1666464484
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_197
timestamp 1666464484
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_209
timestamp 1666464484
transform 1 0 20332 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_213
timestamp 1666464484
transform 1 0 20700 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_231
timestamp 1666464484
transform 1 0 22356 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_102_244
timestamp 1666464484
transform 1 0 23552 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_102_253
timestamp 1666464484
transform 1 0 24380 0 1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_263
timestamp 1666464484
transform 1 0 25300 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_275
timestamp 1666464484
transform 1 0 26404 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_287
timestamp 1666464484
transform 1 0 27508 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_299
timestamp 1666464484
transform 1 0 28612 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_102_307
timestamp 1666464484
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_309
timestamp 1666464484
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_321
timestamp 1666464484
transform 1 0 30636 0 1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_102_346
timestamp 1666464484
transform 1 0 32936 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_358
timestamp 1666464484
transform 1 0 34040 0 1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_102_365
timestamp 1666464484
transform 1 0 34684 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_377
timestamp 1666464484
transform 1 0 35788 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_389
timestamp 1666464484
transform 1 0 36892 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_401
timestamp 1666464484
transform 1 0 37996 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_102_412
timestamp 1666464484
transform 1 0 39008 0 1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_102_421
timestamp 1666464484
transform 1 0 39836 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_433
timestamp 1666464484
transform 1 0 40940 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_445
timestamp 1666464484
transform 1 0 42044 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_102_457
timestamp 1666464484
transform 1 0 43148 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_102_474
timestamp 1666464484
transform 1 0 44712 0 1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_477
timestamp 1666464484
transform 1 0 44988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_489
timestamp 1666464484
transform 1 0 46092 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_501
timestamp 1666464484
transform 1 0 47196 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_513
timestamp 1666464484
transform 1 0 48300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_525
timestamp 1666464484
transform 1 0 49404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_531
timestamp 1666464484
transform 1 0 49956 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_533
timestamp 1666464484
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_545
timestamp 1666464484
transform 1 0 51244 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_557
timestamp 1666464484
transform 1 0 52348 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_569
timestamp 1666464484
transform 1 0 53452 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_575
timestamp 1666464484
transform 1 0 54004 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_584
timestamp 1666464484
transform 1 0 54832 0 1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_102_589
timestamp 1666464484
transform 1 0 55292 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_601
timestamp 1666464484
transform 1 0 56396 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_613
timestamp 1666464484
transform 1 0 57500 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_102_623
timestamp 1666464484
transform 1 0 58420 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_3
timestamp 1666464484
transform 1 0 1380 0 -1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_103_11
timestamp 1666464484
transform 1 0 2116 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_23
timestamp 1666464484
transform 1 0 3220 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_35
timestamp 1666464484
transform 1 0 4324 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_47
timestamp 1666464484
transform 1 0 5428 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1666464484
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1666464484
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_69
timestamp 1666464484
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_81
timestamp 1666464484
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_93
timestamp 1666464484
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1666464484
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1666464484
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_113
timestamp 1666464484
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_125
timestamp 1666464484
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_137
timestamp 1666464484
transform 1 0 13708 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_103_147
timestamp 1666464484
transform 1 0 14628 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_103_157
timestamp 1666464484
transform 1 0 15548 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_103_165
timestamp 1666464484
transform 1 0 16284 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_103_169
timestamp 1666464484
transform 1 0 16652 0 -1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_103_180
timestamp 1666464484
transform 1 0 17664 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_192
timestamp 1666464484
transform 1 0 18768 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_204
timestamp 1666464484
transform 1 0 19872 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_216
timestamp 1666464484
transform 1 0 20976 0 -1 58752
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_103_225
timestamp 1666464484
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_237
timestamp 1666464484
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_249
timestamp 1666464484
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_261
timestamp 1666464484
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_273
timestamp 1666464484
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_279
timestamp 1666464484
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_281
timestamp 1666464484
transform 1 0 26956 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_293
timestamp 1666464484
transform 1 0 28060 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_305
timestamp 1666464484
transform 1 0 29164 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_317
timestamp 1666464484
transform 1 0 30268 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_329
timestamp 1666464484
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_335
timestamp 1666464484
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_337
timestamp 1666464484
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_349
timestamp 1666464484
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_361
timestamp 1666464484
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_373
timestamp 1666464484
transform 1 0 35420 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_385
timestamp 1666464484
transform 1 0 36524 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_391
timestamp 1666464484
transform 1 0 37076 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_393
timestamp 1666464484
transform 1 0 37260 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_405
timestamp 1666464484
transform 1 0 38364 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_425
timestamp 1666464484
transform 1 0 40204 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_437
timestamp 1666464484
transform 1 0 41308 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_103_445
timestamp 1666464484
transform 1 0 42044 0 -1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_103_449
timestamp 1666464484
transform 1 0 42412 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_461
timestamp 1666464484
transform 1 0 43516 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_473
timestamp 1666464484
transform 1 0 44620 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_485
timestamp 1666464484
transform 1 0 45724 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_497
timestamp 1666464484
transform 1 0 46828 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_503
timestamp 1666464484
transform 1 0 47380 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_505
timestamp 1666464484
transform 1 0 47564 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_517
timestamp 1666464484
transform 1 0 48668 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_529
timestamp 1666464484
transform 1 0 49772 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_541
timestamp 1666464484
transform 1 0 50876 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_553
timestamp 1666464484
transform 1 0 51980 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_559
timestamp 1666464484
transform 1 0 52532 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_561
timestamp 1666464484
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_573
timestamp 1666464484
transform 1 0 53820 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_585
timestamp 1666464484
transform 1 0 54924 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_597
timestamp 1666464484
transform 1 0 56028 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_609
timestamp 1666464484
transform 1 0 57132 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_615
timestamp 1666464484
transform 1 0 57684 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_103_617
timestamp 1666464484
transform 1 0 57868 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_623
timestamp 1666464484
transform 1 0 58420 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_104_3
timestamp 1666464484
transform 1 0 1380 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_9
timestamp 1666464484
transform 1 0 1932 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_21
timestamp 1666464484
transform 1 0 3036 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1666464484
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1666464484
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1666464484
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1666464484
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_65
timestamp 1666464484
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1666464484
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1666464484
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_85
timestamp 1666464484
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_97
timestamp 1666464484
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_109
timestamp 1666464484
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_121
timestamp 1666464484
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_133
timestamp 1666464484
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_139
timestamp 1666464484
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_141
timestamp 1666464484
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_153
timestamp 1666464484
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_165
timestamp 1666464484
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_177
timestamp 1666464484
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_189
timestamp 1666464484
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_195
timestamp 1666464484
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_197
timestamp 1666464484
transform 1 0 19228 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_209
timestamp 1666464484
transform 1 0 20332 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_221
timestamp 1666464484
transform 1 0 21436 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_233
timestamp 1666464484
transform 1 0 22540 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_245
timestamp 1666464484
transform 1 0 23644 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_251
timestamp 1666464484
transform 1 0 24196 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_253
timestamp 1666464484
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_265
timestamp 1666464484
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_277
timestamp 1666464484
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_289
timestamp 1666464484
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_301
timestamp 1666464484
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_307
timestamp 1666464484
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_309
timestamp 1666464484
transform 1 0 29532 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_321
timestamp 1666464484
transform 1 0 30636 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_333
timestamp 1666464484
transform 1 0 31740 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_345
timestamp 1666464484
transform 1 0 32844 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_357
timestamp 1666464484
transform 1 0 33948 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_363
timestamp 1666464484
transform 1 0 34500 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_365
timestamp 1666464484
transform 1 0 34684 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_377
timestamp 1666464484
transform 1 0 35788 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_389
timestamp 1666464484
transform 1 0 36892 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_401
timestamp 1666464484
transform 1 0 37996 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_413
timestamp 1666464484
transform 1 0 39100 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_419
timestamp 1666464484
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_421
timestamp 1666464484
transform 1 0 39836 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_433
timestamp 1666464484
transform 1 0 40940 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_445
timestamp 1666464484
transform 1 0 42044 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_104_457
timestamp 1666464484
transform 1 0 43148 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_104_474
timestamp 1666464484
transform 1 0 44712 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_477
timestamp 1666464484
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_489
timestamp 1666464484
transform 1 0 46092 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_501
timestamp 1666464484
transform 1 0 47196 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_513
timestamp 1666464484
transform 1 0 48300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_525
timestamp 1666464484
transform 1 0 49404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_531
timestamp 1666464484
transform 1 0 49956 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_533
timestamp 1666464484
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_545
timestamp 1666464484
transform 1 0 51244 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_557
timestamp 1666464484
transform 1 0 52348 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_569
timestamp 1666464484
transform 1 0 53452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_581
timestamp 1666464484
transform 1 0 54556 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_587
timestamp 1666464484
transform 1 0 55108 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_589
timestamp 1666464484
transform 1 0 55292 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_601
timestamp 1666464484
transform 1 0 56396 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_104_613
timestamp 1666464484
transform 1 0 57500 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_104_623
timestamp 1666464484
transform 1 0 58420 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_3
timestamp 1666464484
transform 1 0 1380 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_105_9
timestamp 1666464484
transform 1 0 1932 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_105_17
timestamp 1666464484
transform 1 0 2668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_29
timestamp 1666464484
transform 1 0 3772 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_41
timestamp 1666464484
transform 1 0 4876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_105_53
timestamp 1666464484
transform 1 0 5980 0 -1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_105_57
timestamp 1666464484
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_69
timestamp 1666464484
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_81
timestamp 1666464484
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_93
timestamp 1666464484
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1666464484
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1666464484
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_113
timestamp 1666464484
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_125
timestamp 1666464484
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_137
timestamp 1666464484
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_149
timestamp 1666464484
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_161
timestamp 1666464484
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_167
timestamp 1666464484
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_169
timestamp 1666464484
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_181
timestamp 1666464484
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_193
timestamp 1666464484
transform 1 0 18860 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_205
timestamp 1666464484
transform 1 0 19964 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_217
timestamp 1666464484
transform 1 0 21068 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_223
timestamp 1666464484
transform 1 0 21620 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_225
timestamp 1666464484
transform 1 0 21804 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_237
timestamp 1666464484
transform 1 0 22908 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_249
timestamp 1666464484
transform 1 0 24012 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_261
timestamp 1666464484
transform 1 0 25116 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_273
timestamp 1666464484
transform 1 0 26220 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_279
timestamp 1666464484
transform 1 0 26772 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_281
timestamp 1666464484
transform 1 0 26956 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_293
timestamp 1666464484
transform 1 0 28060 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_305
timestamp 1666464484
transform 1 0 29164 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_317
timestamp 1666464484
transform 1 0 30268 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_329
timestamp 1666464484
transform 1 0 31372 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_335
timestamp 1666464484
transform 1 0 31924 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_337
timestamp 1666464484
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_349
timestamp 1666464484
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_361
timestamp 1666464484
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_373
timestamp 1666464484
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_385
timestamp 1666464484
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_391
timestamp 1666464484
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_393
timestamp 1666464484
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_405
timestamp 1666464484
transform 1 0 38364 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_417
timestamp 1666464484
transform 1 0 39468 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_429
timestamp 1666464484
transform 1 0 40572 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_441
timestamp 1666464484
transform 1 0 41676 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_447
timestamp 1666464484
transform 1 0 42228 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_449
timestamp 1666464484
transform 1 0 42412 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_461
timestamp 1666464484
transform 1 0 43516 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_473
timestamp 1666464484
transform 1 0 44620 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_485
timestamp 1666464484
transform 1 0 45724 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_497
timestamp 1666464484
transform 1 0 46828 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_503
timestamp 1666464484
transform 1 0 47380 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_505
timestamp 1666464484
transform 1 0 47564 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_517
timestamp 1666464484
transform 1 0 48668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_529
timestamp 1666464484
transform 1 0 49772 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_541
timestamp 1666464484
transform 1 0 50876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_553
timestamp 1666464484
transform 1 0 51980 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_559
timestamp 1666464484
transform 1 0 52532 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_561
timestamp 1666464484
transform 1 0 52716 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_573
timestamp 1666464484
transform 1 0 53820 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_585
timestamp 1666464484
transform 1 0 54924 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_597
timestamp 1666464484
transform 1 0 56028 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_105_605
timestamp 1666464484
transform 1 0 56764 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_105_614
timestamp 1666464484
transform 1 0 57592 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_617
timestamp 1666464484
transform 1 0 57868 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_623
timestamp 1666464484
transform 1 0 58420 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_106_3
timestamp 1666464484
transform 1 0 1380 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_106_10
timestamp 1666464484
transform 1 0 2024 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_106_18
timestamp 1666464484
transform 1 0 2760 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_26
timestamp 1666464484
transform 1 0 3496 0 1 59840
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1666464484
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1666464484
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_53
timestamp 1666464484
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_65
timestamp 1666464484
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1666464484
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1666464484
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_85
timestamp 1666464484
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_97
timestamp 1666464484
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_109
timestamp 1666464484
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_121
timestamp 1666464484
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_133
timestamp 1666464484
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_139
timestamp 1666464484
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_141
timestamp 1666464484
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_153
timestamp 1666464484
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_165
timestamp 1666464484
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_177
timestamp 1666464484
transform 1 0 17388 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_189
timestamp 1666464484
transform 1 0 18492 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_195
timestamp 1666464484
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_197
timestamp 1666464484
transform 1 0 19228 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_209
timestamp 1666464484
transform 1 0 20332 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_221
timestamp 1666464484
transform 1 0 21436 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_233
timestamp 1666464484
transform 1 0 22540 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_245
timestamp 1666464484
transform 1 0 23644 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_251
timestamp 1666464484
transform 1 0 24196 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_253
timestamp 1666464484
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_265
timestamp 1666464484
transform 1 0 25484 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_277
timestamp 1666464484
transform 1 0 26588 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_289
timestamp 1666464484
transform 1 0 27692 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_301
timestamp 1666464484
transform 1 0 28796 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_307
timestamp 1666464484
transform 1 0 29348 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_309
timestamp 1666464484
transform 1 0 29532 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_321
timestamp 1666464484
transform 1 0 30636 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_333
timestamp 1666464484
transform 1 0 31740 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_345
timestamp 1666464484
transform 1 0 32844 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_357
timestamp 1666464484
transform 1 0 33948 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_363
timestamp 1666464484
transform 1 0 34500 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_365
timestamp 1666464484
transform 1 0 34684 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_377
timestamp 1666464484
transform 1 0 35788 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_389
timestamp 1666464484
transform 1 0 36892 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_401
timestamp 1666464484
transform 1 0 37996 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_413
timestamp 1666464484
transform 1 0 39100 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_419
timestamp 1666464484
transform 1 0 39652 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_421
timestamp 1666464484
transform 1 0 39836 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_433
timestamp 1666464484
transform 1 0 40940 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_445
timestamp 1666464484
transform 1 0 42044 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_457
timestamp 1666464484
transform 1 0 43148 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_469
timestamp 1666464484
transform 1 0 44252 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_475
timestamp 1666464484
transform 1 0 44804 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_477
timestamp 1666464484
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_489
timestamp 1666464484
transform 1 0 46092 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_501
timestamp 1666464484
transform 1 0 47196 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_513
timestamp 1666464484
transform 1 0 48300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_525
timestamp 1666464484
transform 1 0 49404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_531
timestamp 1666464484
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_533
timestamp 1666464484
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_545
timestamp 1666464484
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_557
timestamp 1666464484
transform 1 0 52348 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_569
timestamp 1666464484
transform 1 0 53452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_581
timestamp 1666464484
transform 1 0 54556 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_587
timestamp 1666464484
transform 1 0 55108 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_589
timestamp 1666464484
transform 1 0 55292 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_597
timestamp 1666464484
transform 1 0 56028 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_602
timestamp 1666464484
transform 1 0 56488 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_606
timestamp 1666464484
transform 1 0 56856 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_613
timestamp 1666464484
transform 1 0 57500 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_106_623
timestamp 1666464484
transform 1 0 58420 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_3
timestamp 1666464484
transform 1 0 1380 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_107_11
timestamp 1666464484
transform 1 0 2116 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_19
timestamp 1666464484
transform 1 0 2852 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_26
timestamp 1666464484
transform 1 0 3496 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_34
timestamp 1666464484
transform 1 0 4232 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_46
timestamp 1666464484
transform 1 0 5336 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_54
timestamp 1666464484
transform 1 0 6072 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1666464484
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_69
timestamp 1666464484
transform 1 0 7452 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_77
timestamp 1666464484
transform 1 0 8188 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_82
timestamp 1666464484
transform 1 0 8648 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_90
timestamp 1666464484
transform 1 0 9384 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_102
timestamp 1666464484
transform 1 0 10488 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_110
timestamp 1666464484
transform 1 0 11224 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_107_113
timestamp 1666464484
transform 1 0 11500 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_117
timestamp 1666464484
transform 1 0 11868 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_122
timestamp 1666464484
transform 1 0 12328 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_134
timestamp 1666464484
transform 1 0 13432 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_146
timestamp 1666464484
transform 1 0 14536 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_154
timestamp 1666464484
transform 1 0 15272 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_166
timestamp 1666464484
transform 1 0 16376 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_169
timestamp 1666464484
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_181
timestamp 1666464484
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_193
timestamp 1666464484
transform 1 0 18860 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_197
timestamp 1666464484
transform 1 0 19228 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_202
timestamp 1666464484
transform 1 0 19688 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_214
timestamp 1666464484
transform 1 0 20792 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_222
timestamp 1666464484
transform 1 0 21528 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_225
timestamp 1666464484
transform 1 0 21804 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_237
timestamp 1666464484
transform 1 0 22908 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_249
timestamp 1666464484
transform 1 0 24012 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_253
timestamp 1666464484
transform 1 0 24380 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_258
timestamp 1666464484
transform 1 0 24840 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_270
timestamp 1666464484
transform 1 0 25944 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_278
timestamp 1666464484
transform 1 0 26680 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_281
timestamp 1666464484
transform 1 0 26956 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_287
timestamp 1666464484
transform 1 0 27508 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_299
timestamp 1666464484
transform 1 0 28612 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_307
timestamp 1666464484
transform 1 0 29348 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_314
timestamp 1666464484
transform 1 0 29992 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_322
timestamp 1666464484
transform 1 0 30728 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_334
timestamp 1666464484
transform 1 0 31832 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_337
timestamp 1666464484
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_349
timestamp 1666464484
transform 1 0 33212 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_357
timestamp 1666464484
transform 1 0 33948 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_362
timestamp 1666464484
transform 1 0 34408 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_374
timestamp 1666464484
transform 1 0 35512 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_107_386
timestamp 1666464484
transform 1 0 36616 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_393
timestamp 1666464484
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_405
timestamp 1666464484
transform 1 0 38364 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_417
timestamp 1666464484
transform 1 0 39468 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_429
timestamp 1666464484
transform 1 0 40572 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_437
timestamp 1666464484
transform 1 0 41308 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_442
timestamp 1666464484
transform 1 0 41768 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_449
timestamp 1666464484
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_461
timestamp 1666464484
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_473
timestamp 1666464484
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_485
timestamp 1666464484
transform 1 0 45724 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_493
timestamp 1666464484
transform 1 0 46460 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_498
timestamp 1666464484
transform 1 0 46920 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_505
timestamp 1666464484
transform 1 0 47564 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_517
timestamp 1666464484
transform 1 0 48668 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_525
timestamp 1666464484
transform 1 0 49404 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_530
timestamp 1666464484
transform 1 0 49864 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_538
timestamp 1666464484
transform 1 0 50600 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_550
timestamp 1666464484
transform 1 0 51704 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_558
timestamp 1666464484
transform 1 0 52440 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_561
timestamp 1666464484
transform 1 0 52716 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_567
timestamp 1666464484
transform 1 0 53268 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_107_579
timestamp 1666464484
transform 1 0 54372 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_586
timestamp 1666464484
transform 1 0 55016 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_594
timestamp 1666464484
transform 1 0 55752 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_604
timestamp 1666464484
transform 1 0 56672 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_107_614
timestamp 1666464484
transform 1 0 57592 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_617
timestamp 1666464484
transform 1 0 57868 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_623
timestamp 1666464484
transform 1 0 58420 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_3
timestamp 1666464484
transform 1 0 1380 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_11
timestamp 1666464484
transform 1 0 2116 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_108_21
timestamp 1666464484
transform 1 0 3036 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1666464484
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_29
timestamp 1666464484
transform 1 0 3772 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_33
timestamp 1666464484
transform 1 0 4140 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_38
timestamp 1666464484
transform 1 0 4600 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_46
timestamp 1666464484
transform 1 0 5336 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_54
timestamp 1666464484
transform 1 0 6072 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_108_57
timestamp 1666464484
transform 1 0 6348 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_66
timestamp 1666464484
transform 1 0 7176 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_76
timestamp 1666464484
transform 1 0 8096 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_108_85
timestamp 1666464484
transform 1 0 8924 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_89
timestamp 1666464484
transform 1 0 9292 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_94
timestamp 1666464484
transform 1 0 9752 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_102
timestamp 1666464484
transform 1 0 10488 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_110
timestamp 1666464484
transform 1 0 11224 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_113
timestamp 1666464484
transform 1 0 11500 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_121
timestamp 1666464484
transform 1 0 12236 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_128
timestamp 1666464484
transform 1 0 12880 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_138
timestamp 1666464484
transform 1 0 13800 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_141
timestamp 1666464484
transform 1 0 14076 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_149
timestamp 1666464484
transform 1 0 14812 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_153
timestamp 1666464484
transform 1 0 15180 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_158
timestamp 1666464484
transform 1 0 15640 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_166
timestamp 1666464484
transform 1 0 16376 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_169
timestamp 1666464484
transform 1 0 16652 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_173
timestamp 1666464484
transform 1 0 17020 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_178
timestamp 1666464484
transform 1 0 17480 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_186
timestamp 1666464484
transform 1 0 18216 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_194
timestamp 1666464484
transform 1 0 18952 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_197
timestamp 1666464484
transform 1 0 19228 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_201
timestamp 1666464484
transform 1 0 19596 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_206
timestamp 1666464484
transform 1 0 20056 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_214
timestamp 1666464484
transform 1 0 20792 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_222
timestamp 1666464484
transform 1 0 21528 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_225
timestamp 1666464484
transform 1 0 21804 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_229
timestamp 1666464484
transform 1 0 22172 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_234
timestamp 1666464484
transform 1 0 22632 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_242
timestamp 1666464484
transform 1 0 23368 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_250
timestamp 1666464484
transform 1 0 24104 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_253
timestamp 1666464484
transform 1 0 24380 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_261
timestamp 1666464484
transform 1 0 25116 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_266
timestamp 1666464484
transform 1 0 25576 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_276
timestamp 1666464484
transform 1 0 26496 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_281
timestamp 1666464484
transform 1 0 26956 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_285
timestamp 1666464484
transform 1 0 27324 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_292
timestamp 1666464484
transform 1 0 27968 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_300
timestamp 1666464484
transform 1 0 28704 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_309
timestamp 1666464484
transform 1 0 29532 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_317
timestamp 1666464484
transform 1 0 30268 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_325
timestamp 1666464484
transform 1 0 31004 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_330
timestamp 1666464484
transform 1 0 31464 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_108_337
timestamp 1666464484
transform 1 0 32108 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_343
timestamp 1666464484
transform 1 0 32660 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_351
timestamp 1666464484
transform 1 0 33396 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_359
timestamp 1666464484
transform 1 0 34132 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_363
timestamp 1666464484
transform 1 0 34500 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_365
timestamp 1666464484
transform 1 0 34684 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_373
timestamp 1666464484
transform 1 0 35420 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_383
timestamp 1666464484
transform 1 0 36340 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_391
timestamp 1666464484
transform 1 0 37076 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_393
timestamp 1666464484
transform 1 0 37260 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_399
timestamp 1666464484
transform 1 0 37812 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_407
timestamp 1666464484
transform 1 0 38548 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_415
timestamp 1666464484
transform 1 0 39284 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_419
timestamp 1666464484
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_421
timestamp 1666464484
transform 1 0 39836 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_427
timestamp 1666464484
transform 1 0 40388 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_435
timestamp 1666464484
transform 1 0 41124 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_443
timestamp 1666464484
transform 1 0 41860 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_447
timestamp 1666464484
transform 1 0 42228 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_449
timestamp 1666464484
transform 1 0 42412 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_457
timestamp 1666464484
transform 1 0 43148 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_465
timestamp 1666464484
transform 1 0 43884 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_108_473
timestamp 1666464484
transform 1 0 44620 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_108_477
timestamp 1666464484
transform 1 0 44988 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_483
timestamp 1666464484
transform 1 0 45540 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_491
timestamp 1666464484
transform 1 0 46276 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_499
timestamp 1666464484
transform 1 0 47012 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_503
timestamp 1666464484
transform 1 0 47380 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_108_505
timestamp 1666464484
transform 1 0 47564 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_511
timestamp 1666464484
transform 1 0 48116 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_519
timestamp 1666464484
transform 1 0 48852 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_527
timestamp 1666464484
transform 1 0 49588 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_531
timestamp 1666464484
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_533
timestamp 1666464484
transform 1 0 50140 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_541
timestamp 1666464484
transform 1 0 50876 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_548
timestamp 1666464484
transform 1 0 51520 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_558
timestamp 1666464484
transform 1 0 52440 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_561
timestamp 1666464484
transform 1 0 52716 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_565
timestamp 1666464484
transform 1 0 53084 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_572
timestamp 1666464484
transform 1 0 53728 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_580
timestamp 1666464484
transform 1 0 54464 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_108_589
timestamp 1666464484
transform 1 0 55292 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_597
timestamp 1666464484
transform 1 0 56028 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_604
timestamp 1666464484
transform 1 0 56672 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_108_614
timestamp 1666464484
transform 1 0 57592 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_617
timestamp 1666464484
transform 1 0 57868 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_623
timestamp 1666464484
transform 1 0 58420 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666464484
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666464484
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666464484
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666464484
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666464484
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666464484
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666464484
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666464484
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666464484
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666464484
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666464484
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666464484
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666464484
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666464484
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666464484
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666464484
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666464484
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666464484
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666464484
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666464484
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666464484
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666464484
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666464484
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666464484
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666464484
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666464484
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666464484
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666464484
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666464484
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666464484
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666464484
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666464484
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666464484
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666464484
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666464484
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666464484
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1666464484
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1666464484
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1666464484
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1666464484
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1666464484
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1666464484
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1666464484
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1666464484
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1666464484
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1666464484
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1666464484
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1666464484
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1666464484
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1666464484
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1666464484
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1666464484
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1666464484
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1666464484
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1666464484
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1666464484
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1666464484
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1666464484
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1666464484
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1666464484
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1666464484
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1666464484
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1666464484
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1666464484
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1666464484
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1666464484
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1666464484
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1666464484
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1666464484
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1666464484
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1666464484
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1666464484
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1666464484
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1666464484
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1666464484
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1666464484
transform -1 0 58880 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1666464484
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1666464484
transform -1 0 58880 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1666464484
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1666464484
transform -1 0 58880 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1666464484
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1666464484
transform -1 0 58880 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1666464484
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1666464484
transform -1 0 58880 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1666464484
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1666464484
transform -1 0 58880 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1666464484
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1666464484
transform -1 0 58880 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666464484
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666464484
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666464484
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666464484
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666464484
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666464484
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666464484
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666464484
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666464484
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666464484
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666464484
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666464484
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666464484
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666464484
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666464484
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666464484
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666464484
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666464484
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666464484
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666464484
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666464484
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666464484
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666464484
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666464484
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666464484
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666464484
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666464484
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666464484
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666464484
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666464484
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666464484
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666464484
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666464484
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666464484
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666464484
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666464484
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666464484
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666464484
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666464484
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666464484
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666464484
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666464484
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666464484
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666464484
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666464484
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666464484
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666464484
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666464484
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666464484
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666464484
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666464484
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666464484
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666464484
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666464484
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666464484
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666464484
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666464484
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666464484
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666464484
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666464484
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666464484
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666464484
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666464484
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666464484
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666464484
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666464484
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666464484
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666464484
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666464484
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666464484
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666464484
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666464484
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666464484
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666464484
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666464484
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666464484
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666464484
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666464484
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666464484
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666464484
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666464484
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666464484
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666464484
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666464484
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666464484
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666464484
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666464484
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666464484
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666464484
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666464484
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666464484
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666464484
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666464484
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666464484
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666464484
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666464484
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666464484
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666464484
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666464484
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666464484
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666464484
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666464484
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666464484
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666464484
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666464484
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666464484
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666464484
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666464484
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666464484
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666464484
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666464484
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666464484
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666464484
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666464484
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666464484
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666464484
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666464484
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666464484
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666464484
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666464484
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666464484
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666464484
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666464484
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666464484
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666464484
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666464484
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666464484
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666464484
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666464484
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666464484
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666464484
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666464484
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666464484
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666464484
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666464484
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666464484
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666464484
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666464484
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666464484
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666464484
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666464484
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666464484
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666464484
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666464484
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666464484
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666464484
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666464484
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666464484
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666464484
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666464484
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666464484
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666464484
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666464484
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666464484
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666464484
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666464484
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666464484
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666464484
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666464484
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666464484
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666464484
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666464484
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666464484
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666464484
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666464484
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666464484
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666464484
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666464484
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666464484
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666464484
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666464484
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666464484
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666464484
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666464484
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666464484
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666464484
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666464484
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666464484
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666464484
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666464484
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666464484
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666464484
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666464484
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666464484
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666464484
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666464484
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666464484
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666464484
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1666464484
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1666464484
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1666464484
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1666464484
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1666464484
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1666464484
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1666464484
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1666464484
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1666464484
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1666464484
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1666464484
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1666464484
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1666464484
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1666464484
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1666464484
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1666464484
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1666464484
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1666464484
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1666464484
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1666464484
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1666464484
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1666464484
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1666464484
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1666464484
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1666464484
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1666464484
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1666464484
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1666464484
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1666464484
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1666464484
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1666464484
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1666464484
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1666464484
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1666464484
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1666464484
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1666464484
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1666464484
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1666464484
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1666464484
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1666464484
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1666464484
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1666464484
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1666464484
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1666464484
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1666464484
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1666464484
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1666464484
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1666464484
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1666464484
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1666464484
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1666464484
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1666464484
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1666464484
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1666464484
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1666464484
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1666464484
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1666464484
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1666464484
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1666464484
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1666464484
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1666464484
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1666464484
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1666464484
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1666464484
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1666464484
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1666464484
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1666464484
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1666464484
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1666464484
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1666464484
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1666464484
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1666464484
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1666464484
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1666464484
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1666464484
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1666464484
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1666464484
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1666464484
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1666464484
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1666464484
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1666464484
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1666464484
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1666464484
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1666464484
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1666464484
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1666464484
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1666464484
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1666464484
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1666464484
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1666464484
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1666464484
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1666464484
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1666464484
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1666464484
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1666464484
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1666464484
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1666464484
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1666464484
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1666464484
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1666464484
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1666464484
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1666464484
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1666464484
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1666464484
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1666464484
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1666464484
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1666464484
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1666464484
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1666464484
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1666464484
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1666464484
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1666464484
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1666464484
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1666464484
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1666464484
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1666464484
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1666464484
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1666464484
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1666464484
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1666464484
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1666464484
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1666464484
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1666464484
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1666464484
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1666464484
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1666464484
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1666464484
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1666464484
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1666464484
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1666464484
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1666464484
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1666464484
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1666464484
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1666464484
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1666464484
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1666464484
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1666464484
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1666464484
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1666464484
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1666464484
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1666464484
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1666464484
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1666464484
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1666464484
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1666464484
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1666464484
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1666464484
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1666464484
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1666464484
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1666464484
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1666464484
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1666464484
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1666464484
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1666464484
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1666464484
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1666464484
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1666464484
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1666464484
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1666464484
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1666464484
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1666464484
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1666464484
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1666464484
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1666464484
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1666464484
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1666464484
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1666464484
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1666464484
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1666464484
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1666464484
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1666464484
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1666464484
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1666464484
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1666464484
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1666464484
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1666464484
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1666464484
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1666464484
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1666464484
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1666464484
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1666464484
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1666464484
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1666464484
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1666464484
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1666464484
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1666464484
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1666464484
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1666464484
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1666464484
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1666464484
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1666464484
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1666464484
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1666464484
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1666464484
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1666464484
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1666464484
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1666464484
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1666464484
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1666464484
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1666464484
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1666464484
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1666464484
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1666464484
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1666464484
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1666464484
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1666464484
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1666464484
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1666464484
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1666464484
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1666464484
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1666464484
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1666464484
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1666464484
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1666464484
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1666464484
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1666464484
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1666464484
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1666464484
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1666464484
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1666464484
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1666464484
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1666464484
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1666464484
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1666464484
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1666464484
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1666464484
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1666464484
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1666464484
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1666464484
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1666464484
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1666464484
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1666464484
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1666464484
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1666464484
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1666464484
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1666464484
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1666464484
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1666464484
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1666464484
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1666464484
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1666464484
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1666464484
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1666464484
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1666464484
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1666464484
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1666464484
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1666464484
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1666464484
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1666464484
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1666464484
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1666464484
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1666464484
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1666464484
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1666464484
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1666464484
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1666464484
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1666464484
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1666464484
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1666464484
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1666464484
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1666464484
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1666464484
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1666464484
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1666464484
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1666464484
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1666464484
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1666464484
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1666464484
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1666464484
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1666464484
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1666464484
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1666464484
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1666464484
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1666464484
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1666464484
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1666464484
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1666464484
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1666464484
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1666464484
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1666464484
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1666464484
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1666464484
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1666464484
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1666464484
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1666464484
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1666464484
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1666464484
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1666464484
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1666464484
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1666464484
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1666464484
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1666464484
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1666464484
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1666464484
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1666464484
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1666464484
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1666464484
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1666464484
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1666464484
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1666464484
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1666464484
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1666464484
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1666464484
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1666464484
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1666464484
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1666464484
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1666464484
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1666464484
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1666464484
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1666464484
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1666464484
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1666464484
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1666464484
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1666464484
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1666464484
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1666464484
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1666464484
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1666464484
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1666464484
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1666464484
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1666464484
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1666464484
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1666464484
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1666464484
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1666464484
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1666464484
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1666464484
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1666464484
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1666464484
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1666464484
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1666464484
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1666464484
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1666464484
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1666464484
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1666464484
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1666464484
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1666464484
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1666464484
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1666464484
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1666464484
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1666464484
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1666464484
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1666464484
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1666464484
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1666464484
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1666464484
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1666464484
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1666464484
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1666464484
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1666464484
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1666464484
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1666464484
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1666464484
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1666464484
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1666464484
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1666464484
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1666464484
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1666464484
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1666464484
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1666464484
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1666464484
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1666464484
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1666464484
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1666464484
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1666464484
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1666464484
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1666464484
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1666464484
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1666464484
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1666464484
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1666464484
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1666464484
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1666464484
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1666464484
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1666464484
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1666464484
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1666464484
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1666464484
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1666464484
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1666464484
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1666464484
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1666464484
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1666464484
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1666464484
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1666464484
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1666464484
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1666464484
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1666464484
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1666464484
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1666464484
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1666464484
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1666464484
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1666464484
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1666464484
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1666464484
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1666464484
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1666464484
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1666464484
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1666464484
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1666464484
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1666464484
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1666464484
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1666464484
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1666464484
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1666464484
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1666464484
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1666464484
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1666464484
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1666464484
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1666464484
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1666464484
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1666464484
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1666464484
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1666464484
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1666464484
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1666464484
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1666464484
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1666464484
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1666464484
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1666464484
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1666464484
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1666464484
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1666464484
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1666464484
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1666464484
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1666464484
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1666464484
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1666464484
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1666464484
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1666464484
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1666464484
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1666464484
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1666464484
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1666464484
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1666464484
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1666464484
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1666464484
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1666464484
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1666464484
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1666464484
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1666464484
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1666464484
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1666464484
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1666464484
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1666464484
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1666464484
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1666464484
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1666464484
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1666464484
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1666464484
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1666464484
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1666464484
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1666464484
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1666464484
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1666464484
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1666464484
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1666464484
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1666464484
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1666464484
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1666464484
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1666464484
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1666464484
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1666464484
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1666464484
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1666464484
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1666464484
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1666464484
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1666464484
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1666464484
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1666464484
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1666464484
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1666464484
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1666464484
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1666464484
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1666464484
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1666464484
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1666464484
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1666464484
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1666464484
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1666464484
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1666464484
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1666464484
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1666464484
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1666464484
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1666464484
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1666464484
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1666464484
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1666464484
transform 1 0 6256 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1666464484
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1666464484
transform 1 0 11408 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1666464484
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1666464484
transform 1 0 16560 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1666464484
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1666464484
transform 1 0 21712 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1666464484
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1666464484
transform 1 0 26864 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1666464484
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1666464484
transform 1 0 32016 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1666464484
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1666464484
transform 1 0 37168 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1666464484
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1666464484
transform 1 0 42320 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1666464484
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1666464484
transform 1 0 47472 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1666464484
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1666464484
transform 1 0 52624 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1666464484
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1666464484
transform 1 0 57776 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0446_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1666464484
transform 1 0 23276 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0448_
timestamp 1666464484
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0449_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1666464484
transform 1 0 28244 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0451_
timestamp 1666464484
transform 1 0 30912 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0452_
timestamp 1666464484
transform 1 0 29624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0453_
timestamp 1666464484
transform 1 0 37536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0454_
timestamp 1666464484
transform 1 0 39652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0455_
timestamp 1666464484
transform 1 0 37168 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0456_
timestamp 1666464484
transform 1 0 42688 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0457_
timestamp 1666464484
transform 1 0 15640 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _0458_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19872 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor4b_2  _0459_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_4  _0460_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9108 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2b_1  _0461_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15824 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_4  _0462_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18032 0 -1 31552
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_1  _0463_
timestamp 1666464484
transform 1 0 2484 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18308 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_2  _0465_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16744 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_4  _0466_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0467_
timestamp 1666464484
transform 1 0 13524 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _0468_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18584 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0469_
timestamp 1666464484
transform 1 0 16008 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor4b_4  _0470_
timestamp 1666464484
transform 1 0 19412 0 1 29376
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_1  _0471_
timestamp 1666464484
transform 1 0 2024 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0472_
timestamp 1666464484
transform 1 0 17848 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0473_
timestamp 1666464484
transform 1 0 2484 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0474_
timestamp 1666464484
transform 1 0 18124 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0475_
timestamp 1666464484
transform 1 0 2484 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_4  _0476_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19688 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__or3_2  _0477_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 15824 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_2  _0478_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16928 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__nor4b_4  _0479_
timestamp 1666464484
transform 1 0 17204 0 1 31552
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_1  _0480_
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0481_
timestamp 1666464484
transform 1 0 17388 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0482_
timestamp 1666464484
transform 1 0 15548 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_4  _0483_
timestamp 1666464484
transform 1 0 17664 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0484_
timestamp 1666464484
transform 1 0 15180 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_4  _0485_
timestamp 1666464484
transform 1 0 17940 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_1  _0486_
timestamp 1666464484
transform 1 0 2484 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_2  _0487_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18032 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__nand2b_1  _0488_
timestamp 1666464484
transform 1 0 2484 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0489_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0490_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 38088 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0491_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17296 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0492_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17848 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _0493_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0494_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30820 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0495_
timestamp 1666464484
transform 1 0 28980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0496_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28428 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18308 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0498_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18768 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0499_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 12328 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_4  _0500_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 10580 0 1 16320
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_1  _0501_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16928 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _0502_
timestamp 1666464484
transform 1 0 17112 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0503_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0504_
timestamp 1666464484
transform 1 0 34868 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_2  _0505_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16836 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0506_
timestamp 1666464484
transform 1 0 15640 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _0507_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16928 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__nor4_4  _0508_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19412 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__a211o_2  _0509_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0510_
timestamp 1666464484
transform 1 0 35420 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0511_
timestamp 1666464484
transform 1 0 18676 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _0512_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0513_
timestamp 1666464484
transform 1 0 31740 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34316 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 53360 0 1 56576
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0516_
timestamp 1666464484
transform 1 0 33304 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0517_
timestamp 1666464484
transform 1 0 34408 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0518_
timestamp 1666464484
transform 1 0 34868 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0519_
timestamp 1666464484
transform 1 0 53820 0 -1 57664
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_1  _0520_
timestamp 1666464484
transform 1 0 32752 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0521_
timestamp 1666464484
transform 1 0 34960 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0522_
timestamp 1666464484
transform 1 0 32844 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _0523_
timestamp 1666464484
transform 1 0 33764 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_2  _0524_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19596 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _0525_
timestamp 1666464484
transform 1 0 21068 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _0526_
timestamp 1666464484
transform 1 0 33580 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0527_
timestamp 1666464484
transform 1 0 35788 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_4  _0528_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35236 0 -1 57664
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_4  _0529_
timestamp 1666464484
transform 1 0 14996 0 1 43520
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_1  _0530_
timestamp 1666464484
transform 1 0 33672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0531_
timestamp 1666464484
transform 1 0 34960 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0532_
timestamp 1666464484
transform 1 0 35696 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0533_
timestamp 1666464484
transform 1 0 54096 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0534_
timestamp 1666464484
transform 1 0 33580 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0535_
timestamp 1666464484
transform 1 0 15364 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _0536_
timestamp 1666464484
transform 1 0 34592 0 -1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_2  _0537_
timestamp 1666464484
transform 1 0 34868 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0538_
timestamp 1666464484
transform 1 0 45172 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0539_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 46184 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0540_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25484 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0541_
timestamp 1666464484
transform 1 0 14812 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _0542_
timestamp 1666464484
transform 1 0 15732 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__or3_4  _0543_
timestamp 1666464484
transform 1 0 26680 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0544_
timestamp 1666464484
transform 1 0 38088 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0545_
timestamp 1666464484
transform 1 0 38364 0 1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0546_
timestamp 1666464484
transform 1 0 22816 0 1 45696
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0547_
timestamp 1666464484
transform 1 0 16928 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0548_
timestamp 1666464484
transform 1 0 24012 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0549_
timestamp 1666464484
transform 1 0 23000 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0550_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23092 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _0551_
timestamp 1666464484
transform 1 0 25852 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0552_
timestamp 1666464484
transform 1 0 18676 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0553_
timestamp 1666464484
transform 1 0 19412 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0554_
timestamp 1666464484
transform 1 0 20700 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0555_
timestamp 1666464484
transform 1 0 20424 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0556_
timestamp 1666464484
transform 1 0 22724 0 1 57664
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0557_
timestamp 1666464484
transform 1 0 21344 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0558_
timestamp 1666464484
transform 1 0 39468 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0559_
timestamp 1666464484
transform 1 0 40112 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0560_
timestamp 1666464484
transform 1 0 11684 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0561_
timestamp 1666464484
transform 1 0 18216 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0562_
timestamp 1666464484
transform 1 0 2024 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0563_
timestamp 1666464484
transform 1 0 21160 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _0564_
timestamp 1666464484
transform 1 0 21988 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0565_
timestamp 1666464484
transform 1 0 20148 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0566_
timestamp 1666464484
transform 1 0 20792 0 1 57664
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0567_
timestamp 1666464484
transform 1 0 2116 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_4  _0568_
timestamp 1666464484
transform 1 0 1932 0 1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0569_
timestamp 1666464484
transform 1 0 21896 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_4  _0570_
timestamp 1666464484
transform 1 0 21988 0 -1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _0571_
timestamp 1666464484
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _0572_
timestamp 1666464484
transform 1 0 2024 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0573_
timestamp 1666464484
transform 1 0 22632 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0574_
timestamp 1666464484
transform 1 0 19688 0 -1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0575_
timestamp 1666464484
transform 1 0 25024 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0576_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23736 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor4b_4  _0577_
timestamp 1666464484
transform 1 0 23368 0 -1 34816
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0578_
timestamp 1666464484
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0579_
timestamp 1666464484
transform 1 0 22172 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_4  _0580_
timestamp 1666464484
transform 1 0 21528 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _0581_
timestamp 1666464484
transform 1 0 2484 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0582_
timestamp 1666464484
transform 1 0 20792 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0583_
timestamp 1666464484
transform 1 0 21160 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0584_
timestamp 1666464484
transform 1 0 21620 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0585_
timestamp 1666464484
transform 1 0 22080 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0586_
timestamp 1666464484
transform 1 0 22632 0 1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0587_
timestamp 1666464484
transform 1 0 20516 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0588_
timestamp 1666464484
transform 1 0 22908 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0589_
timestamp 1666464484
transform 1 0 21344 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0590_
timestamp 1666464484
transform 1 0 21988 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0591_
timestamp 1666464484
transform 1 0 22356 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_4  _0592_
timestamp 1666464484
transform 1 0 41860 0 1 3264
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _0593_
timestamp 1666464484
transform 1 0 3680 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0594_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 16560 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17020 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_4  _0596_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20976 0 1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__a211oi_4  _0597_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32476 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1666464484
transform 1 0 31556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0599_
timestamp 1666464484
transform 1 0 4416 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0600_
timestamp 1666464484
transform 1 0 22448 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_4  _0601_
timestamp 1666464484
transform 1 0 42596 0 -1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_1  _0602_
timestamp 1666464484
transform 1 0 22632 0 1 41344
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _0603_
timestamp 1666464484
transform 1 0 22908 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _0604_
timestamp 1666464484
transform 1 0 42872 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _0605_
timestamp 1666464484
transform 1 0 5152 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0606_
timestamp 1666464484
transform 1 0 24564 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0607_
timestamp 1666464484
transform 1 0 25392 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0608_
timestamp 1666464484
transform 1 0 24564 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _0609_
timestamp 1666464484
transform 1 0 24564 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0610_
timestamp 1666464484
transform 1 0 24840 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0611_
timestamp 1666464484
transform 1 0 24288 0 -1 35904
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_2  _0612_
timestamp 1666464484
transform 1 0 44712 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _0613_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0614_
timestamp 1666464484
transform 1 0 24748 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0615_
timestamp 1666464484
transform 1 0 24564 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0616_
timestamp 1666464484
transform 1 0 42596 0 -1 54400
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0617_
timestamp 1666464484
transform 1 0 43516 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_2  _0618_
timestamp 1666464484
transform 1 0 33304 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _0619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19964 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0620_
timestamp 1666464484
transform 1 0 43976 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0621_
timestamp 1666464484
transform 1 0 35788 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0622_
timestamp 1666464484
transform 1 0 37996 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0623_
timestamp 1666464484
transform 1 0 42964 0 -1 55488
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_2  _0624_
timestamp 1666464484
transform 1 0 43516 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_2  _0625_
timestamp 1666464484
transform 1 0 33212 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _0626_
timestamp 1666464484
transform 1 0 29440 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _0627_
timestamp 1666464484
transform 1 0 43148 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _0628_
timestamp 1666464484
transform 1 0 29716 0 1 30464
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0629_
timestamp 1666464484
transform 1 0 43424 0 1 56576
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_4  _0630_
timestamp 1666464484
transform 1 0 44068 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__a211o_4  _0631_
timestamp 1666464484
transform 1 0 29716 0 1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__a31o_2  _0632_
timestamp 1666464484
transform 1 0 19964 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0633_
timestamp 1666464484
transform 1 0 42228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0634_
timestamp 1666464484
transform 1 0 36892 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0635_
timestamp 1666464484
transform 1 0 37444 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_4  _0636_
timestamp 1666464484
transform 1 0 43424 0 1 57664
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_4  _0637_
timestamp 1666464484
transform 1 0 45172 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__a211o_2  _0638_
timestamp 1666464484
transform 1 0 32200 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_4  _0639_
timestamp 1666464484
transform 1 0 30268 0 -1 57664
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_2  _0640_
timestamp 1666464484
transform 1 0 45172 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0641_
timestamp 1666464484
transform 1 0 44804 0 -1 25024
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_4  _0642_
timestamp 1666464484
transform 1 0 31372 0 1 57664
box -38 -48 1602 592
use sky130_fd_sc_hd__a22o_1  _0643_
timestamp 1666464484
transform 1 0 45356 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _0644_
timestamp 1666464484
transform 1 0 45172 0 1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__a22o_4  _0645_
timestamp 1666464484
transform 1 0 43424 0 1 58752
box -38 -48 1326 592
use sky130_fd_sc_hd__a221o_4  _0646_
timestamp 1666464484
transform 1 0 44804 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__a211o_2  _0647_
timestamp 1666464484
transform 1 0 32752 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _0648_
timestamp 1666464484
transform 1 0 16836 0 1 23936
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_2  _0649_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20332 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0650_
timestamp 1666464484
transform 1 0 19872 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0651_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0652_
timestamp 1666464484
transform 1 0 28336 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0653_
timestamp 1666464484
transform 1 0 9384 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0654_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0655_
timestamp 1666464484
transform 1 0 9384 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0656_
timestamp 1666464484
transform 1 0 9660 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0657_
timestamp 1666464484
transform 1 0 14260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0658_
timestamp 1666464484
transform 1 0 18676 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0659_
timestamp 1666464484
transform 1 0 10120 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0660_
timestamp 1666464484
transform 1 0 10304 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0661_
timestamp 1666464484
transform 1 0 10672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0662_
timestamp 1666464484
transform 1 0 11592 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0663_
timestamp 1666464484
transform 1 0 12052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0664_
timestamp 1666464484
transform 1 0 10580 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0665_
timestamp 1666464484
transform 1 0 10672 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0666_
timestamp 1666464484
transform 1 0 11040 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0667_
timestamp 1666464484
transform 1 0 11684 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0668_
timestamp 1666464484
transform 1 0 11776 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0669_
timestamp 1666464484
transform 1 0 11592 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0670_
timestamp 1666464484
transform 1 0 11776 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0671_
timestamp 1666464484
transform 1 0 12788 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0672_
timestamp 1666464484
transform 1 0 12788 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0673_
timestamp 1666464484
transform 1 0 12420 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0674_
timestamp 1666464484
transform 1 0 12880 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0675_
timestamp 1666464484
transform 1 0 14260 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0676_
timestamp 1666464484
transform 1 0 32384 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0677_
timestamp 1666464484
transform 1 0 13984 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0678_
timestamp 1666464484
transform 1 0 14720 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0679_
timestamp 1666464484
transform 1 0 12788 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0680_
timestamp 1666464484
transform 1 0 12972 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0681_
timestamp 1666464484
transform 1 0 12972 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0682_
timestamp 1666464484
transform 1 0 13064 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0683_
timestamp 1666464484
transform 1 0 15824 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0684_
timestamp 1666464484
transform 1 0 23460 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0685_
timestamp 1666464484
transform 1 0 13248 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0686_
timestamp 1666464484
transform 1 0 24564 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0687_
timestamp 1666464484
transform 1 0 13616 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0688_
timestamp 1666464484
transform 1 0 23460 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0689_
timestamp 1666464484
transform 1 0 13248 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0690_
timestamp 1666464484
transform 1 0 25576 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0691_
timestamp 1666464484
transform 1 0 13984 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0692_
timestamp 1666464484
transform 1 0 23460 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0693_
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0694_
timestamp 1666464484
transform 1 0 14536 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0695_
timestamp 1666464484
transform 1 0 14720 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0696_
timestamp 1666464484
transform 1 0 22356 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0697_
timestamp 1666464484
transform 1 0 14904 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0698_
timestamp 1666464484
transform 1 0 14812 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0699_
timestamp 1666464484
transform 1 0 21712 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0700_
timestamp 1666464484
transform 1 0 24564 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0701_
timestamp 1666464484
transform 1 0 21528 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _0702_
timestamp 1666464484
transform 1 0 22448 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0703_
timestamp 1666464484
transform 1 0 14904 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0704_
timestamp 1666464484
transform 1 0 15088 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0705_
timestamp 1666464484
transform 1 0 10028 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0706_
timestamp 1666464484
transform 1 0 10764 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _0707_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 57040 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0708_
timestamp 1666464484
transform 1 0 57960 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_4  _0709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 37352 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0710_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30360 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0711_
timestamp 1666464484
transform 1 0 30268 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0712_
timestamp 1666464484
transform 1 0 36524 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0713_
timestamp 1666464484
transform 1 0 36340 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0714_
timestamp 1666464484
transform 1 0 24472 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0715_
timestamp 1666464484
transform 1 0 25576 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0716_
timestamp 1666464484
transform 1 0 28336 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0717_
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0718_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 55384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0719_
timestamp 1666464484
transform 1 0 23552 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0720_
timestamp 1666464484
transform 1 0 21988 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0721_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 37904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0722_
timestamp 1666464484
transform 1 0 38916 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0723_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 38824 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _0724_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 37996 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_1  _0725_
timestamp 1666464484
transform 1 0 29900 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0726_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30728 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0727_
timestamp 1666464484
transform 1 0 27968 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0728_
timestamp 1666464484
transform 1 0 27876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0729_
timestamp 1666464484
transform 1 0 28796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0730_
timestamp 1666464484
transform 1 0 28336 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0731_
timestamp 1666464484
transform 1 0 33948 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0732_
timestamp 1666464484
transform 1 0 34960 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0733_
timestamp 1666464484
transform 1 0 29256 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0734_
timestamp 1666464484
transform 1 0 27140 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0735_
timestamp 1666464484
transform 1 0 33764 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0736_
timestamp 1666464484
transform 1 0 33672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0737_
timestamp 1666464484
transform 1 0 32292 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0738_
timestamp 1666464484
transform 1 0 31188 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0739_
timestamp 1666464484
transform 1 0 32660 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0740_
timestamp 1666464484
transform 1 0 29716 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0741_
timestamp 1666464484
transform 1 0 27140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0742_
timestamp 1666464484
transform 1 0 25760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1666464484
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0744_
timestamp 1666464484
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0745_
timestamp 1666464484
transform 1 0 32292 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0746_
timestamp 1666464484
transform 1 0 27968 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0747_
timestamp 1666464484
transform 1 0 31372 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0748_
timestamp 1666464484
transform 1 0 29808 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0749_
timestamp 1666464484
transform 1 0 33764 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0750_
timestamp 1666464484
transform 1 0 35052 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0751_
timestamp 1666464484
transform 1 0 36432 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0752_
timestamp 1666464484
transform 1 0 36248 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0753_
timestamp 1666464484
transform 1 0 26404 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0754_
timestamp 1666464484
transform 1 0 25576 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0755_
timestamp 1666464484
transform 1 0 29256 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0756_
timestamp 1666464484
transform 1 0 31096 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0757_
timestamp 1666464484
transform 1 0 29716 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0758_
timestamp 1666464484
transform 1 0 27232 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0759_
timestamp 1666464484
transform 1 0 33764 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0760_
timestamp 1666464484
transform 1 0 35420 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0761_
timestamp 1666464484
transform 1 0 32384 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0762_
timestamp 1666464484
transform 1 0 35420 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0763_
timestamp 1666464484
transform 1 0 38824 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0764_
timestamp 1666464484
transform 1 0 38364 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0765_
timestamp 1666464484
transform 1 0 31372 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0766_
timestamp 1666464484
transform 1 0 32292 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0767_
timestamp 1666464484
transform 1 0 37352 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0768_
timestamp 1666464484
transform 1 0 37444 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0769_
timestamp 1666464484
transform 1 0 36524 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0770_
timestamp 1666464484
transform 1 0 36248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0771_
timestamp 1666464484
transform 1 0 28980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0772_
timestamp 1666464484
transform 1 0 29716 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0773_
timestamp 1666464484
transform 1 0 56028 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0774_
timestamp 1666464484
transform 1 0 38732 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0775_
timestamp 1666464484
transform 1 0 29256 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0776_
timestamp 1666464484
transform 1 0 24564 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0777_
timestamp 1666464484
transform 1 0 19504 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0778_
timestamp 1666464484
transform 1 0 19688 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0779_
timestamp 1666464484
transform 1 0 27140 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0780_
timestamp 1666464484
transform 1 0 22448 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0781_
timestamp 1666464484
transform 1 0 24564 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1666464484
transform 1 0 27140 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0783_
timestamp 1666464484
transform 1 0 19964 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0784_
timestamp 1666464484
transform 1 0 25852 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1666464484
transform 1 0 19412 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0786_
timestamp 1666464484
transform 1 0 29716 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0787_
timestamp 1666464484
transform 1 0 33764 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0788_
timestamp 1666464484
transform 1 0 36248 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1666464484
transform 1 0 28980 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0790_
timestamp 1666464484
transform 1 0 30820 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1666464484
transform 1 0 24564 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0792_
timestamp 1666464484
transform 1 0 34776 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1666464484
transform 1 0 34868 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0794_
timestamp 1666464484
transform 1 0 37812 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1666464484
transform 1 0 25760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0796_
timestamp 1666464484
transform 1 0 37628 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1666464484
transform 1 0 33580 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0798_
timestamp 1666464484
transform 1 0 20148 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0799_
timestamp 1666464484
transform 1 0 25576 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0800_
timestamp 1666464484
transform 1 0 25668 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1666464484
transform 1 0 21344 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0802_
timestamp 1666464484
transform 1 0 20148 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0803_
timestamp 1666464484
transform 1 0 18124 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0804_
timestamp 1666464484
transform 1 0 18124 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1666464484
transform 1 0 18400 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0806_
timestamp 1666464484
transform 1 0 17848 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0807_
timestamp 1666464484
transform 1 0 17848 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1666464484
transform 1 0 17848 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1666464484
transform 1 0 17296 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0810_
timestamp 1666464484
transform 1 0 17572 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0811_
timestamp 1666464484
transform 1 0 36984 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0812_
timestamp 1666464484
transform 1 0 40020 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 1666464484
transform 1 0 57316 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0814_
timestamp 1666464484
transform 1 0 32568 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0815_
timestamp 1666464484
transform 1 0 31648 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0816_
timestamp 1666464484
transform 1 0 30728 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0817_
timestamp 1666464484
transform 1 0 32568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _0818_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32936 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0819_
timestamp 1666464484
transform 1 0 58052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0820_
timestamp 1666464484
transform 1 0 55476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0821_
timestamp 1666464484
transform 1 0 29808 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0822_
timestamp 1666464484
transform 1 0 31188 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0823_
timestamp 1666464484
transform 1 0 33120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _0824_
timestamp 1666464484
transform 1 0 33580 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0825_
timestamp 1666464484
transform 1 0 56120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1666464484
transform 1 0 57316 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0827_
timestamp 1666464484
transform 1 0 30268 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0828_
timestamp 1666464484
transform 1 0 31004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0829_
timestamp 1666464484
transform 1 0 32292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _0830_
timestamp 1666464484
transform 1 0 31740 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0831_
timestamp 1666464484
transform 1 0 58052 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0832_
timestamp 1666464484
transform 1 0 34316 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0833_
timestamp 1666464484
transform 1 0 37812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0834_
timestamp 1666464484
transform 1 0 40020 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0835_
timestamp 1666464484
transform 1 0 41032 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0836_
timestamp 1666464484
transform 1 0 58052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_4  _0837_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27140 0 -1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__o221a_1  _0838_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29716 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_2  _0839_
timestamp 1666464484
transform 1 0 30544 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0840_
timestamp 1666464484
transform 1 0 56764 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0841_
timestamp 1666464484
transform 1 0 58052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0842_
timestamp 1666464484
transform 1 0 32292 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_2  _0843_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_2  _0844_
timestamp 1666464484
transform 1 0 31556 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0845_
timestamp 1666464484
transform 1 0 56764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_2  _0846_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29900 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_4  _0847_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 39744 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _0848_
timestamp 1666464484
transform 1 0 41032 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0849_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 40020 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0850_
timestamp 1666464484
transform 1 0 39008 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0851_
timestamp 1666464484
transform 1 0 29716 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0852_
timestamp 1666464484
transform 1 0 56672 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0853_
timestamp 1666464484
transform 1 0 56028 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0854_
timestamp 1666464484
transform 1 0 21988 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31648 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 41768 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0857_
timestamp 1666464484
transform 1 0 41768 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0858_
timestamp 1666464484
transform 1 0 24564 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0859_
timestamp 1666464484
transform 1 0 43792 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0860_
timestamp 1666464484
transform 1 0 42964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0861_
timestamp 1666464484
transform 1 0 31372 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _0862_
timestamp 1666464484
transform 1 0 28336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0863_
timestamp 1666464484
transform 1 0 49772 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0864_
timestamp 1666464484
transform 1 0 50048 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _0865_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30268 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__o2bb2a_1  _0866_
timestamp 1666464484
transform 1 0 43792 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0867_
timestamp 1666464484
transform 1 0 43792 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 36984 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0869_
timestamp 1666464484
transform 1 0 37444 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0870_
timestamp 1666464484
transform 1 0 38456 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0871_
timestamp 1666464484
transform 1 0 38180 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0872_
timestamp 1666464484
transform 1 0 28336 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1666464484
transform 1 0 37904 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0874_
timestamp 1666464484
transform 1 0 40020 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0875_
timestamp 1666464484
transform 1 0 38732 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0876_
timestamp 1666464484
transform 1 0 27048 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0877_
timestamp 1666464484
transform 1 0 27140 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0878_
timestamp 1666464484
transform 1 0 41952 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0879_
timestamp 1666464484
transform 1 0 41860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_4  _0880_
timestamp 1666464484
transform 1 0 27140 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__o2bb2a_1  _0881_
timestamp 1666464484
transform 1 0 43240 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0882_
timestamp 1666464484
transform 1 0 44436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0883_
timestamp 1666464484
transform 1 0 27692 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0884_
timestamp 1666464484
transform 1 0 55476 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0885_
timestamp 1666464484
transform 1 0 55844 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0886_
timestamp 1666464484
transform 1 0 34224 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_1  _0887_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 55936 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0888_
timestamp 1666464484
transform 1 0 56488 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0889_
timestamp 1666464484
transform 1 0 35236 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0890_
timestamp 1666464484
transform 1 0 50324 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1666464484
transform 1 0 50324 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _0892_
timestamp 1666464484
transform 1 0 35604 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_1  _0893_
timestamp 1666464484
transform 1 0 55936 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0894_
timestamp 1666464484
transform 1 0 56396 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0895_
timestamp 1666464484
transform 1 0 32292 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0896_
timestamp 1666464484
transform 1 0 56488 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0897_
timestamp 1666464484
transform 1 0 56672 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0898_
timestamp 1666464484
transform 1 0 30820 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_4  _0899_
timestamp 1666464484
transform 1 0 30268 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__o2bb2a_1  _0900_
timestamp 1666464484
transform 1 0 40388 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0901_
timestamp 1666464484
transform 1 0 40296 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0902_
timestamp 1666464484
transform 1 0 37444 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0903_
timestamp 1666464484
transform 1 0 47472 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0904_
timestamp 1666464484
transform 1 0 48484 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0905_
timestamp 1666464484
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0906_
timestamp 1666464484
transform 1 0 45172 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0907_
timestamp 1666464484
transform 1 0 43148 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0908_
timestamp 1666464484
transform 1 0 51428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0909_
timestamp 1666464484
transform 1 0 52900 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0910_
timestamp 1666464484
transform 1 0 51980 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0911_
timestamp 1666464484
transform 1 0 51980 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0912_
timestamp 1666464484
transform 1 0 58052 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 37720 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0914_
timestamp 1666464484
transform 1 0 56764 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0915_
timestamp 1666464484
transform 1 0 53728 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0916_
timestamp 1666464484
transform 1 0 54464 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0917_
timestamp 1666464484
transform 1 0 16928 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0918_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 18952 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0919_
timestamp 1666464484
transform 1 0 15548 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_2  _0920_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 19504 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0921_
timestamp 1666464484
transform 1 0 17572 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0922_
timestamp 1666464484
transform 1 0 17112 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1666464484
transform 1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0924_
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0925_
timestamp 1666464484
transform 1 0 15548 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0926_
timestamp 1666464484
transform 1 0 14996 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 21988 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0928_
timestamp 1666464484
transform 1 0 22632 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0929_
timestamp 1666464484
transform 1 0 18032 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0930_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 20148 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0931_
timestamp 1666464484
transform 1 0 19412 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0932_
timestamp 1666464484
transform 1 0 22632 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0933_
timestamp 1666464484
transform 1 0 21160 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0934_
timestamp 1666464484
transform 1 0 23644 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0935_
timestamp 1666464484
transform 1 0 24564 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0936_
timestamp 1666464484
transform 1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0937_
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0938_
timestamp 1666464484
transform 1 0 26128 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0939_
timestamp 1666464484
transform 1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _0940_
timestamp 1666464484
transform 1 0 23000 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0941_
timestamp 1666464484
transform 1 0 16652 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0942_
timestamp 1666464484
transform 1 0 17848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0943_
timestamp 1666464484
transform 1 0 21344 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0944_
timestamp 1666464484
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0945_
timestamp 1666464484
transform 1 0 17388 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0946_
timestamp 1666464484
transform 1 0 18308 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0947_
timestamp 1666464484
transform 1 0 19596 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0948_
timestamp 1666464484
transform 1 0 21160 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0949_
timestamp 1666464484
transform 1 0 24656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0950_
timestamp 1666464484
transform 1 0 22264 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0951_
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0952_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23000 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0953_
timestamp 1666464484
transform 1 0 22080 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and4_2  _0954_
timestamp 1666464484
transform 1 0 20424 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0955_
timestamp 1666464484
transform 1 0 19320 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0956_
timestamp 1666464484
transform 1 0 16100 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0957_
timestamp 1666464484
transform 1 0 15456 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0958_
timestamp 1666464484
transform 1 0 15732 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0959_
timestamp 1666464484
transform 1 0 16836 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4_2  _0960_
timestamp 1666464484
transform 1 0 18032 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0961_
timestamp 1666464484
transform 1 0 18124 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0962_
timestamp 1666464484
transform 1 0 20608 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0963_
timestamp 1666464484
transform 1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0964_
timestamp 1666464484
transform 1 0 18308 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0965_
timestamp 1666464484
transform 1 0 25208 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0966_
timestamp 1666464484
transform 1 0 27140 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0967_
timestamp 1666464484
transform 1 0 27140 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0968_
timestamp 1666464484
transform 1 0 20976 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0969_
timestamp 1666464484
transform 1 0 24564 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0970_
timestamp 1666464484
transform 1 0 32844 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0971_
timestamp 1666464484
transform 1 0 32660 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0972_
timestamp 1666464484
transform 1 0 21252 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0973_
timestamp 1666464484
transform 1 0 32292 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0974_
timestamp 1666464484
transform 1 0 32108 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30268 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0976_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 36432 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0977_
timestamp 1666464484
transform 1 0 23368 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0978_
timestamp 1666464484
transform 1 0 27692 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0979_
timestamp 1666464484
transform 1 0 20516 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0980_
timestamp 1666464484
transform 1 0 56028 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _0981_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30912 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0982_
timestamp 1666464484
transform 1 0 28060 0 -1 5440
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0983_
timestamp 1666464484
transform 1 0 28612 0 -1 6528
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0984_
timestamp 1666464484
transform 1 0 34868 0 1 7616
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _0985_
timestamp 1666464484
transform 1 0 27140 0 -1 10880
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _0986_
timestamp 1666464484
transform 1 0 32844 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0987_
timestamp 1666464484
transform 1 0 30268 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1666464484
transform 1 0 29808 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1666464484
transform 1 0 27140 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1666464484
transform 1 0 29900 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1666464484
transform 1 0 27784 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0992_
timestamp 1666464484
transform 1 0 32292 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0993_
timestamp 1666464484
transform 1 0 33672 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _0994_
timestamp 1666464484
transform 1 0 36524 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1666464484
transform 1 0 27140 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _0996_
timestamp 1666464484
transform 1 0 29992 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1666464484
transform 1 0 27692 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _0998_
timestamp 1666464484
transform 1 0 34868 0 1 21760
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _0999_
timestamp 1666464484
transform 1 0 35052 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1000_
timestamp 1666464484
transform 1 0 38732 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1001_
timestamp 1666464484
transform 1 0 31924 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1002_
timestamp 1666464484
transform 1 0 37628 0 1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1666464484
transform 1 0 36524 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1666464484
transform 1 0 29532 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1666464484
transform 1 0 56856 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1666464484
transform 1 0 28520 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1666464484
transform 1 0 23460 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1666464484
transform 1 0 19044 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1666464484
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1666464484
transform 1 0 25760 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1666464484
transform 1 0 21988 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1666464484
transform 1 0 23920 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1666464484
transform 1 0 26404 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1666464484
transform 1 0 19504 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1666464484
transform 1 0 24564 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1666464484
transform 1 0 19412 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1666464484
transform 1 0 27416 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1666464484
transform 1 0 32844 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1019_
timestamp 1666464484
transform 1 0 35420 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1666464484
transform 1 0 27324 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1666464484
transform 1 0 29716 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1666464484
transform 1 0 23644 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1666464484
transform 1 0 34868 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1666464484
transform 1 0 34684 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1666464484
transform 1 0 37444 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1666464484
transform 1 0 25116 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1027_
timestamp 1666464484
transform 1 0 35696 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1666464484
transform 1 0 33856 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1666464484
transform 1 0 19320 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1666464484
transform 1 0 24564 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1666464484
transform 1 0 24932 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1666464484
transform 1 0 20056 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1666464484
transform 1 0 19504 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1666464484
transform 1 0 19412 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1666464484
transform 1 0 19044 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1036_
timestamp 1666464484
transform 1 0 19044 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1037_
timestamp 1666464484
transform 1 0 19412 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1038_
timestamp 1666464484
transform 1 0 56856 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1039_
timestamp 1666464484
transform 1 0 56856 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1040_
timestamp 1666464484
transform 1 0 56856 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1041_
timestamp 1666464484
transform 1 0 40480 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1042_
timestamp 1666464484
transform 1 0 56856 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1043_
timestamp 1666464484
transform 1 0 56856 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1044_
timestamp 1666464484
transform 1 0 39468 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1045_
timestamp 1666464484
transform 1 0 56856 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1046_
timestamp 1666464484
transform 1 0 42596 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1047_
timestamp 1666464484
transform 1 0 43976 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1048_
timestamp 1666464484
transform 1 0 50324 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1049_
timestamp 1666464484
transform 1 0 43976 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1050_
timestamp 1666464484
transform 1 0 38916 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1051_
timestamp 1666464484
transform 1 0 39008 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1052_
timestamp 1666464484
transform 1 0 42596 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1053_
timestamp 1666464484
transform 1 0 43240 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1054_
timestamp 1666464484
transform 1 0 56028 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1055_
timestamp 1666464484
transform 1 0 56120 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1056_
timestamp 1666464484
transform 1 0 50324 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1057_
timestamp 1666464484
transform 1 0 56856 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1058_
timestamp 1666464484
transform 1 0 56856 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1059_
timestamp 1666464484
transform 1 0 40388 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1060_
timestamp 1666464484
transform 1 0 47748 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1061_
timestamp 1666464484
transform 1 0 44436 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1062_
timestamp 1666464484
transform 1 0 52532 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1063_
timestamp 1666464484
transform 1 0 52900 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1064_
timestamp 1666464484
transform 1 0 56856 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1065_
timestamp 1666464484
transform 1 0 53728 0 -1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1066_
timestamp 1666464484
transform 1 0 19596 0 1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1067_
timestamp 1666464484
transform 1 0 16836 0 -1 14144
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1068_
timestamp 1666464484
transform 1 0 14444 0 1 13056
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1069_
timestamp 1666464484
transform 1 0 14628 0 -1 15232
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1070_
timestamp 1666464484
transform 1 0 14628 0 -1 13056
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1071_
timestamp 1666464484
transform 1 0 21988 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1072_
timestamp 1666464484
transform 1 0 19964 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1666464484
transform 1 0 22448 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1666464484
transform 1 0 24564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1666464484
transform 1 0 22448 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1666464484
transform 1 0 22540 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1077_
timestamp 1666464484
transform 1 0 19412 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1078_
timestamp 1666464484
transform 1 0 17204 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1079_
timestamp 1666464484
transform 1 0 22356 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1666464484
transform 1 0 22448 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1081_
timestamp 1666464484
transform 1 0 22356 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1666464484
transform 1 0 19412 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1083_
timestamp 1666464484
transform 1 0 14444 0 1 20672
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _1084_
timestamp 1666464484
transform 1 0 15916 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1085_
timestamp 1666464484
transform 1 0 19780 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1086_
timestamp 1666464484
transform 1 0 22356 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1087_
timestamp 1666464484
transform 1 0 22172 0 -1 19584
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1666464484
transform 1 0 22632 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1666464484
transform 1 0 24564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1090_
timestamp 1666464484
transform 1 0 32752 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1666464484
transform 1 0 20056 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1092_
timestamp 1666464484
transform 1 0 32016 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_2  _1113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1114_
timestamp 1666464484
transform 1 0 31280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1115_
timestamp 1666464484
transform 1 0 32292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1116_
timestamp 1666464484
transform 1 0 33948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1117_
timestamp 1666464484
transform 1 0 33488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1118_
timestamp 1666464484
transform 1 0 34500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1119_
timestamp 1666464484
transform 1 0 34868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1120_
timestamp 1666464484
transform 1 0 35604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1121_
timestamp 1666464484
transform 1 0 38364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1666464484
transform 1 0 39192 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1123_
timestamp 1666464484
transform 1 0 39100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1666464484
transform 1 0 38088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1125_
timestamp 1666464484
transform 1 0 40020 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1126_
timestamp 1666464484
transform 1 0 37444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 38732 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1666464484
transform 1 0 23368 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1666464484
transform 1 0 29900 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1666464484
transform 1 0 27140 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1666464484
transform 1 0 32476 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1666464484
transform 1 0 46828 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1666464484
transform 1 0 49404 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1666464484
transform 1 0 41584 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1666464484
transform 1 0 46828 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout400 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 40020 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout401 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 40020 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout402
timestamp 1666464484
transform 1 0 33396 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout403
timestamp 1666464484
transform 1 0 39836 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout404
timestamp 1666464484
transform 1 0 39744 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout405
timestamp 1666464484
transform 1 0 47932 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout406
timestamp 1666464484
transform 1 0 57040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout407 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26956 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout408
timestamp 1666464484
transform 1 0 28152 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout409
timestamp 1666464484
transform 1 0 38180 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout410
timestamp 1666464484
transform 1 0 38272 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout411
timestamp 1666464484
transform 1 0 30820 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout412
timestamp 1666464484
transform 1 0 38824 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout413
timestamp 1666464484
transform 1 0 35420 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout414 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23552 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout415
timestamp 1666464484
transform 1 0 23552 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout416 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  fanout418
timestamp 1666464484
transform 1 0 19872 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  fanout419
timestamp 1666464484
transform 1 0 19688 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_12  fanout420 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 17940 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_8  fanout421 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 36708 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout422
timestamp 1666464484
transform 1 0 17296 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout423
timestamp 1666464484
transform 1 0 23000 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout424
timestamp 1666464484
transform 1 0 41308 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout425
timestamp 1666464484
transform 1 0 34592 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout426
timestamp 1666464484
transform 1 0 14260 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout427
timestamp 1666464484
transform 1 0 25024 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout428
timestamp 1666464484
transform 1 0 33856 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout429
timestamp 1666464484
transform 1 0 18124 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout430
timestamp 1666464484
transform 1 0 36340 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout431
timestamp 1666464484
transform 1 0 22908 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout432
timestamp 1666464484
transform 1 0 20424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_12  fanout433
timestamp 1666464484
transform 1 0 21988 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  fanout434
timestamp 1666464484
transform 1 0 17572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_12  fanout435
timestamp 1666464484
transform 1 0 22080 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_4  fanout436
timestamp 1666464484
transform 1 0 13800 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout437
timestamp 1666464484
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout438
timestamp 1666464484
transform 1 0 23000 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout439
timestamp 1666464484
transform 1 0 45356 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout440
timestamp 1666464484
transform 1 0 16008 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout441
timestamp 1666464484
transform 1 0 12604 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout442
timestamp 1666464484
transform 1 0 12144 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout443
timestamp 1666464484
transform 1 0 13248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout444
timestamp 1666464484
transform 1 0 14536 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout445
timestamp 1666464484
transform 1 0 18400 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout446
timestamp 1666464484
transform 1 0 17756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout447
timestamp 1666464484
transform 1 0 22632 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout448
timestamp 1666464484
transform 1 0 33488 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout449
timestamp 1666464484
transform 1 0 20148 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout450
timestamp 1666464484
transform 1 0 21528 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout451
timestamp 1666464484
transform 1 0 19596 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout452
timestamp 1666464484
transform 1 0 20148 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout453
timestamp 1666464484
transform 1 0 20516 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout454
timestamp 1666464484
transform 1 0 18308 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout455
timestamp 1666464484
transform 1 0 19412 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout456
timestamp 1666464484
transform 1 0 19228 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout457
timestamp 1666464484
transform 1 0 19412 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout458
timestamp 1666464484
transform 1 0 18124 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout459
timestamp 1666464484
transform 1 0 19412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout460
timestamp 1666464484
transform 1 0 19596 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout461
timestamp 1666464484
transform 1 0 37444 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout462
timestamp 1666464484
transform 1 0 36156 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout463
timestamp 1666464484
transform 1 0 37444 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout464
timestamp 1666464484
transform 1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout465
timestamp 1666464484
transform 1 0 39008 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout466
timestamp 1666464484
transform 1 0 39560 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout467
timestamp 1666464484
transform 1 0 40204 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout468
timestamp 1666464484
transform 1 0 32292 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout469
timestamp 1666464484
transform 1 0 38180 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout470
timestamp 1666464484
transform 1 0 37720 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout471
timestamp 1666464484
transform 1 0 33120 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout472
timestamp 1666464484
transform 1 0 29072 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout473
timestamp 1666464484
transform 1 0 54188 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout474
timestamp 1666464484
transform 1 0 56396 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  fanout475
timestamp 1666464484
transform 1 0 56764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout476
timestamp 1666464484
transform 1 0 56580 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__bufbuf_16  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26128 0 1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold2
timestamp 1666464484
transform 1 0 20240 0 1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold3
timestamp 1666464484
transform 1 0 28612 0 -1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold4
timestamp 1666464484
transform 1 0 21712 0 1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold5
timestamp 1666464484
transform 1 0 24288 0 -1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold6
timestamp 1666464484
transform 1 0 16560 0 1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold7
timestamp 1666464484
transform 1 0 26864 0 1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold8
timestamp 1666464484
transform 1 0 18400 0 -1 22848
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold9
timestamp 1666464484
transform 1 0 25576 0 1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold10
timestamp 1666464484
transform 1 0 15916 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold11
timestamp 1666464484
transform 1 0 31464 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold12
timestamp 1666464484
transform 1 0 24288 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold13
timestamp 1666464484
transform 1 0 26036 0 1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold14
timestamp 1666464484
transform 1 0 19136 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold15
timestamp 1666464484
transform 1 0 23092 0 -1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold16
timestamp 1666464484
transform 1 0 16560 0 1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold17
timestamp 1666464484
transform 1 0 26864 0 1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold18
timestamp 1666464484
transform 1 0 27140 0 -1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold19
timestamp 1666464484
transform 1 0 24564 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold20
timestamp 1666464484
transform 1 0 32292 0 -1 22848
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold21
timestamp 1666464484
transform 1 0 28612 0 -1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold22
timestamp 1666464484
transform 1 0 25300 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold23
timestamp 1666464484
transform 1 0 26680 0 1 22848
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold24
timestamp 1666464484
transform 1 0 24288 0 -1 22848
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold25
timestamp 1666464484
transform 1 0 21712 0 1 22848
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold26
timestamp 1666464484
transform 1 0 26220 0 1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold27
timestamp 1666464484
transform 1 0 22816 0 -1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold28
timestamp 1666464484
transform 1 0 21712 0 1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold29
timestamp 1666464484
transform 1 0 27140 0 -1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold30
timestamp 1666464484
transform 1 0 24288 0 -1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold31
timestamp 1666464484
transform 1 0 24288 0 -1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold32
timestamp 1666464484
transform 1 0 21712 0 1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold33
timestamp 1666464484
transform 1 0 15088 0 1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold34
timestamp 1666464484
transform 1 0 24288 0 -1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold35
timestamp 1666464484
transform 1 0 19780 0 1 17408
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold36
timestamp 1666464484
transform 1 0 19780 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold37
timestamp 1666464484
transform 1 0 26864 0 1 16320
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold38
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold39
timestamp 1666464484
transform 1 0 23368 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold40
timestamp 1666464484
transform 1 0 26404 0 1 23936
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold41
timestamp 1666464484
transform 1 0 21712 0 1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold42
timestamp 1666464484
transform 1 0 29440 0 -1 22848
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold43
timestamp 1666464484
transform 1 0 23552 0 -1 25024
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold44
timestamp 1666464484
transform 1 0 21712 0 1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold45
timestamp 1666464484
transform 1 0 23920 0 -1 23936
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold46
timestamp 1666464484
transform 1 0 19136 0 -1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold47
timestamp 1666464484
transform 1 0 19136 0 -1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold48
timestamp 1666464484
transform 1 0 28060 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold49
timestamp 1666464484
transform 1 0 21712 0 1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold50
timestamp 1666464484
transform 1 0 21068 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold51
timestamp 1666464484
transform 1 0 32292 0 -1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold52
timestamp 1666464484
transform 1 0 19136 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold53
timestamp 1666464484
transform 1 0 19136 0 -1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold54
timestamp 1666464484
transform 1 0 32292 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold55
timestamp 1666464484
transform 1 0 25208 0 1 18496
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold56
timestamp 1666464484
transform 1 0 24288 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold57
timestamp 1666464484
transform 1 0 24564 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold58
timestamp 1666464484
transform 1 0 17480 0 -1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold59
timestamp 1666464484
transform 1 0 16560 0 1 13056
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold60
timestamp 1666464484
transform 1 0 25576 0 1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold61
timestamp 1666464484
transform 1 0 16008 0 1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold62
timestamp 1666464484
transform 1 0 13984 0 -1 14144
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold63
timestamp 1666464484
transform 1 0 29716 0 1 15232
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold64
timestamp 1666464484
transform 1 0 31004 0 1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold65
timestamp 1666464484
transform 1 0 29440 0 -1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold66
timestamp 1666464484
transform 1 0 16560 0 1 21760
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold67
timestamp 1666464484
transform 1 0 31004 0 1 22848
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold68
timestamp 1666464484
transform 1 0 30360 0 1 20672
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold69
timestamp 1666464484
transform 1 0 34868 0 1 19584
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold70
timestamp 1666464484
transform 1 0 29256 0 -1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold71
timestamp 1666464484
transform 1 0 27140 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold72
timestamp 1666464484
transform 1 0 28336 0 -1 23936
box -38 -48 2430 592
use sky130_fd_sc_hd__bufbuf_16  hold73
timestamp 1666464484
transform 1 0 24288 0 -1 11968
box -38 -48 2430 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1666464484
transform 1 0 40572 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input2
timestamp 1666464484
transform 1 0 41584 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input3
timestamp 1666464484
transform 1 0 40940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1666464484
transform 1 0 42228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1666464484
transform 1 0 46000 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1666464484
transform 1 0 46276 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1666464484
transform 1 0 42964 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1666464484
transform 1 0 43884 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1666464484
transform 1 0 46736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1666464484
transform 1 0 43792 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1666464484
transform 1 0 44528 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1666464484
transform 1 0 39652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1666464484
transform 1 0 45172 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1666464484
transform 1 0 47104 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1666464484
transform 1 0 47748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1666464484
transform 1 0 45908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1666464484
transform 1 0 46736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1666464484
transform 1 0 47840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1666464484
transform 1 0 46644 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1666464484
transform 1 0 40756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input21
timestamp 1666464484
transform 1 0 40204 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1666464484
transform 1 0 40388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1666464484
transform 1 0 40940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input24
timestamp 1666464484
transform 1 0 41124 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1666464484
transform 1 0 41492 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input26
timestamp 1666464484
transform 1 0 42596 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input27
timestamp 1666464484
transform 1 0 42596 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1666464484
transform 1 0 54096 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1666464484
transform 1 0 54648 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1666464484
transform 1 0 55384 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1666464484
transform 1 0 56120 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1666464484
transform 1 0 58052 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 1666464484
transform 1 0 57040 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1666464484
transform 1 0 57040 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input35
timestamp 1666464484
transform 1 0 57040 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1666464484
transform 1 0 47748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input37
timestamp 1666464484
transform 1 0 50324 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input38
timestamp 1666464484
transform 1 0 49312 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1666464484
transform 1 0 50324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1666464484
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1666464484
transform 1 0 51796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input42
timestamp 1666464484
transform 1 0 51244 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1666464484
transform 1 0 51060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1666464484
transform 1 0 51796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input45
timestamp 1666464484
transform 1 0 52900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1666464484
transform 1 0 52900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1666464484
transform 1 0 47380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1666464484
transform 1 0 52532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1666464484
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input50
timestamp 1666464484
transform 1 0 53268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1666464484
transform 1 0 54372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1666464484
transform 1 0 55476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1666464484
transform 1 0 54004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1666464484
transform 1 0 55108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1666464484
transform 1 0 48576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1666464484
transform 1 0 48484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input57
timestamp 1666464484
transform 1 0 48116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input58
timestamp 1666464484
transform 1 0 47748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input59
timestamp 1666464484
transform 1 0 48668 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input60
timestamp 1666464484
transform 1 0 50324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input61
timestamp 1666464484
transform 1 0 48484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1666464484
transform 1 0 49404 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input63
timestamp 1666464484
transform 1 0 13248 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1666464484
transform 1 0 20424 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1666464484
transform 1 0 21160 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1666464484
transform 1 0 22264 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1666464484
transform 1 0 23000 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1666464484
transform 1 0 23736 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1666464484
transform 1 0 24472 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1666464484
transform 1 0 25208 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1666464484
transform 1 0 25944 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1666464484
transform 1 0 27140 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input73
timestamp 1666464484
transform 1 0 27416 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input74
timestamp 1666464484
transform 1 0 14260 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1666464484
transform 1 0 28336 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input76
timestamp 1666464484
transform 1 0 29716 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1666464484
transform 1 0 29624 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1666464484
transform 1 0 30360 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1666464484
transform 1 0 31096 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1666464484
transform 1 0 32292 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input81
timestamp 1666464484
transform 1 0 33028 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1666464484
transform 1 0 14904 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1666464484
transform 1 0 15272 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1666464484
transform 1 0 16008 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1666464484
transform 1 0 17112 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1666464484
transform 1 0 17848 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1666464484
transform 1 0 18584 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp 1666464484
transform 1 0 19320 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1666464484
transform 1 0 19688 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input90
timestamp 1666464484
transform 1 0 1564 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input91
timestamp 1666464484
transform 1 0 1564 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input92
timestamp 1666464484
transform 1 0 1564 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1666464484
transform 1 0 1564 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input94
timestamp 1666464484
transform 1 0 1564 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input95
timestamp 1666464484
transform 1 0 1564 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input96
timestamp 1666464484
transform 1 0 1564 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input97
timestamp 1666464484
transform 1 0 1564 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input98
timestamp 1666464484
transform 1 0 1564 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input99
timestamp 1666464484
transform 1 0 1564 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input100
timestamp 1666464484
transform 1 0 1564 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1666464484
transform 1 0 1564 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1666464484
transform 1 0 1564 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input103
timestamp 1666464484
transform 1 0 1564 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1666464484
transform 1 0 1564 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input105
timestamp 1666464484
transform 1 0 1564 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1666464484
transform 1 0 1564 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input107
timestamp 1666464484
transform 1 0 1564 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input108
timestamp 1666464484
transform 1 0 1564 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input109
timestamp 1666464484
transform 1 0 1564 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1666464484
transform 1 0 1564 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input111
timestamp 1666464484
transform 1 0 1564 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input112
timestamp 1666464484
transform 1 0 1564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input113
timestamp 1666464484
transform 1 0 1564 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input114
timestamp 1666464484
transform 1 0 1564 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1666464484
transform 1 0 1564 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1666464484
transform 1 0 1564 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input117
timestamp 1666464484
transform 1 0 1564 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input118
timestamp 1666464484
transform 1 0 33764 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1666464484
transform 1 0 41492 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input120
timestamp 1666464484
transform 1 0 41400 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input121
timestamp 1666464484
transform 1 0 42596 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input122
timestamp 1666464484
transform 1 0 43516 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input123
timestamp 1666464484
transform 1 0 44252 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input124
timestamp 1666464484
transform 1 0 45172 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input125
timestamp 1666464484
transform 1 0 45908 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input126
timestamp 1666464484
transform 1 0 46644 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input127
timestamp 1666464484
transform 1 0 46552 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input128
timestamp 1666464484
transform 1 0 47748 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input129
timestamp 1666464484
transform 1 0 34040 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1666464484
transform 1 0 48484 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input131
timestamp 1666464484
transform 1 0 49220 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input132
timestamp 1666464484
transform 1 0 49496 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input133
timestamp 1666464484
transform 1 0 50232 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input134
timestamp 1666464484
transform 1 0 50968 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input135
timestamp 1666464484
transform 1 0 51888 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input136
timestamp 1666464484
transform 1 0 52900 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input137
timestamp 1666464484
transform 1 0 34868 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input138
timestamp 1666464484
transform 1 0 35788 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input139
timestamp 1666464484
transform 1 0 36248 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input140
timestamp 1666464484
transform 1 0 37444 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input141
timestamp 1666464484
transform 1 0 38180 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input142
timestamp 1666464484
transform 1 0 38916 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input143
timestamp 1666464484
transform 1 0 40020 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input144
timestamp 1666464484
transform 1 0 40756 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input145
timestamp 1666464484
transform 1 0 58052 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input146
timestamp 1666464484
transform 1 0 56120 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input147
timestamp 1666464484
transform 1 0 56948 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input148
timestamp 1666464484
transform 1 0 58052 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input149
timestamp 1666464484
transform 1 0 58052 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input150
timestamp 1666464484
transform 1 0 58052 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input151
timestamp 1666464484
transform 1 0 58052 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input152
timestamp 1666464484
transform 1 0 58052 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input153
timestamp 1666464484
transform 1 0 57868 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input154
timestamp 1666464484
transform 1 0 57132 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input155
timestamp 1666464484
transform 1 0 56120 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input156
timestamp 1666464484
transform 1 0 57868 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input157
timestamp 1666464484
transform 1 0 6624 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input158
timestamp 1666464484
transform 1 0 7544 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input159
timestamp 1666464484
transform 1 0 8280 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input160
timestamp 1666464484
transform 1 0 9016 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input161
timestamp 1666464484
transform 1 0 9384 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input162
timestamp 1666464484
transform 1 0 10120 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input163
timestamp 1666464484
transform 1 0 10856 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input164
timestamp 1666464484
transform 1 0 11960 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input165
timestamp 1666464484
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input166
timestamp 1666464484
transform 1 0 1564 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input167
timestamp 1666464484
transform 1 0 1564 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input168
timestamp 1666464484
transform 1 0 1564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input169
timestamp 1666464484
transform 1 0 1564 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input170
timestamp 1666464484
transform 1 0 1564 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input171
timestamp 1666464484
transform 1 0 1564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input172
timestamp 1666464484
transform 1 0 1564 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input173
timestamp 1666464484
transform 1 0 1564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input174
timestamp 1666464484
transform 1 0 2300 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input175
timestamp 1666464484
transform 1 0 1656 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input176
timestamp 1666464484
transform 1 0 2392 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input177
timestamp 1666464484
transform 1 0 3128 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input178
timestamp 1666464484
transform 1 0 3864 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input179
timestamp 1666464484
transform 1 0 4232 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input180
timestamp 1666464484
transform 1 0 4968 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input181
timestamp 1666464484
transform 1 0 5704 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input182
timestamp 1666464484
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input183
timestamp 1666464484
transform 1 0 38824 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input184
timestamp 1666464484
transform 1 0 39836 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input185
timestamp 1666464484
transform 1 0 38916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input186
timestamp 1666464484
transform 1 0 2300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input187
timestamp 1666464484
transform 1 0 1564 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input188
timestamp 1666464484
transform 1 0 1564 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input189
timestamp 1666464484
transform 1 0 1564 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input190
timestamp 1666464484
transform 1 0 1564 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input191
timestamp 1666464484
transform 1 0 1564 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input192
timestamp 1666464484
transform 1 0 1564 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input193
timestamp 1666464484
transform 1 0 1564 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  input194
timestamp 1666464484
transform 1 0 54004 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  input195
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input196
timestamp 1666464484
transform 1 0 8280 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input197
timestamp 1666464484
transform 1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input198
timestamp 1666464484
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input199
timestamp 1666464484
transform 1 0 7912 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input200
timestamp 1666464484
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input201
timestamp 1666464484
transform 1 0 10120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input202
timestamp 1666464484
transform 1 0 8648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input203
timestamp 1666464484
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input204
timestamp 1666464484
transform 1 0 8280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input205
timestamp 1666464484
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input206
timestamp 1666464484
transform 1 0 10856 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input207
timestamp 1666464484
transform 1 0 11776 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input208
timestamp 1666464484
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input209
timestamp 1666464484
transform 1 0 8188 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input210
timestamp 1666464484
transform 1 0 12604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input211
timestamp 1666464484
transform 1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input212
timestamp 1666464484
transform 1 0 8924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input213
timestamp 1666464484
transform 1 0 13432 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input214
timestamp 1666464484
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input215
timestamp 1666464484
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input216
timestamp 1666464484
transform 1 0 14260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input217
timestamp 1666464484
transform 1 0 11776 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input218
timestamp 1666464484
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input219
timestamp 1666464484
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input220
timestamp 1666464484
transform 1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input221
timestamp 1666464484
transform 1 0 13248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input222
timestamp 1666464484
transform 1 0 15916 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input223
timestamp 1666464484
transform 1 0 13432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input224
timestamp 1666464484
transform 1 0 7360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input225
timestamp 1666464484
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input226
timestamp 1666464484
transform 1 0 7176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input227
timestamp 1666464484
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input228
timestamp 1666464484
transform 1 0 6808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input229
timestamp 1666464484
transform 1 0 40020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input230
timestamp 1666464484
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input231
timestamp 1666464484
transform 1 0 12328 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input232
timestamp 1666464484
transform 1 0 2484 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input233
timestamp 1666464484
transform 1 0 53176 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input234
timestamp 1666464484
transform 1 0 1564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input235
timestamp 1666464484
transform 1 0 56304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input236
timestamp 1666464484
transform 1 0 57868 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input237
timestamp 1666464484
transform 1 0 58052 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input238
timestamp 1666464484
transform 1 0 57868 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input239
timestamp 1666464484
transform 1 0 58052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input240
timestamp 1666464484
transform 1 0 58052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input241
timestamp 1666464484
transform 1 0 57040 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input242
timestamp 1666464484
transform 1 0 58052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input243
timestamp 1666464484
transform 1 0 58052 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input244
timestamp 1666464484
transform 1 0 58052 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input245
timestamp 1666464484
transform 1 0 57868 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input246
timestamp 1666464484
transform 1 0 56948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input247
timestamp 1666464484
transform 1 0 57868 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input248
timestamp 1666464484
transform 1 0 56948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input249
timestamp 1666464484
transform 1 0 57868 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input250
timestamp 1666464484
transform 1 0 57868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input251
timestamp 1666464484
transform 1 0 57868 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input252
timestamp 1666464484
transform 1 0 57868 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input253
timestamp 1666464484
transform 1 0 56948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input254
timestamp 1666464484
transform 1 0 57868 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input255
timestamp 1666464484
transform 1 0 56948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input256
timestamp 1666464484
transform 1 0 57868 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input257
timestamp 1666464484
transform 1 0 57868 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input258
timestamp 1666464484
transform 1 0 57868 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input259
timestamp 1666464484
transform 1 0 57868 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input260
timestamp 1666464484
transform 1 0 56120 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input261
timestamp 1666464484
transform 1 0 56948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input262
timestamp 1666464484
transform 1 0 57040 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input263
timestamp 1666464484
transform 1 0 57868 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input264
timestamp 1666464484
transform 1 0 57868 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input265
timestamp 1666464484
transform 1 0 57868 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input266
timestamp 1666464484
transform 1 0 56948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input267
timestamp 1666464484
transform 1 0 56948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input268
timestamp 1666464484
transform 1 0 58052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input269
timestamp 1666464484
transform 1 0 58052 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  max_cap417
timestamp 1666464484
transform 1 0 19780 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  multiplexer_477 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_478
timestamp 1666464484
transform 1 0 26404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_479
timestamp 1666464484
transform 1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_480
timestamp 1666464484
transform 1 0 25484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_481
timestamp 1666464484
transform 1 0 17480 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_482
timestamp 1666464484
transform 1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_483
timestamp 1666464484
transform 1 0 17572 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_484
timestamp 1666464484
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_485
timestamp 1666464484
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_486
timestamp 1666464484
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_487
timestamp 1666464484
transform 1 0 58144 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_488
timestamp 1666464484
transform 1 0 58144 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_489
timestamp 1666464484
transform 1 0 58144 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_490
timestamp 1666464484
transform 1 0 58144 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_491
timestamp 1666464484
transform 1 0 27048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_492
timestamp 1666464484
transform 1 0 27692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_493
timestamp 1666464484
transform 1 0 28980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_494
timestamp 1666464484
transform 1 0 28336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_495
timestamp 1666464484
transform 1 0 27692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  multiplexer_496
timestamp 1666464484
transform 1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output270
timestamp 1666464484
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output271
timestamp 1666464484
transform 1 0 1564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output272
timestamp 1666464484
transform 1 0 1564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output273
timestamp 1666464484
transform 1 0 1564 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output274
timestamp 1666464484
transform 1 0 1564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output275
timestamp 1666464484
transform 1 0 1564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output276
timestamp 1666464484
transform 1 0 1564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output277
timestamp 1666464484
transform 1 0 1564 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output278
timestamp 1666464484
transform 1 0 1564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output279
timestamp 1666464484
transform 1 0 1564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output280
timestamp 1666464484
transform 1 0 1564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output281
timestamp 1666464484
transform 1 0 1564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output282
timestamp 1666464484
transform 1 0 1564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output283
timestamp 1666464484
transform 1 0 1564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output284
timestamp 1666464484
transform 1 0 1564 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output285
timestamp 1666464484
transform 1 0 1564 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output286
timestamp 1666464484
transform 1 0 1564 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output287
timestamp 1666464484
transform 1 0 1564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output288
timestamp 1666464484
transform 1 0 1564 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output289
timestamp 1666464484
transform 1 0 1564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output290
timestamp 1666464484
transform 1 0 1564 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output291
timestamp 1666464484
transform 1 0 1564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output292
timestamp 1666464484
transform 1 0 1564 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output293
timestamp 1666464484
transform 1 0 1564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output294
timestamp 1666464484
transform 1 0 1564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output295
timestamp 1666464484
transform 1 0 1564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output296
timestamp 1666464484
transform 1 0 1564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output297
timestamp 1666464484
transform 1 0 1564 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output298
timestamp 1666464484
transform 1 0 1564 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output299
timestamp 1666464484
transform 1 0 27140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output300
timestamp 1666464484
transform 1 0 28704 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output301
timestamp 1666464484
transform 1 0 30268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output302
timestamp 1666464484
transform 1 0 30176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output303
timestamp 1666464484
transform 1 0 30820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output304
timestamp 1666464484
transform 1 0 31096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output305
timestamp 1666464484
transform 1 0 32292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output306
timestamp 1666464484
transform 1 0 32292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output307
timestamp 1666464484
transform 1 0 33212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output308
timestamp 1666464484
transform 1 0 33212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output309
timestamp 1666464484
transform 1 0 34132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output310
timestamp 1666464484
transform 1 0 34868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output311
timestamp 1666464484
transform 1 0 35052 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output312
timestamp 1666464484
transform 1 0 35788 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output313
timestamp 1666464484
transform 1 0 34868 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output314
timestamp 1666464484
transform 1 0 35972 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output315
timestamp 1666464484
transform 1 0 35788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output316
timestamp 1666464484
transform 1 0 37444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output317
timestamp 1666464484
transform 1 0 34868 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output318
timestamp 1666464484
transform 1 0 36708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output319
timestamp 1666464484
transform 1 0 37444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output320
timestamp 1666464484
transform 1 0 38364 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output321
timestamp 1666464484
transform 1 0 38364 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output322
timestamp 1666464484
transform 1 0 36064 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output323
timestamp 1666464484
transform 1 0 37444 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output324
timestamp 1666464484
transform 1 0 39284 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output325
timestamp 1666464484
transform 1 0 40020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output326
timestamp 1666464484
transform 1 0 37168 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output327
timestamp 1666464484
transform 1 0 13984 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output328
timestamp 1666464484
transform 1 0 16836 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output329
timestamp 1666464484
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output330
timestamp 1666464484
transform 1 0 16560 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output331
timestamp 1666464484
transform 1 0 15824 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output332
timestamp 1666464484
transform 1 0 15824 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output333
timestamp 1666464484
transform 1 0 17480 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output334
timestamp 1666464484
transform 1 0 17204 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output335
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output336
timestamp 1666464484
transform 1 0 20976 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output337
timestamp 1666464484
transform 1 0 15824 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output338
timestamp 1666464484
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output339
timestamp 1666464484
transform 1 0 18124 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output340
timestamp 1666464484
transform 1 0 22540 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output341
timestamp 1666464484
transform 1 0 18400 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output342
timestamp 1666464484
transform 1 0 20976 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output343
timestamp 1666464484
transform 1 0 22448 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output344
timestamp 1666464484
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output345
timestamp 1666464484
transform 1 0 20976 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output346
timestamp 1666464484
transform 1 0 20976 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output347
timestamp 1666464484
transform 1 0 22540 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output348
timestamp 1666464484
transform 1 0 17020 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output349
timestamp 1666464484
transform 1 0 23552 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output350
timestamp 1666464484
transform 1 0 22632 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output351
timestamp 1666464484
transform 1 0 23552 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output352
timestamp 1666464484
transform 1 0 25760 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output353
timestamp 1666464484
transform 1 0 25208 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output354
timestamp 1666464484
transform 1 0 26128 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output355
timestamp 1666464484
transform 1 0 27140 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output356
timestamp 1666464484
transform 1 0 26128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output357
timestamp 1666464484
transform 1 0 15640 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output358
timestamp 1666464484
transform 1 0 14904 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output359
timestamp 1666464484
transform 1 0 1564 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output360
timestamp 1666464484
transform 1 0 1564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output361
timestamp 1666464484
transform 1 0 1564 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output362
timestamp 1666464484
transform 1 0 1564 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output363
timestamp 1666464484
transform 1 0 1564 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output364
timestamp 1666464484
transform 1 0 1564 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output365
timestamp 1666464484
transform 1 0 1564 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output366
timestamp 1666464484
transform 1 0 1564 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output367
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output368
timestamp 1666464484
transform 1 0 1564 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output369
timestamp 1666464484
transform 1 0 1564 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output370
timestamp 1666464484
transform 1 0 1564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output371
timestamp 1666464484
transform 1 0 57040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output372
timestamp 1666464484
transform 1 0 56948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output373
timestamp 1666464484
transform 1 0 57868 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output374
timestamp 1666464484
transform 1 0 57868 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output375
timestamp 1666464484
transform 1 0 57868 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output376
timestamp 1666464484
transform 1 0 57868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output377
timestamp 1666464484
transform 1 0 57868 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output378
timestamp 1666464484
transform 1 0 57868 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output379
timestamp 1666464484
transform 1 0 57868 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output380
timestamp 1666464484
transform 1 0 57868 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output381
timestamp 1666464484
transform 1 0 57868 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output382
timestamp 1666464484
transform 1 0 57868 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output383
timestamp 1666464484
transform 1 0 56120 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output384
timestamp 1666464484
transform 1 0 56948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output385
timestamp 1666464484
transform 1 0 57868 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output386
timestamp 1666464484
transform 1 0 56948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output387
timestamp 1666464484
transform 1 0 57868 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output388
timestamp 1666464484
transform 1 0 56948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output389
timestamp 1666464484
transform 1 0 57868 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output390
timestamp 1666464484
transform 1 0 56948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output391
timestamp 1666464484
transform 1 0 57868 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output392
timestamp 1666464484
transform 1 0 57040 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output393
timestamp 1666464484
transform 1 0 57868 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output394
timestamp 1666464484
transform 1 0 56948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output395
timestamp 1666464484
transform 1 0 57040 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output396
timestamp 1666464484
transform 1 0 56948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output397
timestamp 1666464484
transform 1 0 57040 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output398
timestamp 1666464484
transform 1 0 57868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output399
timestamp 1666464484
transform 1 0 57868 0 1 19584
box -38 -48 590 592
<< labels >>
flabel metal3 s 0 21360 800 21480 0 FreeSans 480 0 0 0 design_clk_o
port 0 nsew signal tristate
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 dsi_all[0]
port 1 nsew signal tristate
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 dsi_all[10]
port 2 nsew signal tristate
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 dsi_all[11]
port 3 nsew signal tristate
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 dsi_all[12]
port 4 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 dsi_all[13]
port 5 nsew signal tristate
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 dsi_all[14]
port 6 nsew signal tristate
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 dsi_all[15]
port 7 nsew signal tristate
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 dsi_all[16]
port 8 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 dsi_all[17]
port 9 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 dsi_all[18]
port 10 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 dsi_all[19]
port 11 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 dsi_all[1]
port 12 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 dsi_all[20]
port 13 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 dsi_all[21]
port 14 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 dsi_all[22]
port 15 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 dsi_all[23]
port 16 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 dsi_all[24]
port 17 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 dsi_all[25]
port 18 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 dsi_all[26]
port 19 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 dsi_all[27]
port 20 nsew signal tristate
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 dsi_all[2]
port 21 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 dsi_all[3]
port 22 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 dsi_all[4]
port 23 nsew signal tristate
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 dsi_all[5]
port 24 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 dsi_all[6]
port 25 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 dsi_all[7]
port 26 nsew signal tristate
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 dsi_all[8]
port 27 nsew signal tristate
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 dsi_all[9]
port 28 nsew signal tristate
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 dso_6502[0]
port 29 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 dso_6502[10]
port 30 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 dso_6502[11]
port 31 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 dso_6502[12]
port 32 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 dso_6502[13]
port 33 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 dso_6502[14]
port 34 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 dso_6502[15]
port 35 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 dso_6502[16]
port 36 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 dso_6502[17]
port 37 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 dso_6502[18]
port 38 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 dso_6502[19]
port 39 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 dso_6502[1]
port 40 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 dso_6502[20]
port 41 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 dso_6502[21]
port 42 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 dso_6502[22]
port 43 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 dso_6502[23]
port 44 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 dso_6502[24]
port 45 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 dso_6502[25]
port 46 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 dso_6502[26]
port 47 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 dso_6502[2]
port 48 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 dso_6502[3]
port 49 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 dso_6502[4]
port 50 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 dso_6502[5]
port 51 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 dso_6502[6]
port 52 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 dso_6502[7]
port 53 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 dso_6502[8]
port 54 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 dso_6502[9]
port 55 nsew signal input
flabel metal2 s 53838 63200 53894 64000 0 FreeSans 224 90 0 0 dso_LCD[0]
port 56 nsew signal input
flabel metal2 s 54574 63200 54630 64000 0 FreeSans 224 90 0 0 dso_LCD[1]
port 57 nsew signal input
flabel metal2 s 55310 63200 55366 64000 0 FreeSans 224 90 0 0 dso_LCD[2]
port 58 nsew signal input
flabel metal2 s 56046 63200 56102 64000 0 FreeSans 224 90 0 0 dso_LCD[3]
port 59 nsew signal input
flabel metal2 s 56782 63200 56838 64000 0 FreeSans 224 90 0 0 dso_LCD[4]
port 60 nsew signal input
flabel metal2 s 57518 63200 57574 64000 0 FreeSans 224 90 0 0 dso_LCD[5]
port 61 nsew signal input
flabel metal2 s 58254 63200 58310 64000 0 FreeSans 224 90 0 0 dso_LCD[6]
port 62 nsew signal input
flabel metal2 s 58990 63200 59046 64000 0 FreeSans 224 90 0 0 dso_LCD[7]
port 63 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 dso_as1802[0]
port 64 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 dso_as1802[10]
port 65 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 dso_as1802[11]
port 66 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 dso_as1802[12]
port 67 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 dso_as1802[13]
port 68 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 dso_as1802[14]
port 69 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 dso_as1802[15]
port 70 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 dso_as1802[16]
port 71 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 dso_as1802[17]
port 72 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 dso_as1802[18]
port 73 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 dso_as1802[19]
port 74 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 dso_as1802[1]
port 75 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 dso_as1802[20]
port 76 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 dso_as1802[21]
port 77 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 dso_as1802[22]
port 78 nsew signal input
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 dso_as1802[23]
port 79 nsew signal input
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 dso_as1802[24]
port 80 nsew signal input
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 dso_as1802[25]
port 81 nsew signal input
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 dso_as1802[26]
port 82 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 dso_as1802[2]
port 83 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 dso_as1802[3]
port 84 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 dso_as1802[4]
port 85 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 dso_as1802[5]
port 86 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 dso_as1802[6]
port 87 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 dso_as1802[7]
port 88 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 dso_as1802[8]
port 89 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 dso_as1802[9]
port 90 nsew signal input
flabel metal2 s 13358 63200 13414 64000 0 FreeSans 224 90 0 0 dso_as2650[0]
port 91 nsew signal input
flabel metal2 s 20718 63200 20774 64000 0 FreeSans 224 90 0 0 dso_as2650[10]
port 92 nsew signal input
flabel metal2 s 21454 63200 21510 64000 0 FreeSans 224 90 0 0 dso_as2650[11]
port 93 nsew signal input
flabel metal2 s 22190 63200 22246 64000 0 FreeSans 224 90 0 0 dso_as2650[12]
port 94 nsew signal input
flabel metal2 s 22926 63200 22982 64000 0 FreeSans 224 90 0 0 dso_as2650[13]
port 95 nsew signal input
flabel metal2 s 23662 63200 23718 64000 0 FreeSans 224 90 0 0 dso_as2650[14]
port 96 nsew signal input
flabel metal2 s 24398 63200 24454 64000 0 FreeSans 224 90 0 0 dso_as2650[15]
port 97 nsew signal input
flabel metal2 s 25134 63200 25190 64000 0 FreeSans 224 90 0 0 dso_as2650[16]
port 98 nsew signal input
flabel metal2 s 25870 63200 25926 64000 0 FreeSans 224 90 0 0 dso_as2650[17]
port 99 nsew signal input
flabel metal2 s 26606 63200 26662 64000 0 FreeSans 224 90 0 0 dso_as2650[18]
port 100 nsew signal input
flabel metal2 s 27342 63200 27398 64000 0 FreeSans 224 90 0 0 dso_as2650[19]
port 101 nsew signal input
flabel metal2 s 14094 63200 14150 64000 0 FreeSans 224 90 0 0 dso_as2650[1]
port 102 nsew signal input
flabel metal2 s 28078 63200 28134 64000 0 FreeSans 224 90 0 0 dso_as2650[20]
port 103 nsew signal input
flabel metal2 s 28814 63200 28870 64000 0 FreeSans 224 90 0 0 dso_as2650[21]
port 104 nsew signal input
flabel metal2 s 29550 63200 29606 64000 0 FreeSans 224 90 0 0 dso_as2650[22]
port 105 nsew signal input
flabel metal2 s 30286 63200 30342 64000 0 FreeSans 224 90 0 0 dso_as2650[23]
port 106 nsew signal input
flabel metal2 s 31022 63200 31078 64000 0 FreeSans 224 90 0 0 dso_as2650[24]
port 107 nsew signal input
flabel metal2 s 31758 63200 31814 64000 0 FreeSans 224 90 0 0 dso_as2650[25]
port 108 nsew signal input
flabel metal2 s 32494 63200 32550 64000 0 FreeSans 224 90 0 0 dso_as2650[26]
port 109 nsew signal input
flabel metal2 s 14830 63200 14886 64000 0 FreeSans 224 90 0 0 dso_as2650[2]
port 110 nsew signal input
flabel metal2 s 15566 63200 15622 64000 0 FreeSans 224 90 0 0 dso_as2650[3]
port 111 nsew signal input
flabel metal2 s 16302 63200 16358 64000 0 FreeSans 224 90 0 0 dso_as2650[4]
port 112 nsew signal input
flabel metal2 s 17038 63200 17094 64000 0 FreeSans 224 90 0 0 dso_as2650[5]
port 113 nsew signal input
flabel metal2 s 17774 63200 17830 64000 0 FreeSans 224 90 0 0 dso_as2650[6]
port 114 nsew signal input
flabel metal2 s 18510 63200 18566 64000 0 FreeSans 224 90 0 0 dso_as2650[7]
port 115 nsew signal input
flabel metal2 s 19246 63200 19302 64000 0 FreeSans 224 90 0 0 dso_as2650[8]
port 116 nsew signal input
flabel metal2 s 19982 63200 20038 64000 0 FreeSans 224 90 0 0 dso_as2650[9]
port 117 nsew signal input
flabel metal3 s 0 42440 800 42560 0 FreeSans 480 0 0 0 dso_as512512512[0]
port 118 nsew signal input
flabel metal3 s 0 49240 800 49360 0 FreeSans 480 0 0 0 dso_as512512512[10]
port 119 nsew signal input
flabel metal3 s 0 49920 800 50040 0 FreeSans 480 0 0 0 dso_as512512512[11]
port 120 nsew signal input
flabel metal3 s 0 50600 800 50720 0 FreeSans 480 0 0 0 dso_as512512512[12]
port 121 nsew signal input
flabel metal3 s 0 51280 800 51400 0 FreeSans 480 0 0 0 dso_as512512512[13]
port 122 nsew signal input
flabel metal3 s 0 51960 800 52080 0 FreeSans 480 0 0 0 dso_as512512512[14]
port 123 nsew signal input
flabel metal3 s 0 52640 800 52760 0 FreeSans 480 0 0 0 dso_as512512512[15]
port 124 nsew signal input
flabel metal3 s 0 53320 800 53440 0 FreeSans 480 0 0 0 dso_as512512512[16]
port 125 nsew signal input
flabel metal3 s 0 54000 800 54120 0 FreeSans 480 0 0 0 dso_as512512512[17]
port 126 nsew signal input
flabel metal3 s 0 54680 800 54800 0 FreeSans 480 0 0 0 dso_as512512512[18]
port 127 nsew signal input
flabel metal3 s 0 55360 800 55480 0 FreeSans 480 0 0 0 dso_as512512512[19]
port 128 nsew signal input
flabel metal3 s 0 43120 800 43240 0 FreeSans 480 0 0 0 dso_as512512512[1]
port 129 nsew signal input
flabel metal3 s 0 56040 800 56160 0 FreeSans 480 0 0 0 dso_as512512512[20]
port 130 nsew signal input
flabel metal3 s 0 56720 800 56840 0 FreeSans 480 0 0 0 dso_as512512512[21]
port 131 nsew signal input
flabel metal3 s 0 57400 800 57520 0 FreeSans 480 0 0 0 dso_as512512512[22]
port 132 nsew signal input
flabel metal3 s 0 58080 800 58200 0 FreeSans 480 0 0 0 dso_as512512512[23]
port 133 nsew signal input
flabel metal3 s 0 58760 800 58880 0 FreeSans 480 0 0 0 dso_as512512512[24]
port 134 nsew signal input
flabel metal3 s 0 59440 800 59560 0 FreeSans 480 0 0 0 dso_as512512512[25]
port 135 nsew signal input
flabel metal3 s 0 60120 800 60240 0 FreeSans 480 0 0 0 dso_as512512512[26]
port 136 nsew signal input
flabel metal3 s 0 60800 800 60920 0 FreeSans 480 0 0 0 dso_as512512512[27]
port 137 nsew signal input
flabel metal3 s 0 43800 800 43920 0 FreeSans 480 0 0 0 dso_as512512512[2]
port 138 nsew signal input
flabel metal3 s 0 44480 800 44600 0 FreeSans 480 0 0 0 dso_as512512512[3]
port 139 nsew signal input
flabel metal3 s 0 45160 800 45280 0 FreeSans 480 0 0 0 dso_as512512512[4]
port 140 nsew signal input
flabel metal3 s 0 45840 800 45960 0 FreeSans 480 0 0 0 dso_as512512512[5]
port 141 nsew signal input
flabel metal3 s 0 46520 800 46640 0 FreeSans 480 0 0 0 dso_as512512512[6]
port 142 nsew signal input
flabel metal3 s 0 47200 800 47320 0 FreeSans 480 0 0 0 dso_as512512512[7]
port 143 nsew signal input
flabel metal3 s 0 47880 800 48000 0 FreeSans 480 0 0 0 dso_as512512512[8]
port 144 nsew signal input
flabel metal3 s 0 48560 800 48680 0 FreeSans 480 0 0 0 dso_as512512512[9]
port 145 nsew signal input
flabel metal2 s 33230 63200 33286 64000 0 FreeSans 224 90 0 0 dso_as5401[0]
port 146 nsew signal input
flabel metal2 s 40590 63200 40646 64000 0 FreeSans 224 90 0 0 dso_as5401[10]
port 147 nsew signal input
flabel metal2 s 41326 63200 41382 64000 0 FreeSans 224 90 0 0 dso_as5401[11]
port 148 nsew signal input
flabel metal2 s 42062 63200 42118 64000 0 FreeSans 224 90 0 0 dso_as5401[12]
port 149 nsew signal input
flabel metal2 s 42798 63200 42854 64000 0 FreeSans 224 90 0 0 dso_as5401[13]
port 150 nsew signal input
flabel metal2 s 43534 63200 43590 64000 0 FreeSans 224 90 0 0 dso_as5401[14]
port 151 nsew signal input
flabel metal2 s 44270 63200 44326 64000 0 FreeSans 224 90 0 0 dso_as5401[15]
port 152 nsew signal input
flabel metal2 s 45006 63200 45062 64000 0 FreeSans 224 90 0 0 dso_as5401[16]
port 153 nsew signal input
flabel metal2 s 45742 63200 45798 64000 0 FreeSans 224 90 0 0 dso_as5401[17]
port 154 nsew signal input
flabel metal2 s 46478 63200 46534 64000 0 FreeSans 224 90 0 0 dso_as5401[18]
port 155 nsew signal input
flabel metal2 s 47214 63200 47270 64000 0 FreeSans 224 90 0 0 dso_as5401[19]
port 156 nsew signal input
flabel metal2 s 33966 63200 34022 64000 0 FreeSans 224 90 0 0 dso_as5401[1]
port 157 nsew signal input
flabel metal2 s 47950 63200 48006 64000 0 FreeSans 224 90 0 0 dso_as5401[20]
port 158 nsew signal input
flabel metal2 s 48686 63200 48742 64000 0 FreeSans 224 90 0 0 dso_as5401[21]
port 159 nsew signal input
flabel metal2 s 49422 63200 49478 64000 0 FreeSans 224 90 0 0 dso_as5401[22]
port 160 nsew signal input
flabel metal2 s 50158 63200 50214 64000 0 FreeSans 224 90 0 0 dso_as5401[23]
port 161 nsew signal input
flabel metal2 s 50894 63200 50950 64000 0 FreeSans 224 90 0 0 dso_as5401[24]
port 162 nsew signal input
flabel metal2 s 51630 63200 51686 64000 0 FreeSans 224 90 0 0 dso_as5401[25]
port 163 nsew signal input
flabel metal2 s 52366 63200 52422 64000 0 FreeSans 224 90 0 0 dso_as5401[26]
port 164 nsew signal input
flabel metal2 s 34702 63200 34758 64000 0 FreeSans 224 90 0 0 dso_as5401[2]
port 165 nsew signal input
flabel metal2 s 35438 63200 35494 64000 0 FreeSans 224 90 0 0 dso_as5401[3]
port 166 nsew signal input
flabel metal2 s 36174 63200 36230 64000 0 FreeSans 224 90 0 0 dso_as5401[4]
port 167 nsew signal input
flabel metal2 s 36910 63200 36966 64000 0 FreeSans 224 90 0 0 dso_as5401[5]
port 168 nsew signal input
flabel metal2 s 37646 63200 37702 64000 0 FreeSans 224 90 0 0 dso_as5401[6]
port 169 nsew signal input
flabel metal2 s 38382 63200 38438 64000 0 FreeSans 224 90 0 0 dso_as5401[7]
port 170 nsew signal input
flabel metal2 s 39118 63200 39174 64000 0 FreeSans 224 90 0 0 dso_as5401[8]
port 171 nsew signal input
flabel metal2 s 39854 63200 39910 64000 0 FreeSans 224 90 0 0 dso_as5401[9]
port 172 nsew signal input
flabel metal3 s 59200 56584 60000 56704 0 FreeSans 480 0 0 0 dso_counter[0]
port 173 nsew signal input
flabel metal3 s 59200 62024 60000 62144 0 FreeSans 480 0 0 0 dso_counter[10]
port 174 nsew signal input
flabel metal3 s 59200 62568 60000 62688 0 FreeSans 480 0 0 0 dso_counter[11]
port 175 nsew signal input
flabel metal3 s 59200 57128 60000 57248 0 FreeSans 480 0 0 0 dso_counter[1]
port 176 nsew signal input
flabel metal3 s 59200 57672 60000 57792 0 FreeSans 480 0 0 0 dso_counter[2]
port 177 nsew signal input
flabel metal3 s 59200 58216 60000 58336 0 FreeSans 480 0 0 0 dso_counter[3]
port 178 nsew signal input
flabel metal3 s 59200 58760 60000 58880 0 FreeSans 480 0 0 0 dso_counter[4]
port 179 nsew signal input
flabel metal3 s 59200 59304 60000 59424 0 FreeSans 480 0 0 0 dso_counter[5]
port 180 nsew signal input
flabel metal3 s 59200 59848 60000 59968 0 FreeSans 480 0 0 0 dso_counter[6]
port 181 nsew signal input
flabel metal3 s 59200 60392 60000 60512 0 FreeSans 480 0 0 0 dso_counter[7]
port 182 nsew signal input
flabel metal3 s 59200 60936 60000 61056 0 FreeSans 480 0 0 0 dso_counter[8]
port 183 nsew signal input
flabel metal3 s 59200 61480 60000 61600 0 FreeSans 480 0 0 0 dso_counter[9]
port 184 nsew signal input
flabel metal2 s 6734 63200 6790 64000 0 FreeSans 224 90 0 0 dso_diceroll[0]
port 185 nsew signal input
flabel metal2 s 7470 63200 7526 64000 0 FreeSans 224 90 0 0 dso_diceroll[1]
port 186 nsew signal input
flabel metal2 s 8206 63200 8262 64000 0 FreeSans 224 90 0 0 dso_diceroll[2]
port 187 nsew signal input
flabel metal2 s 8942 63200 8998 64000 0 FreeSans 224 90 0 0 dso_diceroll[3]
port 188 nsew signal input
flabel metal2 s 9678 63200 9734 64000 0 FreeSans 224 90 0 0 dso_diceroll[4]
port 189 nsew signal input
flabel metal2 s 10414 63200 10470 64000 0 FreeSans 224 90 0 0 dso_diceroll[5]
port 190 nsew signal input
flabel metal2 s 11150 63200 11206 64000 0 FreeSans 224 90 0 0 dso_diceroll[6]
port 191 nsew signal input
flabel metal2 s 11886 63200 11942 64000 0 FreeSans 224 90 0 0 dso_diceroll[7]
port 192 nsew signal input
flabel metal3 s 0 30200 800 30320 0 FreeSans 480 0 0 0 dso_mc14500[0]
port 193 nsew signal input
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 dso_mc14500[1]
port 194 nsew signal input
flabel metal3 s 0 31560 800 31680 0 FreeSans 480 0 0 0 dso_mc14500[2]
port 195 nsew signal input
flabel metal3 s 0 32240 800 32360 0 FreeSans 480 0 0 0 dso_mc14500[3]
port 196 nsew signal input
flabel metal3 s 0 32920 800 33040 0 FreeSans 480 0 0 0 dso_mc14500[4]
port 197 nsew signal input
flabel metal3 s 0 33600 800 33720 0 FreeSans 480 0 0 0 dso_mc14500[5]
port 198 nsew signal input
flabel metal3 s 0 34280 800 34400 0 FreeSans 480 0 0 0 dso_mc14500[6]
port 199 nsew signal input
flabel metal3 s 0 34960 800 35080 0 FreeSans 480 0 0 0 dso_mc14500[7]
port 200 nsew signal input
flabel metal3 s 0 35640 800 35760 0 FreeSans 480 0 0 0 dso_mc14500[8]
port 201 nsew signal input
flabel metal2 s 846 63200 902 64000 0 FreeSans 224 90 0 0 dso_multiplier[0]
port 202 nsew signal input
flabel metal2 s 1582 63200 1638 64000 0 FreeSans 224 90 0 0 dso_multiplier[1]
port 203 nsew signal input
flabel metal2 s 2318 63200 2374 64000 0 FreeSans 224 90 0 0 dso_multiplier[2]
port 204 nsew signal input
flabel metal2 s 3054 63200 3110 64000 0 FreeSans 224 90 0 0 dso_multiplier[3]
port 205 nsew signal input
flabel metal2 s 3790 63200 3846 64000 0 FreeSans 224 90 0 0 dso_multiplier[4]
port 206 nsew signal input
flabel metal2 s 4526 63200 4582 64000 0 FreeSans 224 90 0 0 dso_multiplier[5]
port 207 nsew signal input
flabel metal2 s 5262 63200 5318 64000 0 FreeSans 224 90 0 0 dso_multiplier[6]
port 208 nsew signal input
flabel metal2 s 5998 63200 6054 64000 0 FreeSans 224 90 0 0 dso_multiplier[7]
port 209 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 dso_posit[0]
port 210 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 dso_posit[1]
port 211 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 dso_posit[2]
port 212 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 dso_posit[3]
port 213 nsew signal input
flabel metal3 s 0 37000 800 37120 0 FreeSans 480 0 0 0 dso_tbb1143[0]
port 214 nsew signal input
flabel metal3 s 0 37680 800 37800 0 FreeSans 480 0 0 0 dso_tbb1143[1]
port 215 nsew signal input
flabel metal3 s 0 38360 800 38480 0 FreeSans 480 0 0 0 dso_tbb1143[2]
port 216 nsew signal input
flabel metal3 s 0 39040 800 39160 0 FreeSans 480 0 0 0 dso_tbb1143[3]
port 217 nsew signal input
flabel metal3 s 0 39720 800 39840 0 FreeSans 480 0 0 0 dso_tbb1143[4]
port 218 nsew signal input
flabel metal3 s 0 40400 800 40520 0 FreeSans 480 0 0 0 dso_tbb1143[5]
port 219 nsew signal input
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 dso_tbb1143[6]
port 220 nsew signal input
flabel metal3 s 0 41760 800 41880 0 FreeSans 480 0 0 0 dso_tbb1143[7]
port 221 nsew signal input
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 dso_tune
port 222 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 io_in[0]
port 223 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 io_in[10]
port 224 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 io_in[11]
port 225 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 io_in[12]
port 226 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 io_in[13]
port 227 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 io_in[14]
port 228 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 io_in[15]
port 229 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 io_in[16]
port 230 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 io_in[17]
port 231 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 io_in[18]
port 232 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 io_in[19]
port 233 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 io_in[1]
port 234 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 io_in[20]
port 235 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 io_in[21]
port 236 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 io_in[22]
port 237 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 io_in[23]
port 238 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 io_in[24]
port 239 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 io_in[25]
port 240 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 io_in[26]
port 241 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 io_in[27]
port 242 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 io_in[28]
port 243 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 io_in[29]
port 244 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 io_in[2]
port 245 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 io_in[30]
port 246 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 io_in[31]
port 247 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 io_in[32]
port 248 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 io_in[33]
port 249 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 io_in[34]
port 250 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 io_in[35]
port 251 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 io_in[36]
port 252 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 io_in[37]
port 253 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 io_in[3]
port 254 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 io_in[4]
port 255 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 io_in[5]
port 256 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 io_in[6]
port 257 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 io_in[7]
port 258 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 io_in[8]
port 259 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 io_in[9]
port 260 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 261 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 262 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 263 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 264 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 265 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 266 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 267 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 268 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 269 nsew signal tristate
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 270 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 271 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 272 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 273 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 274 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 275 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 276 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 277 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 278 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 279 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 280 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 281 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 282 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 283 nsew signal tristate
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 284 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 285 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 286 nsew signal tristate
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 287 nsew signal tristate
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 288 nsew signal tristate
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 289 nsew signal tristate
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 290 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 291 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 292 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 293 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 294 nsew signal tristate
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 295 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 296 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 297 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 298 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 io_out[0]
port 299 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 io_out[10]
port 300 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 io_out[11]
port 301 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 io_out[12]
port 302 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 io_out[13]
port 303 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 io_out[14]
port 304 nsew signal tristate
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 io_out[15]
port 305 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 io_out[16]
port 306 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 io_out[17]
port 307 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 io_out[18]
port 308 nsew signal tristate
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 io_out[19]
port 309 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 io_out[1]
port 310 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 io_out[20]
port 311 nsew signal tristate
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 io_out[21]
port 312 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 io_out[22]
port 313 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 io_out[23]
port 314 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 io_out[24]
port 315 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 io_out[25]
port 316 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 io_out[26]
port 317 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 io_out[27]
port 318 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 io_out[28]
port 319 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 io_out[29]
port 320 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 io_out[2]
port 321 nsew signal tristate
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 io_out[30]
port 322 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 io_out[31]
port 323 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 io_out[32]
port 324 nsew signal tristate
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 io_out[33]
port 325 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 io_out[34]
port 326 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 io_out[35]
port 327 nsew signal tristate
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 io_out[36]
port 328 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 io_out[37]
port 329 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 io_out[3]
port 330 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 io_out[4]
port 331 nsew signal tristate
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 io_out[5]
port 332 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 io_out[6]
port 333 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 io_out[7]
port 334 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 io_out[8]
port 335 nsew signal tristate
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 io_out[9]
port 336 nsew signal tristate
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 oeb_6502
port 337 nsew signal input
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 oeb_as1802
port 338 nsew signal input
flabel metal2 s 12622 63200 12678 64000 0 FreeSans 224 90 0 0 oeb_as2650
port 339 nsew signal input
flabel metal3 s 0 61480 800 61600 0 FreeSans 480 0 0 0 oeb_as512512512
port 340 nsew signal input
flabel metal2 s 53102 63200 53158 64000 0 FreeSans 224 90 0 0 oeb_as5401
port 341 nsew signal input
flabel metal3 s 0 36320 800 36440 0 FreeSans 480 0 0 0 oeb_mc14500
port 342 nsew signal input
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 rst_6502
port 343 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 rst_LCD
port 344 nsew signal tristate
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 rst_as1802
port 345 nsew signal tristate
flabel metal3 s 0 24080 800 24200 0 FreeSans 480 0 0 0 rst_as2650
port 346 nsew signal tristate
flabel metal3 s 0 25440 800 25560 0 FreeSans 480 0 0 0 rst_as512512512
port 347 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 rst_as5401
port 348 nsew signal tristate
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 rst_counter
port 349 nsew signal tristate
flabel metal3 s 0 26800 800 26920 0 FreeSans 480 0 0 0 rst_diceroll
port 350 nsew signal tristate
flabel metal3 s 0 27480 800 27600 0 FreeSans 480 0 0 0 rst_mc14500
port 351 nsew signal tristate
flabel metal3 s 0 28160 800 28280 0 FreeSans 480 0 0 0 rst_posit
port 352 nsew signal tristate
flabel metal3 s 0 28840 800 28960 0 FreeSans 480 0 0 0 rst_tbb1143
port 353 nsew signal tristate
flabel metal3 s 0 29520 800 29640 0 FreeSans 480 0 0 0 rst_tune
port 354 nsew signal tristate
flabel metal4 s 4208 2128 4528 61520 0 FreeSans 1920 90 0 0 vccd1
port 355 nsew power bidirectional
flabel metal4 s 34928 2128 35248 61520 0 FreeSans 1920 90 0 0 vccd1
port 355 nsew power bidirectional
flabel metal4 s 19568 2128 19888 61520 0 FreeSans 1920 90 0 0 vssd1
port 356 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 61520 0 FreeSans 1920 90 0 0 vssd1
port 356 nsew ground bidirectional
flabel metal3 s 59200 1096 60000 1216 0 FreeSans 480 0 0 0 wb_clk_i
port 357 nsew signal input
flabel metal3 s 59200 1640 60000 1760 0 FreeSans 480 0 0 0 wb_rst_i
port 358 nsew signal input
flabel metal3 s 59200 2184 60000 2304 0 FreeSans 480 0 0 0 wbs_ack_o
port 359 nsew signal tristate
flabel metal3 s 59200 4360 60000 4480 0 FreeSans 480 0 0 0 wbs_adr_i[0]
port 360 nsew signal input
flabel metal3 s 59200 20680 60000 20800 0 FreeSans 480 0 0 0 wbs_adr_i[10]
port 361 nsew signal input
flabel metal3 s 59200 22312 60000 22432 0 FreeSans 480 0 0 0 wbs_adr_i[11]
port 362 nsew signal input
flabel metal3 s 59200 23944 60000 24064 0 FreeSans 480 0 0 0 wbs_adr_i[12]
port 363 nsew signal input
flabel metal3 s 59200 25576 60000 25696 0 FreeSans 480 0 0 0 wbs_adr_i[13]
port 364 nsew signal input
flabel metal3 s 59200 27208 60000 27328 0 FreeSans 480 0 0 0 wbs_adr_i[14]
port 365 nsew signal input
flabel metal3 s 59200 28840 60000 28960 0 FreeSans 480 0 0 0 wbs_adr_i[15]
port 366 nsew signal input
flabel metal3 s 59200 30472 60000 30592 0 FreeSans 480 0 0 0 wbs_adr_i[16]
port 367 nsew signal input
flabel metal3 s 59200 32104 60000 32224 0 FreeSans 480 0 0 0 wbs_adr_i[17]
port 368 nsew signal input
flabel metal3 s 59200 33736 60000 33856 0 FreeSans 480 0 0 0 wbs_adr_i[18]
port 369 nsew signal input
flabel metal3 s 59200 35368 60000 35488 0 FreeSans 480 0 0 0 wbs_adr_i[19]
port 370 nsew signal input
flabel metal3 s 59200 5992 60000 6112 0 FreeSans 480 0 0 0 wbs_adr_i[1]
port 371 nsew signal input
flabel metal3 s 59200 37000 60000 37120 0 FreeSans 480 0 0 0 wbs_adr_i[20]
port 372 nsew signal input
flabel metal3 s 59200 38632 60000 38752 0 FreeSans 480 0 0 0 wbs_adr_i[21]
port 373 nsew signal input
flabel metal3 s 59200 40264 60000 40384 0 FreeSans 480 0 0 0 wbs_adr_i[22]
port 374 nsew signal input
flabel metal3 s 59200 41896 60000 42016 0 FreeSans 480 0 0 0 wbs_adr_i[23]
port 375 nsew signal input
flabel metal3 s 59200 43528 60000 43648 0 FreeSans 480 0 0 0 wbs_adr_i[24]
port 376 nsew signal input
flabel metal3 s 59200 45160 60000 45280 0 FreeSans 480 0 0 0 wbs_adr_i[25]
port 377 nsew signal input
flabel metal3 s 59200 46792 60000 46912 0 FreeSans 480 0 0 0 wbs_adr_i[26]
port 378 nsew signal input
flabel metal3 s 59200 48424 60000 48544 0 FreeSans 480 0 0 0 wbs_adr_i[27]
port 379 nsew signal input
flabel metal3 s 59200 50056 60000 50176 0 FreeSans 480 0 0 0 wbs_adr_i[28]
port 380 nsew signal input
flabel metal3 s 59200 51688 60000 51808 0 FreeSans 480 0 0 0 wbs_adr_i[29]
port 381 nsew signal input
flabel metal3 s 59200 7624 60000 7744 0 FreeSans 480 0 0 0 wbs_adr_i[2]
port 382 nsew signal input
flabel metal3 s 59200 53320 60000 53440 0 FreeSans 480 0 0 0 wbs_adr_i[30]
port 383 nsew signal input
flabel metal3 s 59200 54952 60000 55072 0 FreeSans 480 0 0 0 wbs_adr_i[31]
port 384 nsew signal input
flabel metal3 s 59200 9256 60000 9376 0 FreeSans 480 0 0 0 wbs_adr_i[3]
port 385 nsew signal input
flabel metal3 s 59200 10888 60000 11008 0 FreeSans 480 0 0 0 wbs_adr_i[4]
port 386 nsew signal input
flabel metal3 s 59200 12520 60000 12640 0 FreeSans 480 0 0 0 wbs_adr_i[5]
port 387 nsew signal input
flabel metal3 s 59200 14152 60000 14272 0 FreeSans 480 0 0 0 wbs_adr_i[6]
port 388 nsew signal input
flabel metal3 s 59200 15784 60000 15904 0 FreeSans 480 0 0 0 wbs_adr_i[7]
port 389 nsew signal input
flabel metal3 s 59200 17416 60000 17536 0 FreeSans 480 0 0 0 wbs_adr_i[8]
port 390 nsew signal input
flabel metal3 s 59200 19048 60000 19168 0 FreeSans 480 0 0 0 wbs_adr_i[9]
port 391 nsew signal input
flabel metal3 s 59200 2728 60000 2848 0 FreeSans 480 0 0 0 wbs_cyc_i
port 392 nsew signal input
flabel metal3 s 59200 4904 60000 5024 0 FreeSans 480 0 0 0 wbs_dat_i[0]
port 393 nsew signal input
flabel metal3 s 59200 21224 60000 21344 0 FreeSans 480 0 0 0 wbs_dat_i[10]
port 394 nsew signal input
flabel metal3 s 59200 22856 60000 22976 0 FreeSans 480 0 0 0 wbs_dat_i[11]
port 395 nsew signal input
flabel metal3 s 59200 24488 60000 24608 0 FreeSans 480 0 0 0 wbs_dat_i[12]
port 396 nsew signal input
flabel metal3 s 59200 26120 60000 26240 0 FreeSans 480 0 0 0 wbs_dat_i[13]
port 397 nsew signal input
flabel metal3 s 59200 27752 60000 27872 0 FreeSans 480 0 0 0 wbs_dat_i[14]
port 398 nsew signal input
flabel metal3 s 59200 29384 60000 29504 0 FreeSans 480 0 0 0 wbs_dat_i[15]
port 399 nsew signal input
flabel metal3 s 59200 31016 60000 31136 0 FreeSans 480 0 0 0 wbs_dat_i[16]
port 400 nsew signal input
flabel metal3 s 59200 32648 60000 32768 0 FreeSans 480 0 0 0 wbs_dat_i[17]
port 401 nsew signal input
flabel metal3 s 59200 34280 60000 34400 0 FreeSans 480 0 0 0 wbs_dat_i[18]
port 402 nsew signal input
flabel metal3 s 59200 35912 60000 36032 0 FreeSans 480 0 0 0 wbs_dat_i[19]
port 403 nsew signal input
flabel metal3 s 59200 6536 60000 6656 0 FreeSans 480 0 0 0 wbs_dat_i[1]
port 404 nsew signal input
flabel metal3 s 59200 37544 60000 37664 0 FreeSans 480 0 0 0 wbs_dat_i[20]
port 405 nsew signal input
flabel metal3 s 59200 39176 60000 39296 0 FreeSans 480 0 0 0 wbs_dat_i[21]
port 406 nsew signal input
flabel metal3 s 59200 40808 60000 40928 0 FreeSans 480 0 0 0 wbs_dat_i[22]
port 407 nsew signal input
flabel metal3 s 59200 42440 60000 42560 0 FreeSans 480 0 0 0 wbs_dat_i[23]
port 408 nsew signal input
flabel metal3 s 59200 44072 60000 44192 0 FreeSans 480 0 0 0 wbs_dat_i[24]
port 409 nsew signal input
flabel metal3 s 59200 45704 60000 45824 0 FreeSans 480 0 0 0 wbs_dat_i[25]
port 410 nsew signal input
flabel metal3 s 59200 47336 60000 47456 0 FreeSans 480 0 0 0 wbs_dat_i[26]
port 411 nsew signal input
flabel metal3 s 59200 48968 60000 49088 0 FreeSans 480 0 0 0 wbs_dat_i[27]
port 412 nsew signal input
flabel metal3 s 59200 50600 60000 50720 0 FreeSans 480 0 0 0 wbs_dat_i[28]
port 413 nsew signal input
flabel metal3 s 59200 52232 60000 52352 0 FreeSans 480 0 0 0 wbs_dat_i[29]
port 414 nsew signal input
flabel metal3 s 59200 8168 60000 8288 0 FreeSans 480 0 0 0 wbs_dat_i[2]
port 415 nsew signal input
flabel metal3 s 59200 53864 60000 53984 0 FreeSans 480 0 0 0 wbs_dat_i[30]
port 416 nsew signal input
flabel metal3 s 59200 55496 60000 55616 0 FreeSans 480 0 0 0 wbs_dat_i[31]
port 417 nsew signal input
flabel metal3 s 59200 9800 60000 9920 0 FreeSans 480 0 0 0 wbs_dat_i[3]
port 418 nsew signal input
flabel metal3 s 59200 11432 60000 11552 0 FreeSans 480 0 0 0 wbs_dat_i[4]
port 419 nsew signal input
flabel metal3 s 59200 13064 60000 13184 0 FreeSans 480 0 0 0 wbs_dat_i[5]
port 420 nsew signal input
flabel metal3 s 59200 14696 60000 14816 0 FreeSans 480 0 0 0 wbs_dat_i[6]
port 421 nsew signal input
flabel metal3 s 59200 16328 60000 16448 0 FreeSans 480 0 0 0 wbs_dat_i[7]
port 422 nsew signal input
flabel metal3 s 59200 17960 60000 18080 0 FreeSans 480 0 0 0 wbs_dat_i[8]
port 423 nsew signal input
flabel metal3 s 59200 19592 60000 19712 0 FreeSans 480 0 0 0 wbs_dat_i[9]
port 424 nsew signal input
flabel metal3 s 59200 5448 60000 5568 0 FreeSans 480 0 0 0 wbs_dat_o[0]
port 425 nsew signal tristate
flabel metal3 s 59200 21768 60000 21888 0 FreeSans 480 0 0 0 wbs_dat_o[10]
port 426 nsew signal tristate
flabel metal3 s 59200 23400 60000 23520 0 FreeSans 480 0 0 0 wbs_dat_o[11]
port 427 nsew signal tristate
flabel metal3 s 59200 25032 60000 25152 0 FreeSans 480 0 0 0 wbs_dat_o[12]
port 428 nsew signal tristate
flabel metal3 s 59200 26664 60000 26784 0 FreeSans 480 0 0 0 wbs_dat_o[13]
port 429 nsew signal tristate
flabel metal3 s 59200 28296 60000 28416 0 FreeSans 480 0 0 0 wbs_dat_o[14]
port 430 nsew signal tristate
flabel metal3 s 59200 29928 60000 30048 0 FreeSans 480 0 0 0 wbs_dat_o[15]
port 431 nsew signal tristate
flabel metal3 s 59200 31560 60000 31680 0 FreeSans 480 0 0 0 wbs_dat_o[16]
port 432 nsew signal tristate
flabel metal3 s 59200 33192 60000 33312 0 FreeSans 480 0 0 0 wbs_dat_o[17]
port 433 nsew signal tristate
flabel metal3 s 59200 34824 60000 34944 0 FreeSans 480 0 0 0 wbs_dat_o[18]
port 434 nsew signal tristate
flabel metal3 s 59200 36456 60000 36576 0 FreeSans 480 0 0 0 wbs_dat_o[19]
port 435 nsew signal tristate
flabel metal3 s 59200 7080 60000 7200 0 FreeSans 480 0 0 0 wbs_dat_o[1]
port 436 nsew signal tristate
flabel metal3 s 59200 38088 60000 38208 0 FreeSans 480 0 0 0 wbs_dat_o[20]
port 437 nsew signal tristate
flabel metal3 s 59200 39720 60000 39840 0 FreeSans 480 0 0 0 wbs_dat_o[21]
port 438 nsew signal tristate
flabel metal3 s 59200 41352 60000 41472 0 FreeSans 480 0 0 0 wbs_dat_o[22]
port 439 nsew signal tristate
flabel metal3 s 59200 42984 60000 43104 0 FreeSans 480 0 0 0 wbs_dat_o[23]
port 440 nsew signal tristate
flabel metal3 s 59200 44616 60000 44736 0 FreeSans 480 0 0 0 wbs_dat_o[24]
port 441 nsew signal tristate
flabel metal3 s 59200 46248 60000 46368 0 FreeSans 480 0 0 0 wbs_dat_o[25]
port 442 nsew signal tristate
flabel metal3 s 59200 47880 60000 48000 0 FreeSans 480 0 0 0 wbs_dat_o[26]
port 443 nsew signal tristate
flabel metal3 s 59200 49512 60000 49632 0 FreeSans 480 0 0 0 wbs_dat_o[27]
port 444 nsew signal tristate
flabel metal3 s 59200 51144 60000 51264 0 FreeSans 480 0 0 0 wbs_dat_o[28]
port 445 nsew signal tristate
flabel metal3 s 59200 52776 60000 52896 0 FreeSans 480 0 0 0 wbs_dat_o[29]
port 446 nsew signal tristate
flabel metal3 s 59200 8712 60000 8832 0 FreeSans 480 0 0 0 wbs_dat_o[2]
port 447 nsew signal tristate
flabel metal3 s 59200 54408 60000 54528 0 FreeSans 480 0 0 0 wbs_dat_o[30]
port 448 nsew signal tristate
flabel metal3 s 59200 56040 60000 56160 0 FreeSans 480 0 0 0 wbs_dat_o[31]
port 449 nsew signal tristate
flabel metal3 s 59200 10344 60000 10464 0 FreeSans 480 0 0 0 wbs_dat_o[3]
port 450 nsew signal tristate
flabel metal3 s 59200 11976 60000 12096 0 FreeSans 480 0 0 0 wbs_dat_o[4]
port 451 nsew signal tristate
flabel metal3 s 59200 13608 60000 13728 0 FreeSans 480 0 0 0 wbs_dat_o[5]
port 452 nsew signal tristate
flabel metal3 s 59200 15240 60000 15360 0 FreeSans 480 0 0 0 wbs_dat_o[6]
port 453 nsew signal tristate
flabel metal3 s 59200 16872 60000 16992 0 FreeSans 480 0 0 0 wbs_dat_o[7]
port 454 nsew signal tristate
flabel metal3 s 59200 18504 60000 18624 0 FreeSans 480 0 0 0 wbs_dat_o[8]
port 455 nsew signal tristate
flabel metal3 s 59200 20136 60000 20256 0 FreeSans 480 0 0 0 wbs_dat_o[9]
port 456 nsew signal tristate
flabel metal3 s 59200 3272 60000 3392 0 FreeSans 480 0 0 0 wbs_stb_i
port 457 nsew signal input
flabel metal3 s 59200 3816 60000 3936 0 FreeSans 480 0 0 0 wbs_we_i
port 458 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 64000
<< end >>
