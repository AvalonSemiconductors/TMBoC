VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tholin_avalonsemi_5401
  CLASS BLOCK ;
  FOREIGN tholin_avalonsemi_5401 ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 146.000 6.810 150.000 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 146.000 31.650 150.000 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 146.000 44.070 150.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 146.000 56.490 150.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 146.000 68.910 150.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 146.000 81.330 150.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 146.000 93.750 150.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 146.000 106.170 150.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 146.000 118.590 150.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 146.000 131.010 150.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 146.000 143.430 150.000 ;
    END
  END io_in[9]
  PIN io_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 74.160 150.000 74.760 ;
    END
  END io_oeb
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 146.000 19.230 150.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.085 10.640 23.685 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.815 10.640 58.415 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.545 10.640 93.145 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.275 10.640 127.875 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.450 10.640 41.050 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.180 10.640 75.780 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.910 10.640 110.510 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.640 10.640 145.240 138.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 0.070 9.900 146.670 138.960 ;
      LAYER met2 ;
        RECT 0.100 145.720 6.250 146.610 ;
        RECT 7.090 145.720 18.670 146.610 ;
        RECT 19.510 145.720 31.090 146.610 ;
        RECT 31.930 145.720 43.510 146.610 ;
        RECT 44.350 145.720 55.930 146.610 ;
        RECT 56.770 145.720 68.350 146.610 ;
        RECT 69.190 145.720 80.770 146.610 ;
        RECT 81.610 145.720 93.190 146.610 ;
        RECT 94.030 145.720 105.610 146.610 ;
        RECT 106.450 145.720 118.030 146.610 ;
        RECT 118.870 145.720 130.450 146.610 ;
        RECT 131.290 145.720 142.870 146.610 ;
        RECT 143.710 145.720 146.640 146.610 ;
        RECT 0.100 4.280 146.640 145.720 ;
        RECT 0.100 3.670 2.570 4.280 ;
        RECT 3.410 3.670 8.090 4.280 ;
        RECT 8.930 3.670 13.610 4.280 ;
        RECT 14.450 3.670 19.130 4.280 ;
        RECT 19.970 3.670 24.650 4.280 ;
        RECT 25.490 3.670 30.170 4.280 ;
        RECT 31.010 3.670 35.690 4.280 ;
        RECT 36.530 3.670 41.210 4.280 ;
        RECT 42.050 3.670 46.730 4.280 ;
        RECT 47.570 3.670 52.250 4.280 ;
        RECT 53.090 3.670 57.770 4.280 ;
        RECT 58.610 3.670 63.290 4.280 ;
        RECT 64.130 3.670 68.810 4.280 ;
        RECT 69.650 3.670 74.330 4.280 ;
        RECT 75.170 3.670 79.850 4.280 ;
        RECT 80.690 3.670 85.370 4.280 ;
        RECT 86.210 3.670 90.890 4.280 ;
        RECT 91.730 3.670 96.410 4.280 ;
        RECT 97.250 3.670 101.930 4.280 ;
        RECT 102.770 3.670 107.450 4.280 ;
        RECT 108.290 3.670 112.970 4.280 ;
        RECT 113.810 3.670 118.490 4.280 ;
        RECT 119.330 3.670 124.010 4.280 ;
        RECT 124.850 3.670 129.530 4.280 ;
        RECT 130.370 3.670 135.050 4.280 ;
        RECT 135.890 3.670 140.570 4.280 ;
        RECT 141.410 3.670 146.090 4.280 ;
      LAYER met3 ;
        RECT 9.265 75.160 146.000 138.885 ;
        RECT 9.265 73.760 145.600 75.160 ;
        RECT 9.265 10.715 146.000 73.760 ;
      LAYER met4 ;
        RECT 20.535 18.535 21.685 131.745 ;
        RECT 24.085 18.535 39.050 131.745 ;
        RECT 41.450 18.535 56.415 131.745 ;
        RECT 58.815 18.535 73.780 131.745 ;
        RECT 76.180 18.535 91.145 131.745 ;
        RECT 93.545 18.535 98.145 131.745 ;
  END
END tholin_avalonsemi_5401
END LIBRARY

