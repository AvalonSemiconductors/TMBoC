// This is the unpowered netlist.
module tt2_tholin_diceroll (clk,
    io_in,
    rst,
    io_out);
 input clk;
 input io_in;
 input rst;
 output [7:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire \dice.bcd[0] ;
 wire \dice.bcd[1] ;
 wire \dice.bcd[2] ;
 wire \dice.clkdiv[0] ;
 wire \dice.clkdiv[1] ;
 wire \dice.clkdiv[2] ;
 wire \dice.clkdiv[3] ;
 wire \dice.clkdiv[4] ;
 wire \dice.clkdiv[5] ;
 wire \dice.clkdiv[6] ;
 wire \dice.clkdiv[7] ;
 wire \dice.counter[0] ;
 wire \dice.counter[10] ;
 wire \dice.counter[11] ;
 wire \dice.counter[12] ;
 wire \dice.counter[13] ;
 wire \dice.counter[14] ;
 wire \dice.counter[15] ;
 wire \dice.counter[1] ;
 wire \dice.counter[2] ;
 wire \dice.counter[3] ;
 wire \dice.counter[4] ;
 wire \dice.counter[5] ;
 wire \dice.counter[6] ;
 wire \dice.counter[7] ;
 wire \dice.counter[8] ;
 wire \dice.counter[9] ;
 wire \dice.lfsr[0] ;
 wire \dice.lfsr[10] ;
 wire \dice.lfsr[11] ;
 wire \dice.lfsr[12] ;
 wire \dice.lfsr[13] ;
 wire \dice.lfsr[14] ;
 wire \dice.lfsr[15] ;
 wire \dice.lfsr[1] ;
 wire \dice.lfsr[2] ;
 wire \dice.lfsr[3] ;
 wire \dice.lfsr[4] ;
 wire \dice.lfsr[5] ;
 wire \dice.lfsr[6] ;
 wire \dice.lfsr[7] ;
 wire \dice.lfsr[8] ;
 wire \dice.lfsr[9] ;
 wire \dice.r_counter[0] ;
 wire \dice.r_counter[1] ;
 wire \dice.r_counter[2] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__inv_2 _181_ (.A(\dice.bcd[2] ),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _182_ (.A(\dice.bcd[0] ),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _183_ (.A(net19),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _184_ (.A(\dice.clkdiv[5] ),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _185_ (.A(\dice.counter[13] ),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _186_ (.A(net15),
    .Y(_059_));
 sky130_fd_sc_hd__and2_1 _187_ (.A(\dice.lfsr[1] ),
    .B(\dice.r_counter[1] ),
    .X(_060_));
 sky130_fd_sc_hd__xor2_4 _188_ (.A(\dice.lfsr[1] ),
    .B(\dice.r_counter[1] ),
    .X(_061_));
 sky130_fd_sc_hd__nand2_2 _189_ (.A(\dice.lfsr[0] ),
    .B(\dice.r_counter[0] ),
    .Y(_062_));
 sky130_fd_sc_hd__xor2_2 _190_ (.A(_061_),
    .B(_062_),
    .X(_063_));
 sky130_fd_sc_hd__a31o_1 _191_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.r_counter[0] ),
    .A3(_061_),
    .B1(_060_),
    .X(_064_));
 sky130_fd_sc_hd__xnor2_2 _192_ (.A(\dice.lfsr[2] ),
    .B(\dice.r_counter[2] ),
    .Y(_065_));
 sky130_fd_sc_hd__xnor2_2 _193_ (.A(_064_),
    .B(_065_),
    .Y(_066_));
 sky130_fd_sc_hd__nand2_1 _194_ (.A(_063_),
    .B(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__or3_1 _195_ (.A(net20),
    .B(\dice.counter[1] ),
    .C(\dice.clkdiv[1] ),
    .X(_068_));
 sky130_fd_sc_hd__nand3b_1 _196_ (.A_N(net20),
    .B(\dice.counter[1] ),
    .C(\dice.clkdiv[1] ),
    .Y(_069_));
 sky130_fd_sc_hd__o21ba_1 _197_ (.A1(\dice.counter[6] ),
    .A2(\dice.clkdiv[6] ),
    .B1_N(net20),
    .X(_070_));
 sky130_fd_sc_hd__nand3b_1 _198_ (.A_N(net20),
    .B(\dice.counter[6] ),
    .C(\dice.clkdiv[6] ),
    .Y(_071_));
 sky130_fd_sc_hd__a22o_1 _199_ (.A1(_068_),
    .A2(_069_),
    .B1(_070_),
    .B2(_071_),
    .X(_072_));
 sky130_fd_sc_hd__and2_1 _200_ (.A(net13),
    .B(\dice.counter[12] ),
    .X(_073_));
 sky130_fd_sc_hd__and2_1 _201_ (.A(net13),
    .B(\dice.counter[10] ),
    .X(_074_));
 sky130_fd_sc_hd__nand2b_2 _202_ (.A_N(net19),
    .B(\dice.clkdiv[2] ),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _203_ (.A(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__and2_1 _204_ (.A(net13),
    .B(\dice.counter[8] ),
    .X(_077_));
 sky130_fd_sc_hd__and2_1 _205_ (.A(net13),
    .B(\dice.counter[9] ),
    .X(_078_));
 sky130_fd_sc_hd__xor2_1 _206_ (.A(\dice.counter[0] ),
    .B(\dice.clkdiv[0] ),
    .X(_079_));
 sky130_fd_sc_hd__and2b_1 _207_ (.A_N(\dice.clkdiv[2] ),
    .B(\dice.counter[2] ),
    .X(_080_));
 sky130_fd_sc_hd__o41a_1 _208_ (.A1(\dice.counter[14] ),
    .A2(\dice.counter[15] ),
    .A3(_079_),
    .A4(_080_),
    .B1(net13),
    .X(_081_));
 sky130_fd_sc_hd__and2b_1 _209_ (.A_N(\dice.counter[4] ),
    .B(\dice.clkdiv[4] ),
    .X(_082_));
 sky130_fd_sc_hd__nand2b_2 _210_ (.A_N(net19),
    .B(\dice.clkdiv[7] ),
    .Y(_083_));
 sky130_fd_sc_hd__or3b_1 _211_ (.A(net20),
    .B(\dice.clkdiv[4] ),
    .C_N(\dice.counter[4] ),
    .X(_084_));
 sky130_fd_sc_hd__or3b_1 _212_ (.A(net19),
    .B(\dice.clkdiv[7] ),
    .C_N(\dice.counter[7] ),
    .X(_085_));
 sky130_fd_sc_hd__nand2b_2 _213_ (.A_N(net21),
    .B(\dice.counter[3] ),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _214_ (.A(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__nand2b_1 _215_ (.A_N(net20),
    .B(\dice.clkdiv[3] ),
    .Y(_088_));
 sky130_fd_sc_hd__mux2_1 _216_ (.A0(\dice.clkdiv[3] ),
    .A1(_088_),
    .S(_086_),
    .X(_089_));
 sky130_fd_sc_hd__and2b_2 _217_ (.A_N(net19),
    .B(\dice.counter[5] ),
    .X(_090_));
 sky130_fd_sc_hd__o41a_1 _218_ (.A1(\dice.counter[8] ),
    .A2(\dice.counter[9] ),
    .A3(\dice.counter[11] ),
    .A4(\dice.counter[13] ),
    .B1(net14),
    .X(_091_));
 sky130_fd_sc_hd__or4b_4 _219_ (.A(_072_),
    .B(_091_),
    .C(_081_),
    .D_N(_089_),
    .X(_092_));
 sky130_fd_sc_hd__o21ai_1 _220_ (.A1(\dice.counter[2] ),
    .A2(_075_),
    .B1(_084_),
    .Y(_093_));
 sky130_fd_sc_hd__a2bb2o_1 _221_ (.A1_N(\dice.counter[7] ),
    .A2_N(_083_),
    .B1(_090_),
    .B2(_057_),
    .X(_094_));
 sky130_fd_sc_hd__o31ai_1 _222_ (.A1(net19),
    .A2(\dice.counter[5] ),
    .A3(_057_),
    .B1(_085_),
    .Y(_095_));
 sky130_fd_sc_hd__o31a_1 _223_ (.A1(\dice.counter[10] ),
    .A2(\dice.counter[12] ),
    .A3(_082_),
    .B1(net13),
    .X(_096_));
 sky130_fd_sc_hd__or4_4 _224_ (.A(_093_),
    .B(_094_),
    .C(_095_),
    .D(_096_),
    .X(_097_));
 sky130_fd_sc_hd__or3b_1 _225_ (.A(\dice.clkdiv[4] ),
    .B(\dice.clkdiv[6] ),
    .C_N(\dice.clkdiv[5] ),
    .X(_098_));
 sky130_fd_sc_hd__or4_1 _226_ (.A(\dice.clkdiv[0] ),
    .B(\dice.clkdiv[1] ),
    .C(\dice.clkdiv[2] ),
    .D(\dice.clkdiv[3] ),
    .X(_099_));
 sky130_fd_sc_hd__nor3_2 _227_ (.A(_083_),
    .B(_098_),
    .C(_099_),
    .Y(_100_));
 sky130_fd_sc_hd__or3_4 _228_ (.A(\dice.clkdiv[2] ),
    .B(\dice.clkdiv[4] ),
    .C(\dice.clkdiv[6] ),
    .X(_101_));
 sky130_fd_sc_hd__and2b_2 _229_ (.A_N(net19),
    .B(\dice.clkdiv[0] ),
    .X(_102_));
 sky130_fd_sc_hd__or3b_4 _230_ (.A(net20),
    .B(\dice.clkdiv[3] ),
    .C_N(\dice.clkdiv[7] ),
    .X(_103_));
 sky130_fd_sc_hd__or3b_4 _231_ (.A(net19),
    .B(\dice.clkdiv[1] ),
    .C_N(\dice.clkdiv[5] ),
    .X(_104_));
 sky130_fd_sc_hd__nor4_4 _232_ (.A(_101_),
    .B(_102_),
    .C(_103_),
    .D(_104_),
    .Y(_105_));
 sky130_fd_sc_hd__or4_4 _233_ (.A(_101_),
    .B(_102_),
    .C(_103_),
    .D(_104_),
    .X(_106_));
 sky130_fd_sc_hd__nor3_4 _234_ (.A(_092_),
    .B(_097_),
    .C(_105_),
    .Y(_107_));
 sky130_fd_sc_hd__or2_1 _235_ (.A(\dice.lfsr[0] ),
    .B(\dice.r_counter[0] ),
    .X(_108_));
 sky130_fd_sc_hd__and2_1 _236_ (.A(_062_),
    .B(_108_),
    .X(_109_));
 sky130_fd_sc_hd__nand2_1 _237_ (.A(_062_),
    .B(_108_),
    .Y(_110_));
 sky130_fd_sc_hd__nand2_1 _238_ (.A(_061_),
    .B(_109_),
    .Y(_111_));
 sky130_fd_sc_hd__or2_1 _239_ (.A(_066_),
    .B(_111_),
    .X(_112_));
 sky130_fd_sc_hd__o31a_1 _240_ (.A1(_092_),
    .A2(_097_),
    .A3(_105_),
    .B1(_054_),
    .X(_113_));
 sky130_fd_sc_hd__a311o_4 _241_ (.A1(_067_),
    .A2(_107_),
    .A3(_112_),
    .B1(_113_),
    .C1(net15),
    .X(_114_));
 sky130_fd_sc_hd__inv_2 _242_ (.A(_114_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_4 _243_ (.A(net16),
    .B(_107_),
    .Y(_115_));
 sky130_fd_sc_hd__o311a_1 _244_ (.A1(_092_),
    .A2(_097_),
    .A3(_105_),
    .B1(net11),
    .C1(_055_),
    .X(_116_));
 sky130_fd_sc_hd__mux2_2 _245_ (.A0(_109_),
    .A1(_111_),
    .S(_066_),
    .X(_117_));
 sky130_fd_sc_hd__nand2_1 _246_ (.A(_063_),
    .B(_110_),
    .Y(_118_));
 sky130_fd_sc_hd__a211o_1 _247_ (.A1(_063_),
    .A2(_110_),
    .B1(_100_),
    .C1(net15),
    .X(_119_));
 sky130_fd_sc_hd__nor3_2 _248_ (.A(_092_),
    .B(_097_),
    .C(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__a21oi_4 _249_ (.A1(_117_),
    .A2(_120_),
    .B1(_116_),
    .Y(_051_));
 sky130_fd_sc_hd__o31a_1 _250_ (.A1(_092_),
    .A2(_097_),
    .A3(_105_),
    .B1(\dice.bcd[1] ),
    .X(_121_));
 sky130_fd_sc_hd__a31o_2 _251_ (.A1(_107_),
    .A2(_112_),
    .A3(_118_),
    .B1(_121_),
    .X(_122_));
 sky130_fd_sc_hd__nand2_1 _252_ (.A(net11),
    .B(_122_),
    .Y(_123_));
 sky130_fd_sc_hd__inv_2 _253_ (.A(_123_),
    .Y(_052_));
 sky130_fd_sc_hd__nand2_1 _254_ (.A(_114_),
    .B(_052_),
    .Y(_124_));
 sky130_fd_sc_hd__a21o_1 _255_ (.A1(_051_),
    .A2(_123_),
    .B1(_053_),
    .X(_125_));
 sky130_fd_sc_hd__a21bo_1 _256_ (.A1(_053_),
    .A2(_051_),
    .B1_N(_125_),
    .X(_000_));
 sky130_fd_sc_hd__a31o_1 _257_ (.A1(net11),
    .A2(_051_),
    .A3(_122_),
    .B1(_114_),
    .X(_126_));
 sky130_fd_sc_hd__o21bai_2 _258_ (.A1(_051_),
    .A2(_122_),
    .B1_N(_126_),
    .Y(_009_));
 sky130_fd_sc_hd__nand2_1 _259_ (.A(_125_),
    .B(_009_),
    .Y(_001_));
 sky130_fd_sc_hd__o21ba_1 _260_ (.A1(_114_),
    .A2(_122_),
    .B1_N(_051_),
    .X(_002_));
 sky130_fd_sc_hd__o21ai_1 _261_ (.A1(_051_),
    .A2(_122_),
    .B1(_126_),
    .Y(_003_));
 sky130_fd_sc_hd__nand2_1 _262_ (.A(_124_),
    .B(_126_),
    .Y(_004_));
 sky130_fd_sc_hd__or2_1 _263_ (.A(_051_),
    .B(_124_),
    .X(_005_));
 sky130_fd_sc_hd__nor2_1 _264_ (.A(\dice.r_counter[0] ),
    .B(net15),
    .Y(_006_));
 sky130_fd_sc_hd__a21oi_1 _265_ (.A1(\dice.r_counter[1] ),
    .A2(\dice.r_counter[0] ),
    .B1(net15),
    .Y(_127_));
 sky130_fd_sc_hd__o21a_1 _266_ (.A1(\dice.r_counter[1] ),
    .A2(\dice.r_counter[0] ),
    .B1(_127_),
    .X(_007_));
 sky130_fd_sc_hd__a21oi_1 _267_ (.A1(\dice.r_counter[1] ),
    .A2(\dice.r_counter[0] ),
    .B1(\dice.r_counter[2] ),
    .Y(_128_));
 sky130_fd_sc_hd__a31o_1 _268_ (.A1(\dice.r_counter[2] ),
    .A2(\dice.r_counter[1] ),
    .A3(\dice.r_counter[0] ),
    .B1(net15),
    .X(_129_));
 sky130_fd_sc_hd__nor2_1 _269_ (.A(_128_),
    .B(_129_),
    .Y(_008_));
 sky130_fd_sc_hd__a211o_1 _270_ (.A1(net10),
    .A2(net14),
    .B1(net16),
    .C1(_105_),
    .X(_010_));
 sky130_fd_sc_hd__and4bb_2 _271_ (.A_N(_092_),
    .B_N(_097_),
    .C(_102_),
    .D(_106_),
    .X(_130_));
 sky130_fd_sc_hd__nor2_1 _272_ (.A(net16),
    .B(_130_),
    .Y(_131_));
 sky130_fd_sc_hd__o21a_1 _273_ (.A1(_102_),
    .A2(_107_),
    .B1(_131_),
    .X(_011_));
 sky130_fd_sc_hd__or3_1 _274_ (.A(net19),
    .B(\dice.clkdiv[1] ),
    .C(_130_),
    .X(_132_));
 sky130_fd_sc_hd__nand2_1 _275_ (.A(\dice.clkdiv[1] ),
    .B(_130_),
    .Y(_133_));
 sky130_fd_sc_hd__and3_1 _276_ (.A(net11),
    .B(_132_),
    .C(_133_),
    .X(_012_));
 sky130_fd_sc_hd__a31o_1 _277_ (.A1(\dice.clkdiv[1] ),
    .A2(_076_),
    .A3(_130_),
    .B1(net16),
    .X(_134_));
 sky130_fd_sc_hd__a21oi_1 _278_ (.A1(_075_),
    .A2(_133_),
    .B1(_134_),
    .Y(_013_));
 sky130_fd_sc_hd__o21a_1 _279_ (.A1(_075_),
    .A2(_133_),
    .B1(_088_),
    .X(_135_));
 sky130_fd_sc_hd__and4_2 _280_ (.A(\dice.clkdiv[1] ),
    .B(\dice.clkdiv[3] ),
    .C(_076_),
    .D(_130_),
    .X(_136_));
 sky130_fd_sc_hd__nor3_1 _281_ (.A(net16),
    .B(_135_),
    .C(_136_),
    .Y(_014_));
 sky130_fd_sc_hd__a21oi_1 _282_ (.A1(net14),
    .A2(\dice.clkdiv[4] ),
    .B1(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__a211oi_1 _283_ (.A1(\dice.clkdiv[4] ),
    .A2(_136_),
    .B1(_137_),
    .C1(net16),
    .Y(_015_));
 sky130_fd_sc_hd__and4_2 _284_ (.A(net14),
    .B(\dice.clkdiv[4] ),
    .C(\dice.clkdiv[5] ),
    .D(_136_),
    .X(_138_));
 sky130_fd_sc_hd__o2bb2a_1 _285_ (.A1_N(\dice.clkdiv[4] ),
    .A2_N(_136_),
    .B1(_057_),
    .B2(net19),
    .X(_139_));
 sky130_fd_sc_hd__o21ai_1 _286_ (.A1(_138_),
    .A2(_139_),
    .B1(net12),
    .Y(_016_));
 sky130_fd_sc_hd__a21oi_1 _287_ (.A1(net14),
    .A2(\dice.clkdiv[6] ),
    .B1(_138_),
    .Y(_140_));
 sky130_fd_sc_hd__a211oi_1 _288_ (.A1(\dice.clkdiv[6] ),
    .A2(_138_),
    .B1(_140_),
    .C1(net15),
    .Y(_017_));
 sky130_fd_sc_hd__and3_1 _289_ (.A(\dice.clkdiv[6] ),
    .B(_083_),
    .C(_138_),
    .X(_141_));
 sky130_fd_sc_hd__a21oi_1 _290_ (.A1(\dice.clkdiv[6] ),
    .A2(_138_),
    .B1(_083_),
    .Y(_142_));
 sky130_fd_sc_hd__or3_1 _291_ (.A(net16),
    .B(_141_),
    .C(_142_),
    .X(_018_));
 sky130_fd_sc_hd__and2b_1 _292_ (.A_N(net20),
    .B(\dice.counter[0] ),
    .X(_143_));
 sky130_fd_sc_hd__nand2_1 _293_ (.A(_106_),
    .B(_143_),
    .Y(_144_));
 sky130_fd_sc_hd__or2_1 _294_ (.A(_106_),
    .B(_143_),
    .X(_145_));
 sky130_fd_sc_hd__and3_1 _295_ (.A(_115_),
    .B(_144_),
    .C(_145_),
    .X(_019_));
 sky130_fd_sc_hd__nand2_1 _296_ (.A(\dice.counter[1] ),
    .B(_143_),
    .Y(_146_));
 sky130_fd_sc_hd__o21a_1 _297_ (.A1(\dice.counter[0] ),
    .A2(\dice.counter[1] ),
    .B1(net14),
    .X(_147_));
 sky130_fd_sc_hd__o211a_1 _298_ (.A1(_092_),
    .A2(_097_),
    .B1(_146_),
    .C1(_147_),
    .X(_148_));
 sky130_fd_sc_hd__and3_1 _299_ (.A(\dice.counter[0] ),
    .B(_100_),
    .C(_148_),
    .X(_149_));
 sky130_fd_sc_hd__a21oi_1 _300_ (.A1(\dice.counter[0] ),
    .A2(_105_),
    .B1(_148_),
    .Y(_150_));
 sky130_fd_sc_hd__nor3_1 _301_ (.A(net16),
    .B(_149_),
    .C(_150_),
    .Y(_020_));
 sky130_fd_sc_hd__and3_1 _302_ (.A(\dice.counter[1] ),
    .B(\dice.counter[2] ),
    .C(_143_),
    .X(_151_));
 sky130_fd_sc_hd__nand2_1 _303_ (.A(_106_),
    .B(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__a2bb2o_1 _304_ (.A1_N(_146_),
    .A2_N(_100_),
    .B1(\dice.counter[2] ),
    .B2(net14),
    .X(_153_));
 sky130_fd_sc_hd__and3_1 _305_ (.A(_115_),
    .B(_152_),
    .C(_153_),
    .X(_021_));
 sky130_fd_sc_hd__nor2_1 _306_ (.A(_086_),
    .B(_152_),
    .Y(_154_));
 sky130_fd_sc_hd__nand2_1 _307_ (.A(_086_),
    .B(_152_),
    .Y(_155_));
 sky130_fd_sc_hd__and3b_1 _308_ (.A_N(_154_),
    .B(_155_),
    .C(_115_),
    .X(_022_));
 sky130_fd_sc_hd__a21o_1 _309_ (.A1(net13),
    .A2(\dice.counter[4] ),
    .B1(_154_),
    .X(_156_));
 sky130_fd_sc_hd__and4_2 _310_ (.A(\dice.counter[4] ),
    .B(_087_),
    .C(_106_),
    .D(_151_),
    .X(_157_));
 sky130_fd_sc_hd__and3b_1 _311_ (.A_N(_157_),
    .B(_115_),
    .C(_156_),
    .X(_023_));
 sky130_fd_sc_hd__o21ai_1 _312_ (.A1(_090_),
    .A2(_157_),
    .B1(_115_),
    .Y(_158_));
 sky130_fd_sc_hd__a21oi_1 _313_ (.A1(_090_),
    .A2(_157_),
    .B1(_158_),
    .Y(_024_));
 sky130_fd_sc_hd__a22o_1 _314_ (.A1(net13),
    .A2(\dice.counter[6] ),
    .B1(_090_),
    .B2(_157_),
    .X(_159_));
 sky130_fd_sc_hd__and2_1 _315_ (.A(\dice.counter[6] ),
    .B(_090_),
    .X(_160_));
 sky130_fd_sc_hd__and2_1 _316_ (.A(_157_),
    .B(_160_),
    .X(_161_));
 sky130_fd_sc_hd__and3b_1 _317_ (.A_N(_161_),
    .B(_115_),
    .C(_159_),
    .X(_025_));
 sky130_fd_sc_hd__and3_1 _318_ (.A(\dice.counter[7] ),
    .B(_157_),
    .C(_160_),
    .X(_162_));
 sky130_fd_sc_hd__a21o_1 _319_ (.A1(net13),
    .A2(\dice.counter[7] ),
    .B1(_161_),
    .X(_163_));
 sky130_fd_sc_hd__and3b_1 _320_ (.A_N(_162_),
    .B(_163_),
    .C(_115_),
    .X(_026_));
 sky130_fd_sc_hd__and4_2 _321_ (.A(\dice.counter[7] ),
    .B(_077_),
    .C(_157_),
    .D(_160_),
    .X(_164_));
 sky130_fd_sc_hd__inv_2 _322_ (.A(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__o211a_1 _323_ (.A1(_077_),
    .A2(_162_),
    .B1(_165_),
    .C1(_115_),
    .X(_027_));
 sky130_fd_sc_hd__nand2_1 _324_ (.A(\dice.counter[9] ),
    .B(_164_),
    .Y(_166_));
 sky130_fd_sc_hd__o211a_1 _325_ (.A1(_078_),
    .A2(_164_),
    .B1(_166_),
    .C1(net12),
    .X(_028_));
 sky130_fd_sc_hd__a21oi_1 _326_ (.A1(\dice.counter[9] ),
    .A2(_164_),
    .B1(_074_),
    .Y(_167_));
 sky130_fd_sc_hd__and3_1 _327_ (.A(\dice.counter[9] ),
    .B(_074_),
    .C(_164_),
    .X(_168_));
 sky130_fd_sc_hd__nor3_1 _328_ (.A(net16),
    .B(_167_),
    .C(_168_),
    .Y(_029_));
 sky130_fd_sc_hd__a21oi_1 _329_ (.A1(net13),
    .A2(\dice.counter[11] ),
    .B1(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__and4_2 _330_ (.A(\dice.counter[9] ),
    .B(\dice.counter[11] ),
    .C(_074_),
    .D(_164_),
    .X(_170_));
 sky130_fd_sc_hd__nor3_1 _331_ (.A(net16),
    .B(_169_),
    .C(_170_),
    .Y(_030_));
 sky130_fd_sc_hd__or2_1 _332_ (.A(_073_),
    .B(_170_),
    .X(_171_));
 sky130_fd_sc_hd__nand2_1 _333_ (.A(_073_),
    .B(_170_),
    .Y(_172_));
 sky130_fd_sc_hd__and3_1 _334_ (.A(net12),
    .B(_171_),
    .C(_172_),
    .X(_031_));
 sky130_fd_sc_hd__o21ai_1 _335_ (.A1(net21),
    .A2(_058_),
    .B1(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__o211a_1 _336_ (.A1(_058_),
    .A2(_172_),
    .B1(_173_),
    .C1(net12),
    .X(_032_));
 sky130_fd_sc_hd__a31oi_1 _337_ (.A1(\dice.counter[13] ),
    .A2(_073_),
    .A3(_170_),
    .B1(\dice.counter[14] ),
    .Y(_174_));
 sky130_fd_sc_hd__and4_1 _338_ (.A(\dice.counter[13] ),
    .B(\dice.counter[14] ),
    .C(_073_),
    .D(_170_),
    .X(_175_));
 sky130_fd_sc_hd__nor4_1 _339_ (.A(net21),
    .B(net17),
    .C(_174_),
    .D(_175_),
    .Y(_033_));
 sky130_fd_sc_hd__nand2_1 _340_ (.A(net14),
    .B(\dice.counter[15] ),
    .Y(_176_));
 sky130_fd_sc_hd__mux2_1 _341_ (.A0(_176_),
    .A1(\dice.counter[15] ),
    .S(_175_),
    .X(_177_));
 sky130_fd_sc_hd__nor2_1 _342_ (.A(net17),
    .B(_177_),
    .Y(_034_));
 sky130_fd_sc_hd__and2_1 _343_ (.A(\dice.lfsr[1] ),
    .B(net11),
    .X(_035_));
 sky130_fd_sc_hd__or2_1 _344_ (.A(\dice.lfsr[2] ),
    .B(net15),
    .X(_036_));
 sky130_fd_sc_hd__and2_1 _345_ (.A(net11),
    .B(\dice.lfsr[3] ),
    .X(_037_));
 sky130_fd_sc_hd__or2_1 _346_ (.A(net15),
    .B(\dice.lfsr[4] ),
    .X(_038_));
 sky130_fd_sc_hd__or2_1 _347_ (.A(net17),
    .B(\dice.lfsr[5] ),
    .X(_039_));
 sky130_fd_sc_hd__and2_1 _348_ (.A(net12),
    .B(\dice.lfsr[6] ),
    .X(_040_));
 sky130_fd_sc_hd__or2_1 _349_ (.A(net17),
    .B(\dice.lfsr[7] ),
    .X(_041_));
 sky130_fd_sc_hd__or2_1 _350_ (.A(net17),
    .B(\dice.lfsr[8] ),
    .X(_042_));
 sky130_fd_sc_hd__and2_1 _351_ (.A(net12),
    .B(\dice.lfsr[9] ),
    .X(_043_));
 sky130_fd_sc_hd__and2_1 _352_ (.A(net11),
    .B(\dice.lfsr[10] ),
    .X(_044_));
 sky130_fd_sc_hd__a21oi_1 _353_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[11] ),
    .B1(net15),
    .Y(_178_));
 sky130_fd_sc_hd__o21a_1 _354_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[11] ),
    .B1(_178_),
    .X(_045_));
 sky130_fd_sc_hd__and2_1 _355_ (.A(net11),
    .B(\dice.lfsr[12] ),
    .X(_046_));
 sky130_fd_sc_hd__a21oi_1 _356_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[13] ),
    .B1(net18),
    .Y(_179_));
 sky130_fd_sc_hd__o21a_1 _357_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[13] ),
    .B1(_179_),
    .X(_047_));
 sky130_fd_sc_hd__a21oi_1 _358_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[14] ),
    .B1(net18),
    .Y(_180_));
 sky130_fd_sc_hd__o21a_1 _359_ (.A1(\dice.lfsr[0] ),
    .A2(\dice.lfsr[14] ),
    .B1(_180_),
    .X(_048_));
 sky130_fd_sc_hd__and2_1 _360_ (.A(net11),
    .B(\dice.lfsr[15] ),
    .X(_049_));
 sky130_fd_sc_hd__and2_1 _361_ (.A(\dice.lfsr[0] ),
    .B(net11),
    .X(_050_));
 sky130_fd_sc_hd__dfxtp_1 _362_ (.CLK(clknet_2_0__leaf_clk),
    .D(_005_),
    .Q(net5));
 sky130_fd_sc_hd__dfxtp_4 _363_ (.CLK(clknet_2_0__leaf_clk),
    .D(_006_),
    .Q(\dice.r_counter[0] ));
 sky130_fd_sc_hd__dfxtp_4 _364_ (.CLK(clknet_2_0__leaf_clk),
    .D(_007_),
    .Q(\dice.r_counter[1] ));
 sky130_fd_sc_hd__dfxtp_2 _365_ (.CLK(clknet_2_0__leaf_clk),
    .D(_008_),
    .Q(\dice.r_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _366_ (.CLK(clknet_2_0__leaf_clk),
    .D(_009_),
    .Q(net4));
 sky130_fd_sc_hd__dfxtp_1 _367_ (.CLK(clknet_2_0__leaf_clk),
    .D(_000_),
    .Q(net3));
 sky130_fd_sc_hd__dfxtp_1 _368_ (.CLK(clknet_2_0__leaf_clk),
    .D(_001_),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_1 _369_ (.CLK(clknet_2_0__leaf_clk),
    .D(_002_),
    .Q(net7));
 sky130_fd_sc_hd__dfxtp_1 _370_ (.CLK(clknet_2_0__leaf_clk),
    .D(_003_),
    .Q(net8));
 sky130_fd_sc_hd__dfxtp_1 _371_ (.CLK(clknet_2_0__leaf_clk),
    .D(_004_),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_2 _372_ (.CLK(clknet_2_2__leaf_clk),
    .D(_010_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _373_ (.CLK(clknet_2_1__leaf_clk),
    .D(_011_),
    .Q(\dice.clkdiv[0] ));
 sky130_fd_sc_hd__dfxtp_4 _374_ (.CLK(clknet_2_0__leaf_clk),
    .D(_012_),
    .Q(\dice.clkdiv[1] ));
 sky130_fd_sc_hd__dfxtp_2 _375_ (.CLK(clknet_2_1__leaf_clk),
    .D(_013_),
    .Q(\dice.clkdiv[2] ));
 sky130_fd_sc_hd__dfxtp_2 _376_ (.CLK(clknet_2_1__leaf_clk),
    .D(_014_),
    .Q(\dice.clkdiv[3] ));
 sky130_fd_sc_hd__dfxtp_4 _377_ (.CLK(clknet_2_3__leaf_clk),
    .D(_015_),
    .Q(\dice.clkdiv[4] ));
 sky130_fd_sc_hd__dfxtp_1 _378_ (.CLK(clknet_2_1__leaf_clk),
    .D(_016_),
    .Q(\dice.clkdiv[5] ));
 sky130_fd_sc_hd__dfxtp_4 _379_ (.CLK(clknet_2_0__leaf_clk),
    .D(_017_),
    .Q(\dice.clkdiv[6] ));
 sky130_fd_sc_hd__dfxtp_1 _380_ (.CLK(clknet_2_1__leaf_clk),
    .D(_018_),
    .Q(\dice.clkdiv[7] ));
 sky130_fd_sc_hd__dfxtp_2 _381_ (.CLK(clknet_2_3__leaf_clk),
    .D(_019_),
    .Q(\dice.counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _382_ (.CLK(clknet_2_1__leaf_clk),
    .D(_020_),
    .Q(\dice.counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _383_ (.CLK(clknet_2_1__leaf_clk),
    .D(_021_),
    .Q(\dice.counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _384_ (.CLK(clknet_2_1__leaf_clk),
    .D(_022_),
    .Q(\dice.counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _385_ (.CLK(clknet_2_3__leaf_clk),
    .D(_023_),
    .Q(\dice.counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _386_ (.CLK(clknet_2_1__leaf_clk),
    .D(_024_),
    .Q(\dice.counter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _387_ (.CLK(clknet_2_1__leaf_clk),
    .D(_025_),
    .Q(\dice.counter[6] ));
 sky130_fd_sc_hd__dfxtp_2 _388_ (.CLK(clknet_2_1__leaf_clk),
    .D(_026_),
    .Q(\dice.counter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _389_ (.CLK(clknet_2_1__leaf_clk),
    .D(_027_),
    .Q(\dice.counter[8] ));
 sky130_fd_sc_hd__dfxtp_2 _390_ (.CLK(clknet_2_3__leaf_clk),
    .D(_028_),
    .Q(\dice.counter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _391_ (.CLK(clknet_2_3__leaf_clk),
    .D(_029_),
    .Q(\dice.counter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _392_ (.CLK(clknet_2_3__leaf_clk),
    .D(_030_),
    .Q(\dice.counter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _393_ (.CLK(clknet_2_2__leaf_clk),
    .D(_031_),
    .Q(\dice.counter[12] ));
 sky130_fd_sc_hd__dfxtp_2 _394_ (.CLK(clknet_2_3__leaf_clk),
    .D(_032_),
    .Q(\dice.counter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _395_ (.CLK(clknet_2_3__leaf_clk),
    .D(_033_),
    .Q(\dice.counter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _396_ (.CLK(clknet_2_3__leaf_clk),
    .D(_034_),
    .Q(\dice.counter[15] ));
 sky130_fd_sc_hd__dfxtp_4 _397_ (.CLK(clknet_2_2__leaf_clk),
    .D(_035_),
    .Q(\dice.lfsr[0] ));
 sky130_fd_sc_hd__dfxtp_4 _398_ (.CLK(clknet_2_0__leaf_clk),
    .D(_036_),
    .Q(\dice.lfsr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _399_ (.CLK(clknet_2_2__leaf_clk),
    .D(_037_),
    .Q(\dice.lfsr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _400_ (.CLK(clknet_2_2__leaf_clk),
    .D(_038_),
    .Q(\dice.lfsr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _401_ (.CLK(clknet_2_2__leaf_clk),
    .D(_039_),
    .Q(\dice.lfsr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _402_ (.CLK(clknet_2_3__leaf_clk),
    .D(_040_),
    .Q(\dice.lfsr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _403_ (.CLK(clknet_2_3__leaf_clk),
    .D(_041_),
    .Q(\dice.lfsr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _404_ (.CLK(clknet_2_2__leaf_clk),
    .D(_042_),
    .Q(\dice.lfsr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _405_ (.CLK(clknet_2_3__leaf_clk),
    .D(_043_),
    .Q(\dice.lfsr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _406_ (.CLK(clknet_2_2__leaf_clk),
    .D(_044_),
    .Q(\dice.lfsr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _407_ (.CLK(clknet_2_2__leaf_clk),
    .D(_045_),
    .Q(\dice.lfsr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _408_ (.CLK(clknet_2_2__leaf_clk),
    .D(_046_),
    .Q(\dice.lfsr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _409_ (.CLK(clknet_2_2__leaf_clk),
    .D(_047_),
    .Q(\dice.lfsr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _410_ (.CLK(clknet_2_2__leaf_clk),
    .D(_048_),
    .Q(\dice.lfsr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _411_ (.CLK(clknet_2_0__leaf_clk),
    .D(_049_),
    .Q(\dice.lfsr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _412_ (.CLK(clknet_2_2__leaf_clk),
    .D(_050_),
    .Q(\dice.lfsr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _413_ (.CLK(clknet_2_0__leaf_clk),
    .D(_051_),
    .Q(\dice.bcd[0] ));
 sky130_fd_sc_hd__dfxtp_1 _414_ (.CLK(clknet_2_0__leaf_clk),
    .D(_052_),
    .Q(\dice.bcd[1] ));
 sky130_fd_sc_hd__dfxtp_1 _415_ (.CLK(clknet_2_0__leaf_clk),
    .D(_053_),
    .Q(\dice.bcd[2] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_in),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(rst),
    .X(net2));
 sky130_fd_sc_hd__buf_4 output3 (.A(net3),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_4 output4 (.A(net4),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_4 output5 (.A(net5),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_4 output6 (.A(net6),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_4 output7 (.A(net7),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_4 output8 (.A(net8),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_4 output9 (.A(net9),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_4 output10 (.A(net10),
    .X(io_out[7]));
 sky130_fd_sc_hd__clkbuf_4 fanout11 (.A(_059_),
    .X(net11));
 sky130_fd_sc_hd__buf_2 fanout12 (.A(_059_),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__buf_4 fanout14 (.A(_056_),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_8 fanout15 (.A(net18),
    .X(net15));
 sky130_fd_sc_hd__buf_6 fanout16 (.A(net18),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 fanout17 (.A(net18),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 fanout18 (.A(net2),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 fanout19 (.A(net21),
    .X(net19));
 sky130_fd_sc_hd__buf_2 fanout20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__buf_2 fanout21 (.A(net1),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_209 ();
endmodule

