VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiplexer
  CLASS BLOCK ;
  FOREIGN multiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 320.000 ;
  PIN design_clk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END design_clk_o
  PIN dsi_all[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END dsi_all[0]
  PIN dsi_all[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END dsi_all[10]
  PIN dsi_all[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END dsi_all[11]
  PIN dsi_all[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END dsi_all[12]
  PIN dsi_all[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END dsi_all[13]
  PIN dsi_all[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END dsi_all[14]
  PIN dsi_all[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END dsi_all[15]
  PIN dsi_all[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END dsi_all[16]
  PIN dsi_all[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END dsi_all[17]
  PIN dsi_all[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END dsi_all[18]
  PIN dsi_all[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 4.000 74.760 ;
    END
  END dsi_all[19]
  PIN dsi_all[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END dsi_all[1]
  PIN dsi_all[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END dsi_all[20]
  PIN dsi_all[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END dsi_all[21]
  PIN dsi_all[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END dsi_all[22]
  PIN dsi_all[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END dsi_all[23]
  PIN dsi_all[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END dsi_all[24]
  PIN dsi_all[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END dsi_all[25]
  PIN dsi_all[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END dsi_all[26]
  PIN dsi_all[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END dsi_all[27]
  PIN dsi_all[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END dsi_all[2]
  PIN dsi_all[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END dsi_all[3]
  PIN dsi_all[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END dsi_all[4]
  PIN dsi_all[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END dsi_all[5]
  PIN dsi_all[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END dsi_all[6]
  PIN dsi_all[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END dsi_all[7]
  PIN dsi_all[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END dsi_all[8]
  PIN dsi_all[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END dsi_all[9]
  PIN dso_6502[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END dso_6502[0]
  PIN dso_6502[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END dso_6502[10]
  PIN dso_6502[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END dso_6502[11]
  PIN dso_6502[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END dso_6502[12]
  PIN dso_6502[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END dso_6502[13]
  PIN dso_6502[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END dso_6502[14]
  PIN dso_6502[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END dso_6502[15]
  PIN dso_6502[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END dso_6502[16]
  PIN dso_6502[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END dso_6502[17]
  PIN dso_6502[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END dso_6502[18]
  PIN dso_6502[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END dso_6502[19]
  PIN dso_6502[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END dso_6502[1]
  PIN dso_6502[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END dso_6502[20]
  PIN dso_6502[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END dso_6502[21]
  PIN dso_6502[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END dso_6502[22]
  PIN dso_6502[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END dso_6502[23]
  PIN dso_6502[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END dso_6502[24]
  PIN dso_6502[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 0.000 221.630 4.000 ;
    END
  END dso_6502[25]
  PIN dso_6502[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END dso_6502[26]
  PIN dso_6502[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END dso_6502[2]
  PIN dso_6502[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END dso_6502[3]
  PIN dso_6502[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END dso_6502[4]
  PIN dso_6502[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END dso_6502[5]
  PIN dso_6502[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END dso_6502[6]
  PIN dso_6502[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END dso_6502[7]
  PIN dso_6502[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END dso_6502[8]
  PIN dso_6502[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END dso_6502[9]
  PIN dso_LCD[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 316.000 269.470 320.000 ;
    END
  END dso_LCD[0]
  PIN dso_LCD[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 316.000 273.150 320.000 ;
    END
  END dso_LCD[1]
  PIN dso_LCD[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 316.000 276.830 320.000 ;
    END
  END dso_LCD[2]
  PIN dso_LCD[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 316.000 280.510 320.000 ;
    END
  END dso_LCD[3]
  PIN dso_LCD[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 316.000 284.190 320.000 ;
    END
  END dso_LCD[4]
  PIN dso_LCD[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 316.000 287.870 320.000 ;
    END
  END dso_LCD[5]
  PIN dso_LCD[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 316.000 291.550 320.000 ;
    END
  END dso_LCD[6]
  PIN dso_LCD[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 316.000 295.230 320.000 ;
    END
  END dso_LCD[7]
  PIN dso_as1802[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END dso_as1802[0]
  PIN dso_as1802[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END dso_as1802[10]
  PIN dso_as1802[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END dso_as1802[11]
  PIN dso_as1802[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END dso_as1802[12]
  PIN dso_as1802[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END dso_as1802[13]
  PIN dso_as1802[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END dso_as1802[14]
  PIN dso_as1802[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END dso_as1802[15]
  PIN dso_as1802[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END dso_as1802[16]
  PIN dso_as1802[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END dso_as1802[17]
  PIN dso_as1802[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END dso_as1802[18]
  PIN dso_as1802[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END dso_as1802[19]
  PIN dso_as1802[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END dso_as1802[1]
  PIN dso_as1802[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END dso_as1802[20]
  PIN dso_as1802[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END dso_as1802[21]
  PIN dso_as1802[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END dso_as1802[22]
  PIN dso_as1802[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END dso_as1802[23]
  PIN dso_as1802[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END dso_as1802[24]
  PIN dso_as1802[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END dso_as1802[25]
  PIN dso_as1802[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END dso_as1802[26]
  PIN dso_as1802[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END dso_as1802[2]
  PIN dso_as1802[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END dso_as1802[3]
  PIN dso_as1802[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END dso_as1802[4]
  PIN dso_as1802[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END dso_as1802[5]
  PIN dso_as1802[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END dso_as1802[6]
  PIN dso_as1802[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END dso_as1802[7]
  PIN dso_as1802[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END dso_as1802[8]
  PIN dso_as1802[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END dso_as1802[9]
  PIN dso_as2650[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 316.000 67.070 320.000 ;
    END
  END dso_as2650[0]
  PIN dso_as2650[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 316.000 103.870 320.000 ;
    END
  END dso_as2650[10]
  PIN dso_as2650[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 316.000 107.550 320.000 ;
    END
  END dso_as2650[11]
  PIN dso_as2650[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 316.000 111.230 320.000 ;
    END
  END dso_as2650[12]
  PIN dso_as2650[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 316.000 114.910 320.000 ;
    END
  END dso_as2650[13]
  PIN dso_as2650[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 316.000 118.590 320.000 ;
    END
  END dso_as2650[14]
  PIN dso_as2650[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 316.000 122.270 320.000 ;
    END
  END dso_as2650[15]
  PIN dso_as2650[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 316.000 125.950 320.000 ;
    END
  END dso_as2650[16]
  PIN dso_as2650[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 316.000 129.630 320.000 ;
    END
  END dso_as2650[17]
  PIN dso_as2650[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 316.000 133.310 320.000 ;
    END
  END dso_as2650[18]
  PIN dso_as2650[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 316.000 136.990 320.000 ;
    END
  END dso_as2650[19]
  PIN dso_as2650[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 316.000 70.750 320.000 ;
    END
  END dso_as2650[1]
  PIN dso_as2650[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 316.000 140.670 320.000 ;
    END
  END dso_as2650[20]
  PIN dso_as2650[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 316.000 144.350 320.000 ;
    END
  END dso_as2650[21]
  PIN dso_as2650[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 316.000 148.030 320.000 ;
    END
  END dso_as2650[22]
  PIN dso_as2650[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 316.000 151.710 320.000 ;
    END
  END dso_as2650[23]
  PIN dso_as2650[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 316.000 155.390 320.000 ;
    END
  END dso_as2650[24]
  PIN dso_as2650[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 316.000 159.070 320.000 ;
    END
  END dso_as2650[25]
  PIN dso_as2650[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 316.000 162.750 320.000 ;
    END
  END dso_as2650[26]
  PIN dso_as2650[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 316.000 74.430 320.000 ;
    END
  END dso_as2650[2]
  PIN dso_as2650[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 316.000 78.110 320.000 ;
    END
  END dso_as2650[3]
  PIN dso_as2650[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 316.000 81.790 320.000 ;
    END
  END dso_as2650[4]
  PIN dso_as2650[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 316.000 85.470 320.000 ;
    END
  END dso_as2650[5]
  PIN dso_as2650[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 316.000 89.150 320.000 ;
    END
  END dso_as2650[6]
  PIN dso_as2650[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 316.000 92.830 320.000 ;
    END
  END dso_as2650[7]
  PIN dso_as2650[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 316.000 96.510 320.000 ;
    END
  END dso_as2650[8]
  PIN dso_as2650[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 316.000 100.190 320.000 ;
    END
  END dso_as2650[9]
  PIN dso_as512512512[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END dso_as512512512[0]
  PIN dso_as512512512[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END dso_as512512512[10]
  PIN dso_as512512512[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END dso_as512512512[11]
  PIN dso_as512512512[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END dso_as512512512[12]
  PIN dso_as512512512[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END dso_as512512512[13]
  PIN dso_as512512512[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END dso_as512512512[14]
  PIN dso_as512512512[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END dso_as512512512[15]
  PIN dso_as512512512[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END dso_as512512512[16]
  PIN dso_as512512512[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END dso_as512512512[17]
  PIN dso_as512512512[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END dso_as512512512[18]
  PIN dso_as512512512[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END dso_as512512512[19]
  PIN dso_as512512512[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END dso_as512512512[1]
  PIN dso_as512512512[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END dso_as512512512[20]
  PIN dso_as512512512[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END dso_as512512512[21]
  PIN dso_as512512512[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END dso_as512512512[22]
  PIN dso_as512512512[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END dso_as512512512[23]
  PIN dso_as512512512[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END dso_as512512512[24]
  PIN dso_as512512512[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END dso_as512512512[25]
  PIN dso_as512512512[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END dso_as512512512[26]
  PIN dso_as512512512[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END dso_as512512512[27]
  PIN dso_as512512512[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END dso_as512512512[2]
  PIN dso_as512512512[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END dso_as512512512[3]
  PIN dso_as512512512[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END dso_as512512512[4]
  PIN dso_as512512512[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END dso_as512512512[5]
  PIN dso_as512512512[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END dso_as512512512[6]
  PIN dso_as512512512[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END dso_as512512512[7]
  PIN dso_as512512512[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END dso_as512512512[8]
  PIN dso_as512512512[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END dso_as512512512[9]
  PIN dso_as5401[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 316.000 166.430 320.000 ;
    END
  END dso_as5401[0]
  PIN dso_as5401[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 316.000 203.230 320.000 ;
    END
  END dso_as5401[10]
  PIN dso_as5401[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 316.000 206.910 320.000 ;
    END
  END dso_as5401[11]
  PIN dso_as5401[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 316.000 210.590 320.000 ;
    END
  END dso_as5401[12]
  PIN dso_as5401[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 316.000 214.270 320.000 ;
    END
  END dso_as5401[13]
  PIN dso_as5401[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 316.000 217.950 320.000 ;
    END
  END dso_as5401[14]
  PIN dso_as5401[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 316.000 221.630 320.000 ;
    END
  END dso_as5401[15]
  PIN dso_as5401[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 316.000 225.310 320.000 ;
    END
  END dso_as5401[16]
  PIN dso_as5401[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 316.000 228.990 320.000 ;
    END
  END dso_as5401[17]
  PIN dso_as5401[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 316.000 232.670 320.000 ;
    END
  END dso_as5401[18]
  PIN dso_as5401[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 316.000 236.350 320.000 ;
    END
  END dso_as5401[19]
  PIN dso_as5401[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 316.000 170.110 320.000 ;
    END
  END dso_as5401[1]
  PIN dso_as5401[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 316.000 240.030 320.000 ;
    END
  END dso_as5401[20]
  PIN dso_as5401[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 316.000 243.710 320.000 ;
    END
  END dso_as5401[21]
  PIN dso_as5401[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 316.000 247.390 320.000 ;
    END
  END dso_as5401[22]
  PIN dso_as5401[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 316.000 251.070 320.000 ;
    END
  END dso_as5401[23]
  PIN dso_as5401[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 316.000 254.750 320.000 ;
    END
  END dso_as5401[24]
  PIN dso_as5401[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 316.000 258.430 320.000 ;
    END
  END dso_as5401[25]
  PIN dso_as5401[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 316.000 262.110 320.000 ;
    END
  END dso_as5401[26]
  PIN dso_as5401[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 316.000 173.790 320.000 ;
    END
  END dso_as5401[2]
  PIN dso_as5401[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 316.000 177.470 320.000 ;
    END
  END dso_as5401[3]
  PIN dso_as5401[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 316.000 181.150 320.000 ;
    END
  END dso_as5401[4]
  PIN dso_as5401[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 316.000 184.830 320.000 ;
    END
  END dso_as5401[5]
  PIN dso_as5401[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 316.000 188.510 320.000 ;
    END
  END dso_as5401[6]
  PIN dso_as5401[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 316.000 192.190 320.000 ;
    END
  END dso_as5401[7]
  PIN dso_as5401[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 316.000 195.870 320.000 ;
    END
  END dso_as5401[8]
  PIN dso_as5401[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 316.000 199.550 320.000 ;
    END
  END dso_as5401[9]
  PIN dso_counter[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 282.920 300.000 283.520 ;
    END
  END dso_counter[0]
  PIN dso_counter[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 310.120 300.000 310.720 ;
    END
  END dso_counter[10]
  PIN dso_counter[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 312.840 300.000 313.440 ;
    END
  END dso_counter[11]
  PIN dso_counter[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 285.640 300.000 286.240 ;
    END
  END dso_counter[1]
  PIN dso_counter[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 288.360 300.000 288.960 ;
    END
  END dso_counter[2]
  PIN dso_counter[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 291.080 300.000 291.680 ;
    END
  END dso_counter[3]
  PIN dso_counter[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 293.800 300.000 294.400 ;
    END
  END dso_counter[4]
  PIN dso_counter[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 296.520 300.000 297.120 ;
    END
  END dso_counter[5]
  PIN dso_counter[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 299.240 300.000 299.840 ;
    END
  END dso_counter[6]
  PIN dso_counter[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 301.960 300.000 302.560 ;
    END
  END dso_counter[7]
  PIN dso_counter[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 304.680 300.000 305.280 ;
    END
  END dso_counter[8]
  PIN dso_counter[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 307.400 300.000 308.000 ;
    END
  END dso_counter[9]
  PIN dso_diceroll[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 316.000 33.950 320.000 ;
    END
  END dso_diceroll[0]
  PIN dso_diceroll[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 316.000 37.630 320.000 ;
    END
  END dso_diceroll[1]
  PIN dso_diceroll[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 316.000 41.310 320.000 ;
    END
  END dso_diceroll[2]
  PIN dso_diceroll[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 316.000 44.990 320.000 ;
    END
  END dso_diceroll[3]
  PIN dso_diceroll[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 316.000 48.670 320.000 ;
    END
  END dso_diceroll[4]
  PIN dso_diceroll[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 316.000 52.350 320.000 ;
    END
  END dso_diceroll[5]
  PIN dso_diceroll[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 316.000 56.030 320.000 ;
    END
  END dso_diceroll[6]
  PIN dso_diceroll[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 316.000 59.710 320.000 ;
    END
  END dso_diceroll[7]
  PIN dso_mc14500[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END dso_mc14500[0]
  PIN dso_mc14500[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END dso_mc14500[1]
  PIN dso_mc14500[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END dso_mc14500[2]
  PIN dso_mc14500[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END dso_mc14500[3]
  PIN dso_mc14500[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END dso_mc14500[4]
  PIN dso_mc14500[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END dso_mc14500[5]
  PIN dso_mc14500[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END dso_mc14500[6]
  PIN dso_mc14500[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END dso_mc14500[7]
  PIN dso_mc14500[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END dso_mc14500[8]
  PIN dso_multiplier[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 316.000 4.510 320.000 ;
    END
  END dso_multiplier[0]
  PIN dso_multiplier[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 316.000 8.190 320.000 ;
    END
  END dso_multiplier[1]
  PIN dso_multiplier[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 316.000 11.870 320.000 ;
    END
  END dso_multiplier[2]
  PIN dso_multiplier[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 316.000 15.550 320.000 ;
    END
  END dso_multiplier[3]
  PIN dso_multiplier[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 316.000 19.230 320.000 ;
    END
  END dso_multiplier[4]
  PIN dso_multiplier[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 316.000 22.910 320.000 ;
    END
  END dso_multiplier[5]
  PIN dso_multiplier[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 316.000 26.590 320.000 ;
    END
  END dso_multiplier[6]
  PIN dso_multiplier[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 316.000 30.270 320.000 ;
    END
  END dso_multiplier[7]
  PIN dso_posit[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END dso_posit[0]
  PIN dso_posit[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END dso_posit[1]
  PIN dso_posit[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END dso_posit[2]
  PIN dso_posit[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END dso_posit[3]
  PIN dso_tbb1143[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END dso_tbb1143[0]
  PIN dso_tbb1143[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END dso_tbb1143[1]
  PIN dso_tbb1143[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END dso_tbb1143[2]
  PIN dso_tbb1143[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END dso_tbb1143[3]
  PIN dso_tbb1143[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END dso_tbb1143[4]
  PIN dso_tbb1143[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END dso_tbb1143[5]
  PIN dso_tbb1143[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END dso_tbb1143[6]
  PIN dso_tbb1143[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END dso_tbb1143[7]
  PIN dso_tune
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END dso_tune
  PIN dso_vgatest[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END dso_vgatest[0]
  PIN dso_vgatest[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END dso_vgatest[1]
  PIN dso_vgatest[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END dso_vgatest[2]
  PIN dso_vgatest[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END dso_vgatest[3]
  PIN dso_vgatest[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END dso_vgatest[4]
  PIN dso_vgatest[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 0.000 271.310 4.000 ;
    END
  END dso_vgatest[5]
  PIN dso_vgatest[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END dso_vgatest[6]
  PIN dso_vgatest[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END dso_vgatest[7]
  PIN dso_vgatest[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END dso_vgatest[8]
  PIN dso_vgatest[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END dso_vgatest[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END io_out[9]
  PIN oeb_6502
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END oeb_6502
  PIN oeb_as1802
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END oeb_as1802
  PIN oeb_as2650
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 316.000 63.390 320.000 ;
    END
  END oeb_as2650
  PIN oeb_as512512512
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END oeb_as512512512
  PIN oeb_as5401
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 316.000 265.790 320.000 ;
    END
  END oeb_as5401
  PIN oeb_mc14500
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END oeb_mc14500
  PIN rst_6502
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END rst_6502
  PIN rst_LCD
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END rst_LCD
  PIN rst_as1802
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END rst_as1802
  PIN rst_as2650
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END rst_as2650
  PIN rst_as512512512
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END rst_as512512512
  PIN rst_as5401
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END rst_as5401
  PIN rst_counter
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END rst_counter
  PIN rst_diceroll
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END rst_diceroll
  PIN rst_mc14500
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END rst_mc14500
  PIN rst_posit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END rst_posit
  PIN rst_tbb1143
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END rst_tbb1143
  PIN rst_tune
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END rst_tune
  PIN rst_vgatest
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END rst_vgatest
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 307.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 307.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 307.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 307.600 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 5.480 300.000 6.080 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.200 300.000 8.800 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.920 300.000 11.520 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 21.800 300.000 22.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 103.400 300.000 104.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.560 300.000 112.160 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 119.720 300.000 120.320 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 127.880 300.000 128.480 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.040 300.000 136.640 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 144.200 300.000 144.800 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 152.360 300.000 152.960 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 160.520 300.000 161.120 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 168.680 300.000 169.280 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 176.840 300.000 177.440 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 29.960 300.000 30.560 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 185.000 300.000 185.600 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 193.160 300.000 193.760 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.320 300.000 201.920 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 209.480 300.000 210.080 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 217.640 300.000 218.240 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 225.800 300.000 226.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 233.960 300.000 234.560 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 242.120 300.000 242.720 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 250.280 300.000 250.880 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.440 300.000 259.040 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 38.120 300.000 38.720 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.600 300.000 267.200 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 274.760 300.000 275.360 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 46.280 300.000 46.880 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 54.440 300.000 55.040 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 62.600 300.000 63.200 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 70.760 300.000 71.360 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 78.920 300.000 79.520 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 87.080 300.000 87.680 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 95.240 300.000 95.840 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 13.640 300.000 14.240 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 24.520 300.000 25.120 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 106.120 300.000 106.720 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 114.280 300.000 114.880 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.440 300.000 123.040 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 130.600 300.000 131.200 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 138.760 300.000 139.360 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.920 300.000 147.520 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 155.080 300.000 155.680 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 163.240 300.000 163.840 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 171.400 300.000 172.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.560 300.000 180.160 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 32.680 300.000 33.280 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 187.720 300.000 188.320 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 195.880 300.000 196.480 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 204.040 300.000 204.640 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 212.200 300.000 212.800 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 220.360 300.000 220.960 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 228.520 300.000 229.120 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 236.680 300.000 237.280 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 244.840 300.000 245.440 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 253.000 300.000 253.600 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 261.160 300.000 261.760 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 40.840 300.000 41.440 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 269.320 300.000 269.920 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 277.480 300.000 278.080 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 49.000 300.000 49.600 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.160 300.000 57.760 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.320 300.000 65.920 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.480 300.000 74.080 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 81.640 300.000 82.240 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 89.800 300.000 90.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 97.960 300.000 98.560 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 27.240 300.000 27.840 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 108.840 300.000 109.440 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 117.000 300.000 117.600 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.160 300.000 125.760 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 133.320 300.000 133.920 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.480 300.000 142.080 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 149.640 300.000 150.240 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 157.800 300.000 158.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 165.960 300.000 166.560 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 174.120 300.000 174.720 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.280 300.000 182.880 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 35.400 300.000 36.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.440 300.000 191.040 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 198.600 300.000 199.200 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 206.760 300.000 207.360 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 214.920 300.000 215.520 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 223.080 300.000 223.680 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 231.240 300.000 231.840 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 239.400 300.000 240.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 247.560 300.000 248.160 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.720 300.000 256.320 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 263.880 300.000 264.480 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 43.560 300.000 44.160 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 272.040 300.000 272.640 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 280.200 300.000 280.800 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 51.720 300.000 52.320 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 59.880 300.000 60.480 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 68.040 300.000 68.640 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.200 300.000 76.800 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 84.360 300.000 84.960 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 92.520 300.000 93.120 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 100.680 300.000 101.280 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.360 300.000 16.960 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 19.080 300.000 19.680 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 307.445 ;
      LAYER met1 ;
        RECT 4.210 0.380 298.010 316.500 ;
      LAYER met2 ;
        RECT 4.790 315.720 7.630 316.610 ;
        RECT 8.470 315.720 11.310 316.610 ;
        RECT 12.150 315.720 14.990 316.610 ;
        RECT 15.830 315.720 18.670 316.610 ;
        RECT 19.510 315.720 22.350 316.610 ;
        RECT 23.190 315.720 26.030 316.610 ;
        RECT 26.870 315.720 29.710 316.610 ;
        RECT 30.550 315.720 33.390 316.610 ;
        RECT 34.230 315.720 37.070 316.610 ;
        RECT 37.910 315.720 40.750 316.610 ;
        RECT 41.590 315.720 44.430 316.610 ;
        RECT 45.270 315.720 48.110 316.610 ;
        RECT 48.950 315.720 51.790 316.610 ;
        RECT 52.630 315.720 55.470 316.610 ;
        RECT 56.310 315.720 59.150 316.610 ;
        RECT 59.990 315.720 62.830 316.610 ;
        RECT 63.670 315.720 66.510 316.610 ;
        RECT 67.350 315.720 70.190 316.610 ;
        RECT 71.030 315.720 73.870 316.610 ;
        RECT 74.710 315.720 77.550 316.610 ;
        RECT 78.390 315.720 81.230 316.610 ;
        RECT 82.070 315.720 84.910 316.610 ;
        RECT 85.750 315.720 88.590 316.610 ;
        RECT 89.430 315.720 92.270 316.610 ;
        RECT 93.110 315.720 95.950 316.610 ;
        RECT 96.790 315.720 99.630 316.610 ;
        RECT 100.470 315.720 103.310 316.610 ;
        RECT 104.150 315.720 106.990 316.610 ;
        RECT 107.830 315.720 110.670 316.610 ;
        RECT 111.510 315.720 114.350 316.610 ;
        RECT 115.190 315.720 118.030 316.610 ;
        RECT 118.870 315.720 121.710 316.610 ;
        RECT 122.550 315.720 125.390 316.610 ;
        RECT 126.230 315.720 129.070 316.610 ;
        RECT 129.910 315.720 132.750 316.610 ;
        RECT 133.590 315.720 136.430 316.610 ;
        RECT 137.270 315.720 140.110 316.610 ;
        RECT 140.950 315.720 143.790 316.610 ;
        RECT 144.630 315.720 147.470 316.610 ;
        RECT 148.310 315.720 151.150 316.610 ;
        RECT 151.990 315.720 154.830 316.610 ;
        RECT 155.670 315.720 158.510 316.610 ;
        RECT 159.350 315.720 162.190 316.610 ;
        RECT 163.030 315.720 165.870 316.610 ;
        RECT 166.710 315.720 169.550 316.610 ;
        RECT 170.390 315.720 173.230 316.610 ;
        RECT 174.070 315.720 176.910 316.610 ;
        RECT 177.750 315.720 180.590 316.610 ;
        RECT 181.430 315.720 184.270 316.610 ;
        RECT 185.110 315.720 187.950 316.610 ;
        RECT 188.790 315.720 191.630 316.610 ;
        RECT 192.470 315.720 195.310 316.610 ;
        RECT 196.150 315.720 198.990 316.610 ;
        RECT 199.830 315.720 202.670 316.610 ;
        RECT 203.510 315.720 206.350 316.610 ;
        RECT 207.190 315.720 210.030 316.610 ;
        RECT 210.870 315.720 213.710 316.610 ;
        RECT 214.550 315.720 217.390 316.610 ;
        RECT 218.230 315.720 221.070 316.610 ;
        RECT 221.910 315.720 224.750 316.610 ;
        RECT 225.590 315.720 228.430 316.610 ;
        RECT 229.270 315.720 232.110 316.610 ;
        RECT 232.950 315.720 235.790 316.610 ;
        RECT 236.630 315.720 239.470 316.610 ;
        RECT 240.310 315.720 243.150 316.610 ;
        RECT 243.990 315.720 246.830 316.610 ;
        RECT 247.670 315.720 250.510 316.610 ;
        RECT 251.350 315.720 254.190 316.610 ;
        RECT 255.030 315.720 257.870 316.610 ;
        RECT 258.710 315.720 261.550 316.610 ;
        RECT 262.390 315.720 265.230 316.610 ;
        RECT 266.070 315.720 268.910 316.610 ;
        RECT 269.750 315.720 272.590 316.610 ;
        RECT 273.430 315.720 276.270 316.610 ;
        RECT 277.110 315.720 279.950 316.610 ;
        RECT 280.790 315.720 283.630 316.610 ;
        RECT 284.470 315.720 287.310 316.610 ;
        RECT 288.150 315.720 290.990 316.610 ;
        RECT 291.830 315.720 294.670 316.610 ;
        RECT 295.510 315.720 297.980 316.610 ;
        RECT 4.240 4.280 297.980 315.720 ;
        RECT 4.240 0.350 22.350 4.280 ;
        RECT 23.190 0.350 23.730 4.280 ;
        RECT 24.570 0.350 25.110 4.280 ;
        RECT 25.950 0.350 26.490 4.280 ;
        RECT 27.330 0.350 27.870 4.280 ;
        RECT 28.710 0.350 29.250 4.280 ;
        RECT 30.090 0.350 30.630 4.280 ;
        RECT 31.470 0.350 32.010 4.280 ;
        RECT 32.850 0.350 33.390 4.280 ;
        RECT 34.230 0.350 34.770 4.280 ;
        RECT 35.610 0.350 36.150 4.280 ;
        RECT 36.990 0.350 37.530 4.280 ;
        RECT 38.370 0.350 38.910 4.280 ;
        RECT 39.750 0.350 40.290 4.280 ;
        RECT 41.130 0.350 41.670 4.280 ;
        RECT 42.510 0.350 43.050 4.280 ;
        RECT 43.890 0.350 44.430 4.280 ;
        RECT 45.270 0.350 45.810 4.280 ;
        RECT 46.650 0.350 47.190 4.280 ;
        RECT 48.030 0.350 48.570 4.280 ;
        RECT 49.410 0.350 49.950 4.280 ;
        RECT 50.790 0.350 51.330 4.280 ;
        RECT 52.170 0.350 52.710 4.280 ;
        RECT 53.550 0.350 54.090 4.280 ;
        RECT 54.930 0.350 55.470 4.280 ;
        RECT 56.310 0.350 56.850 4.280 ;
        RECT 57.690 0.350 58.230 4.280 ;
        RECT 59.070 0.350 59.610 4.280 ;
        RECT 60.450 0.350 60.990 4.280 ;
        RECT 61.830 0.350 62.370 4.280 ;
        RECT 63.210 0.350 63.750 4.280 ;
        RECT 64.590 0.350 65.130 4.280 ;
        RECT 65.970 0.350 66.510 4.280 ;
        RECT 67.350 0.350 67.890 4.280 ;
        RECT 68.730 0.350 69.270 4.280 ;
        RECT 70.110 0.350 70.650 4.280 ;
        RECT 71.490 0.350 72.030 4.280 ;
        RECT 72.870 0.350 73.410 4.280 ;
        RECT 74.250 0.350 74.790 4.280 ;
        RECT 75.630 0.350 76.170 4.280 ;
        RECT 77.010 0.350 77.550 4.280 ;
        RECT 78.390 0.350 78.930 4.280 ;
        RECT 79.770 0.350 80.310 4.280 ;
        RECT 81.150 0.350 81.690 4.280 ;
        RECT 82.530 0.350 83.070 4.280 ;
        RECT 83.910 0.350 84.450 4.280 ;
        RECT 85.290 0.350 85.830 4.280 ;
        RECT 86.670 0.350 87.210 4.280 ;
        RECT 88.050 0.350 88.590 4.280 ;
        RECT 89.430 0.350 89.970 4.280 ;
        RECT 90.810 0.350 91.350 4.280 ;
        RECT 92.190 0.350 92.730 4.280 ;
        RECT 93.570 0.350 94.110 4.280 ;
        RECT 94.950 0.350 95.490 4.280 ;
        RECT 96.330 0.350 96.870 4.280 ;
        RECT 97.710 0.350 98.250 4.280 ;
        RECT 99.090 0.350 99.630 4.280 ;
        RECT 100.470 0.350 101.010 4.280 ;
        RECT 101.850 0.350 102.390 4.280 ;
        RECT 103.230 0.350 103.770 4.280 ;
        RECT 104.610 0.350 105.150 4.280 ;
        RECT 105.990 0.350 106.530 4.280 ;
        RECT 107.370 0.350 107.910 4.280 ;
        RECT 108.750 0.350 109.290 4.280 ;
        RECT 110.130 0.350 110.670 4.280 ;
        RECT 111.510 0.350 112.050 4.280 ;
        RECT 112.890 0.350 113.430 4.280 ;
        RECT 114.270 0.350 114.810 4.280 ;
        RECT 115.650 0.350 116.190 4.280 ;
        RECT 117.030 0.350 117.570 4.280 ;
        RECT 118.410 0.350 118.950 4.280 ;
        RECT 119.790 0.350 120.330 4.280 ;
        RECT 121.170 0.350 121.710 4.280 ;
        RECT 122.550 0.350 123.090 4.280 ;
        RECT 123.930 0.350 124.470 4.280 ;
        RECT 125.310 0.350 125.850 4.280 ;
        RECT 126.690 0.350 127.230 4.280 ;
        RECT 128.070 0.350 128.610 4.280 ;
        RECT 129.450 0.350 129.990 4.280 ;
        RECT 130.830 0.350 131.370 4.280 ;
        RECT 132.210 0.350 132.750 4.280 ;
        RECT 133.590 0.350 134.130 4.280 ;
        RECT 134.970 0.350 135.510 4.280 ;
        RECT 136.350 0.350 136.890 4.280 ;
        RECT 137.730 0.350 138.270 4.280 ;
        RECT 139.110 0.350 139.650 4.280 ;
        RECT 140.490 0.350 141.030 4.280 ;
        RECT 141.870 0.350 142.410 4.280 ;
        RECT 143.250 0.350 143.790 4.280 ;
        RECT 144.630 0.350 145.170 4.280 ;
        RECT 146.010 0.350 146.550 4.280 ;
        RECT 147.390 0.350 147.930 4.280 ;
        RECT 148.770 0.350 149.310 4.280 ;
        RECT 150.150 0.350 150.690 4.280 ;
        RECT 151.530 0.350 152.070 4.280 ;
        RECT 152.910 0.350 153.450 4.280 ;
        RECT 154.290 0.350 154.830 4.280 ;
        RECT 155.670 0.350 156.210 4.280 ;
        RECT 157.050 0.350 157.590 4.280 ;
        RECT 158.430 0.350 158.970 4.280 ;
        RECT 159.810 0.350 160.350 4.280 ;
        RECT 161.190 0.350 161.730 4.280 ;
        RECT 162.570 0.350 163.110 4.280 ;
        RECT 163.950 0.350 164.490 4.280 ;
        RECT 165.330 0.350 165.870 4.280 ;
        RECT 166.710 0.350 167.250 4.280 ;
        RECT 168.090 0.350 168.630 4.280 ;
        RECT 169.470 0.350 170.010 4.280 ;
        RECT 170.850 0.350 171.390 4.280 ;
        RECT 172.230 0.350 172.770 4.280 ;
        RECT 173.610 0.350 174.150 4.280 ;
        RECT 174.990 0.350 175.530 4.280 ;
        RECT 176.370 0.350 176.910 4.280 ;
        RECT 177.750 0.350 178.290 4.280 ;
        RECT 179.130 0.350 179.670 4.280 ;
        RECT 180.510 0.350 181.050 4.280 ;
        RECT 181.890 0.350 182.430 4.280 ;
        RECT 183.270 0.350 183.810 4.280 ;
        RECT 184.650 0.350 185.190 4.280 ;
        RECT 186.030 0.350 186.570 4.280 ;
        RECT 187.410 0.350 187.950 4.280 ;
        RECT 188.790 0.350 189.330 4.280 ;
        RECT 190.170 0.350 190.710 4.280 ;
        RECT 191.550 0.350 192.090 4.280 ;
        RECT 192.930 0.350 193.470 4.280 ;
        RECT 194.310 0.350 194.850 4.280 ;
        RECT 195.690 0.350 196.230 4.280 ;
        RECT 197.070 0.350 197.610 4.280 ;
        RECT 198.450 0.350 198.990 4.280 ;
        RECT 199.830 0.350 200.370 4.280 ;
        RECT 201.210 0.350 201.750 4.280 ;
        RECT 202.590 0.350 203.130 4.280 ;
        RECT 203.970 0.350 204.510 4.280 ;
        RECT 205.350 0.350 205.890 4.280 ;
        RECT 206.730 0.350 207.270 4.280 ;
        RECT 208.110 0.350 208.650 4.280 ;
        RECT 209.490 0.350 210.030 4.280 ;
        RECT 210.870 0.350 211.410 4.280 ;
        RECT 212.250 0.350 212.790 4.280 ;
        RECT 213.630 0.350 214.170 4.280 ;
        RECT 215.010 0.350 215.550 4.280 ;
        RECT 216.390 0.350 216.930 4.280 ;
        RECT 217.770 0.350 218.310 4.280 ;
        RECT 219.150 0.350 219.690 4.280 ;
        RECT 220.530 0.350 221.070 4.280 ;
        RECT 221.910 0.350 222.450 4.280 ;
        RECT 223.290 0.350 223.830 4.280 ;
        RECT 224.670 0.350 225.210 4.280 ;
        RECT 226.050 0.350 226.590 4.280 ;
        RECT 227.430 0.350 227.970 4.280 ;
        RECT 228.810 0.350 229.350 4.280 ;
        RECT 230.190 0.350 230.730 4.280 ;
        RECT 231.570 0.350 232.110 4.280 ;
        RECT 232.950 0.350 233.490 4.280 ;
        RECT 234.330 0.350 234.870 4.280 ;
        RECT 235.710 0.350 236.250 4.280 ;
        RECT 237.090 0.350 237.630 4.280 ;
        RECT 238.470 0.350 239.010 4.280 ;
        RECT 239.850 0.350 240.390 4.280 ;
        RECT 241.230 0.350 241.770 4.280 ;
        RECT 242.610 0.350 243.150 4.280 ;
        RECT 243.990 0.350 244.530 4.280 ;
        RECT 245.370 0.350 245.910 4.280 ;
        RECT 246.750 0.350 247.290 4.280 ;
        RECT 248.130 0.350 248.670 4.280 ;
        RECT 249.510 0.350 250.050 4.280 ;
        RECT 250.890 0.350 251.430 4.280 ;
        RECT 252.270 0.350 252.810 4.280 ;
        RECT 253.650 0.350 254.190 4.280 ;
        RECT 255.030 0.350 255.570 4.280 ;
        RECT 256.410 0.350 256.950 4.280 ;
        RECT 257.790 0.350 258.330 4.280 ;
        RECT 259.170 0.350 259.710 4.280 ;
        RECT 260.550 0.350 261.090 4.280 ;
        RECT 261.930 0.350 262.470 4.280 ;
        RECT 263.310 0.350 263.850 4.280 ;
        RECT 264.690 0.350 265.230 4.280 ;
        RECT 266.070 0.350 266.610 4.280 ;
        RECT 267.450 0.350 267.990 4.280 ;
        RECT 268.830 0.350 269.370 4.280 ;
        RECT 270.210 0.350 270.750 4.280 ;
        RECT 271.590 0.350 272.130 4.280 ;
        RECT 272.970 0.350 273.510 4.280 ;
        RECT 274.350 0.350 274.890 4.280 ;
        RECT 275.730 0.350 276.270 4.280 ;
        RECT 277.110 0.350 297.980 4.280 ;
      LAYER met3 ;
        RECT 4.000 312.440 295.600 313.305 ;
        RECT 4.000 311.120 296.000 312.440 ;
        RECT 4.000 309.760 295.600 311.120 ;
        RECT 4.400 309.720 295.600 309.760 ;
        RECT 4.400 308.400 296.000 309.720 ;
        RECT 4.400 308.360 295.600 308.400 ;
        RECT 4.000 307.000 295.600 308.360 ;
        RECT 4.000 306.360 296.000 307.000 ;
        RECT 4.400 305.680 296.000 306.360 ;
        RECT 4.400 304.960 295.600 305.680 ;
        RECT 4.000 304.280 295.600 304.960 ;
        RECT 4.000 302.960 296.000 304.280 ;
        RECT 4.400 301.560 295.600 302.960 ;
        RECT 4.000 300.240 296.000 301.560 ;
        RECT 4.000 299.560 295.600 300.240 ;
        RECT 4.400 298.840 295.600 299.560 ;
        RECT 4.400 298.160 296.000 298.840 ;
        RECT 4.000 297.520 296.000 298.160 ;
        RECT 4.000 296.160 295.600 297.520 ;
        RECT 4.400 296.120 295.600 296.160 ;
        RECT 4.400 294.800 296.000 296.120 ;
        RECT 4.400 294.760 295.600 294.800 ;
        RECT 4.000 293.400 295.600 294.760 ;
        RECT 4.000 292.760 296.000 293.400 ;
        RECT 4.400 292.080 296.000 292.760 ;
        RECT 4.400 291.360 295.600 292.080 ;
        RECT 4.000 290.680 295.600 291.360 ;
        RECT 4.000 289.360 296.000 290.680 ;
        RECT 4.400 287.960 295.600 289.360 ;
        RECT 4.000 286.640 296.000 287.960 ;
        RECT 4.000 285.960 295.600 286.640 ;
        RECT 4.400 285.240 295.600 285.960 ;
        RECT 4.400 284.560 296.000 285.240 ;
        RECT 4.000 283.920 296.000 284.560 ;
        RECT 4.000 282.560 295.600 283.920 ;
        RECT 4.400 282.520 295.600 282.560 ;
        RECT 4.400 281.200 296.000 282.520 ;
        RECT 4.400 281.160 295.600 281.200 ;
        RECT 4.000 279.800 295.600 281.160 ;
        RECT 4.000 279.160 296.000 279.800 ;
        RECT 4.400 278.480 296.000 279.160 ;
        RECT 4.400 277.760 295.600 278.480 ;
        RECT 4.000 277.080 295.600 277.760 ;
        RECT 4.000 275.760 296.000 277.080 ;
        RECT 4.400 274.360 295.600 275.760 ;
        RECT 4.000 273.040 296.000 274.360 ;
        RECT 4.000 272.360 295.600 273.040 ;
        RECT 4.400 271.640 295.600 272.360 ;
        RECT 4.400 270.960 296.000 271.640 ;
        RECT 4.000 270.320 296.000 270.960 ;
        RECT 4.000 268.960 295.600 270.320 ;
        RECT 4.400 268.920 295.600 268.960 ;
        RECT 4.400 267.600 296.000 268.920 ;
        RECT 4.400 267.560 295.600 267.600 ;
        RECT 4.000 266.200 295.600 267.560 ;
        RECT 4.000 265.560 296.000 266.200 ;
        RECT 4.400 264.880 296.000 265.560 ;
        RECT 4.400 264.160 295.600 264.880 ;
        RECT 4.000 263.480 295.600 264.160 ;
        RECT 4.000 262.160 296.000 263.480 ;
        RECT 4.400 260.760 295.600 262.160 ;
        RECT 4.000 259.440 296.000 260.760 ;
        RECT 4.000 258.760 295.600 259.440 ;
        RECT 4.400 258.040 295.600 258.760 ;
        RECT 4.400 257.360 296.000 258.040 ;
        RECT 4.000 256.720 296.000 257.360 ;
        RECT 4.000 255.360 295.600 256.720 ;
        RECT 4.400 255.320 295.600 255.360 ;
        RECT 4.400 254.000 296.000 255.320 ;
        RECT 4.400 253.960 295.600 254.000 ;
        RECT 4.000 252.600 295.600 253.960 ;
        RECT 4.000 251.960 296.000 252.600 ;
        RECT 4.400 251.280 296.000 251.960 ;
        RECT 4.400 250.560 295.600 251.280 ;
        RECT 4.000 249.880 295.600 250.560 ;
        RECT 4.000 248.560 296.000 249.880 ;
        RECT 4.400 247.160 295.600 248.560 ;
        RECT 4.000 245.840 296.000 247.160 ;
        RECT 4.000 245.160 295.600 245.840 ;
        RECT 4.400 244.440 295.600 245.160 ;
        RECT 4.400 243.760 296.000 244.440 ;
        RECT 4.000 243.120 296.000 243.760 ;
        RECT 4.000 241.760 295.600 243.120 ;
        RECT 4.400 241.720 295.600 241.760 ;
        RECT 4.400 240.400 296.000 241.720 ;
        RECT 4.400 240.360 295.600 240.400 ;
        RECT 4.000 239.000 295.600 240.360 ;
        RECT 4.000 238.360 296.000 239.000 ;
        RECT 4.400 237.680 296.000 238.360 ;
        RECT 4.400 236.960 295.600 237.680 ;
        RECT 4.000 236.280 295.600 236.960 ;
        RECT 4.000 234.960 296.000 236.280 ;
        RECT 4.400 233.560 295.600 234.960 ;
        RECT 4.000 232.240 296.000 233.560 ;
        RECT 4.000 231.560 295.600 232.240 ;
        RECT 4.400 230.840 295.600 231.560 ;
        RECT 4.400 230.160 296.000 230.840 ;
        RECT 4.000 229.520 296.000 230.160 ;
        RECT 4.000 228.160 295.600 229.520 ;
        RECT 4.400 228.120 295.600 228.160 ;
        RECT 4.400 226.800 296.000 228.120 ;
        RECT 4.400 226.760 295.600 226.800 ;
        RECT 4.000 225.400 295.600 226.760 ;
        RECT 4.000 224.760 296.000 225.400 ;
        RECT 4.400 224.080 296.000 224.760 ;
        RECT 4.400 223.360 295.600 224.080 ;
        RECT 4.000 222.680 295.600 223.360 ;
        RECT 4.000 221.360 296.000 222.680 ;
        RECT 4.400 219.960 295.600 221.360 ;
        RECT 4.000 218.640 296.000 219.960 ;
        RECT 4.000 217.960 295.600 218.640 ;
        RECT 4.400 217.240 295.600 217.960 ;
        RECT 4.400 216.560 296.000 217.240 ;
        RECT 4.000 215.920 296.000 216.560 ;
        RECT 4.000 214.560 295.600 215.920 ;
        RECT 4.400 214.520 295.600 214.560 ;
        RECT 4.400 213.200 296.000 214.520 ;
        RECT 4.400 213.160 295.600 213.200 ;
        RECT 4.000 211.800 295.600 213.160 ;
        RECT 4.000 211.160 296.000 211.800 ;
        RECT 4.400 210.480 296.000 211.160 ;
        RECT 4.400 209.760 295.600 210.480 ;
        RECT 4.000 209.080 295.600 209.760 ;
        RECT 4.000 207.760 296.000 209.080 ;
        RECT 4.400 206.360 295.600 207.760 ;
        RECT 4.000 205.040 296.000 206.360 ;
        RECT 4.000 204.360 295.600 205.040 ;
        RECT 4.400 203.640 295.600 204.360 ;
        RECT 4.400 202.960 296.000 203.640 ;
        RECT 4.000 202.320 296.000 202.960 ;
        RECT 4.000 200.960 295.600 202.320 ;
        RECT 4.400 200.920 295.600 200.960 ;
        RECT 4.400 199.600 296.000 200.920 ;
        RECT 4.400 199.560 295.600 199.600 ;
        RECT 4.000 198.200 295.600 199.560 ;
        RECT 4.000 197.560 296.000 198.200 ;
        RECT 4.400 196.880 296.000 197.560 ;
        RECT 4.400 196.160 295.600 196.880 ;
        RECT 4.000 195.480 295.600 196.160 ;
        RECT 4.000 194.160 296.000 195.480 ;
        RECT 4.400 192.760 295.600 194.160 ;
        RECT 4.000 191.440 296.000 192.760 ;
        RECT 4.000 190.760 295.600 191.440 ;
        RECT 4.400 190.040 295.600 190.760 ;
        RECT 4.400 189.360 296.000 190.040 ;
        RECT 4.000 188.720 296.000 189.360 ;
        RECT 4.000 187.360 295.600 188.720 ;
        RECT 4.400 187.320 295.600 187.360 ;
        RECT 4.400 186.000 296.000 187.320 ;
        RECT 4.400 185.960 295.600 186.000 ;
        RECT 4.000 184.600 295.600 185.960 ;
        RECT 4.000 183.960 296.000 184.600 ;
        RECT 4.400 183.280 296.000 183.960 ;
        RECT 4.400 182.560 295.600 183.280 ;
        RECT 4.000 181.880 295.600 182.560 ;
        RECT 4.000 180.560 296.000 181.880 ;
        RECT 4.400 179.160 295.600 180.560 ;
        RECT 4.000 177.840 296.000 179.160 ;
        RECT 4.000 177.160 295.600 177.840 ;
        RECT 4.400 176.440 295.600 177.160 ;
        RECT 4.400 175.760 296.000 176.440 ;
        RECT 4.000 175.120 296.000 175.760 ;
        RECT 4.000 173.760 295.600 175.120 ;
        RECT 4.400 173.720 295.600 173.760 ;
        RECT 4.400 172.400 296.000 173.720 ;
        RECT 4.400 172.360 295.600 172.400 ;
        RECT 4.000 171.000 295.600 172.360 ;
        RECT 4.000 170.360 296.000 171.000 ;
        RECT 4.400 169.680 296.000 170.360 ;
        RECT 4.400 168.960 295.600 169.680 ;
        RECT 4.000 168.280 295.600 168.960 ;
        RECT 4.000 166.960 296.000 168.280 ;
        RECT 4.400 165.560 295.600 166.960 ;
        RECT 4.000 164.240 296.000 165.560 ;
        RECT 4.000 163.560 295.600 164.240 ;
        RECT 4.400 162.840 295.600 163.560 ;
        RECT 4.400 162.160 296.000 162.840 ;
        RECT 4.000 161.520 296.000 162.160 ;
        RECT 4.000 160.160 295.600 161.520 ;
        RECT 4.400 160.120 295.600 160.160 ;
        RECT 4.400 158.800 296.000 160.120 ;
        RECT 4.400 158.760 295.600 158.800 ;
        RECT 4.000 157.400 295.600 158.760 ;
        RECT 4.000 156.760 296.000 157.400 ;
        RECT 4.400 156.080 296.000 156.760 ;
        RECT 4.400 155.360 295.600 156.080 ;
        RECT 4.000 154.680 295.600 155.360 ;
        RECT 4.000 153.360 296.000 154.680 ;
        RECT 4.400 151.960 295.600 153.360 ;
        RECT 4.000 150.640 296.000 151.960 ;
        RECT 4.000 149.960 295.600 150.640 ;
        RECT 4.400 149.240 295.600 149.960 ;
        RECT 4.400 148.560 296.000 149.240 ;
        RECT 4.000 147.920 296.000 148.560 ;
        RECT 4.000 146.560 295.600 147.920 ;
        RECT 4.400 146.520 295.600 146.560 ;
        RECT 4.400 145.200 296.000 146.520 ;
        RECT 4.400 145.160 295.600 145.200 ;
        RECT 4.000 143.800 295.600 145.160 ;
        RECT 4.000 143.160 296.000 143.800 ;
        RECT 4.400 142.480 296.000 143.160 ;
        RECT 4.400 141.760 295.600 142.480 ;
        RECT 4.000 141.080 295.600 141.760 ;
        RECT 4.000 139.760 296.000 141.080 ;
        RECT 4.400 138.360 295.600 139.760 ;
        RECT 4.000 137.040 296.000 138.360 ;
        RECT 4.000 136.360 295.600 137.040 ;
        RECT 4.400 135.640 295.600 136.360 ;
        RECT 4.400 134.960 296.000 135.640 ;
        RECT 4.000 134.320 296.000 134.960 ;
        RECT 4.000 132.960 295.600 134.320 ;
        RECT 4.400 132.920 295.600 132.960 ;
        RECT 4.400 131.600 296.000 132.920 ;
        RECT 4.400 131.560 295.600 131.600 ;
        RECT 4.000 130.200 295.600 131.560 ;
        RECT 4.000 129.560 296.000 130.200 ;
        RECT 4.400 128.880 296.000 129.560 ;
        RECT 4.400 128.160 295.600 128.880 ;
        RECT 4.000 127.480 295.600 128.160 ;
        RECT 4.000 126.160 296.000 127.480 ;
        RECT 4.400 124.760 295.600 126.160 ;
        RECT 4.000 123.440 296.000 124.760 ;
        RECT 4.000 122.760 295.600 123.440 ;
        RECT 4.400 122.040 295.600 122.760 ;
        RECT 4.400 121.360 296.000 122.040 ;
        RECT 4.000 120.720 296.000 121.360 ;
        RECT 4.000 119.360 295.600 120.720 ;
        RECT 4.400 119.320 295.600 119.360 ;
        RECT 4.400 118.000 296.000 119.320 ;
        RECT 4.400 117.960 295.600 118.000 ;
        RECT 4.000 116.600 295.600 117.960 ;
        RECT 4.000 115.960 296.000 116.600 ;
        RECT 4.400 115.280 296.000 115.960 ;
        RECT 4.400 114.560 295.600 115.280 ;
        RECT 4.000 113.880 295.600 114.560 ;
        RECT 4.000 112.560 296.000 113.880 ;
        RECT 4.400 111.160 295.600 112.560 ;
        RECT 4.000 109.840 296.000 111.160 ;
        RECT 4.000 109.160 295.600 109.840 ;
        RECT 4.400 108.440 295.600 109.160 ;
        RECT 4.400 107.760 296.000 108.440 ;
        RECT 4.000 107.120 296.000 107.760 ;
        RECT 4.000 105.760 295.600 107.120 ;
        RECT 4.400 105.720 295.600 105.760 ;
        RECT 4.400 104.400 296.000 105.720 ;
        RECT 4.400 104.360 295.600 104.400 ;
        RECT 4.000 103.000 295.600 104.360 ;
        RECT 4.000 102.360 296.000 103.000 ;
        RECT 4.400 101.680 296.000 102.360 ;
        RECT 4.400 100.960 295.600 101.680 ;
        RECT 4.000 100.280 295.600 100.960 ;
        RECT 4.000 98.960 296.000 100.280 ;
        RECT 4.400 97.560 295.600 98.960 ;
        RECT 4.000 96.240 296.000 97.560 ;
        RECT 4.000 95.560 295.600 96.240 ;
        RECT 4.400 94.840 295.600 95.560 ;
        RECT 4.400 94.160 296.000 94.840 ;
        RECT 4.000 93.520 296.000 94.160 ;
        RECT 4.000 92.160 295.600 93.520 ;
        RECT 4.400 92.120 295.600 92.160 ;
        RECT 4.400 90.800 296.000 92.120 ;
        RECT 4.400 90.760 295.600 90.800 ;
        RECT 4.000 89.400 295.600 90.760 ;
        RECT 4.000 88.760 296.000 89.400 ;
        RECT 4.400 88.080 296.000 88.760 ;
        RECT 4.400 87.360 295.600 88.080 ;
        RECT 4.000 86.680 295.600 87.360 ;
        RECT 4.000 85.360 296.000 86.680 ;
        RECT 4.400 83.960 295.600 85.360 ;
        RECT 4.000 82.640 296.000 83.960 ;
        RECT 4.000 81.960 295.600 82.640 ;
        RECT 4.400 81.240 295.600 81.960 ;
        RECT 4.400 80.560 296.000 81.240 ;
        RECT 4.000 79.920 296.000 80.560 ;
        RECT 4.000 78.560 295.600 79.920 ;
        RECT 4.400 78.520 295.600 78.560 ;
        RECT 4.400 77.200 296.000 78.520 ;
        RECT 4.400 77.160 295.600 77.200 ;
        RECT 4.000 75.800 295.600 77.160 ;
        RECT 4.000 75.160 296.000 75.800 ;
        RECT 4.400 74.480 296.000 75.160 ;
        RECT 4.400 73.760 295.600 74.480 ;
        RECT 4.000 73.080 295.600 73.760 ;
        RECT 4.000 71.760 296.000 73.080 ;
        RECT 4.400 70.360 295.600 71.760 ;
        RECT 4.000 69.040 296.000 70.360 ;
        RECT 4.000 68.360 295.600 69.040 ;
        RECT 4.400 67.640 295.600 68.360 ;
        RECT 4.400 66.960 296.000 67.640 ;
        RECT 4.000 66.320 296.000 66.960 ;
        RECT 4.000 64.960 295.600 66.320 ;
        RECT 4.400 64.920 295.600 64.960 ;
        RECT 4.400 63.600 296.000 64.920 ;
        RECT 4.400 63.560 295.600 63.600 ;
        RECT 4.000 62.200 295.600 63.560 ;
        RECT 4.000 61.560 296.000 62.200 ;
        RECT 4.400 60.880 296.000 61.560 ;
        RECT 4.400 60.160 295.600 60.880 ;
        RECT 4.000 59.480 295.600 60.160 ;
        RECT 4.000 58.160 296.000 59.480 ;
        RECT 4.400 56.760 295.600 58.160 ;
        RECT 4.000 55.440 296.000 56.760 ;
        RECT 4.000 54.760 295.600 55.440 ;
        RECT 4.400 54.040 295.600 54.760 ;
        RECT 4.400 53.360 296.000 54.040 ;
        RECT 4.000 52.720 296.000 53.360 ;
        RECT 4.000 51.360 295.600 52.720 ;
        RECT 4.400 51.320 295.600 51.360 ;
        RECT 4.400 50.000 296.000 51.320 ;
        RECT 4.400 49.960 295.600 50.000 ;
        RECT 4.000 48.600 295.600 49.960 ;
        RECT 4.000 47.960 296.000 48.600 ;
        RECT 4.400 47.280 296.000 47.960 ;
        RECT 4.400 46.560 295.600 47.280 ;
        RECT 4.000 45.880 295.600 46.560 ;
        RECT 4.000 44.560 296.000 45.880 ;
        RECT 4.400 43.160 295.600 44.560 ;
        RECT 4.000 41.840 296.000 43.160 ;
        RECT 4.000 41.160 295.600 41.840 ;
        RECT 4.400 40.440 295.600 41.160 ;
        RECT 4.400 39.760 296.000 40.440 ;
        RECT 4.000 39.120 296.000 39.760 ;
        RECT 4.000 37.760 295.600 39.120 ;
        RECT 4.400 37.720 295.600 37.760 ;
        RECT 4.400 36.400 296.000 37.720 ;
        RECT 4.400 36.360 295.600 36.400 ;
        RECT 4.000 35.000 295.600 36.360 ;
        RECT 4.000 34.360 296.000 35.000 ;
        RECT 4.400 33.680 296.000 34.360 ;
        RECT 4.400 32.960 295.600 33.680 ;
        RECT 4.000 32.280 295.600 32.960 ;
        RECT 4.000 30.960 296.000 32.280 ;
        RECT 4.400 29.560 295.600 30.960 ;
        RECT 4.000 28.240 296.000 29.560 ;
        RECT 4.000 27.560 295.600 28.240 ;
        RECT 4.400 26.840 295.600 27.560 ;
        RECT 4.400 26.160 296.000 26.840 ;
        RECT 4.000 25.520 296.000 26.160 ;
        RECT 4.000 24.160 295.600 25.520 ;
        RECT 4.400 24.120 295.600 24.160 ;
        RECT 4.400 22.800 296.000 24.120 ;
        RECT 4.400 22.760 295.600 22.800 ;
        RECT 4.000 21.400 295.600 22.760 ;
        RECT 4.000 20.760 296.000 21.400 ;
        RECT 4.400 20.080 296.000 20.760 ;
        RECT 4.400 19.360 295.600 20.080 ;
        RECT 4.000 18.680 295.600 19.360 ;
        RECT 4.000 17.360 296.000 18.680 ;
        RECT 4.400 15.960 295.600 17.360 ;
        RECT 4.000 14.640 296.000 15.960 ;
        RECT 4.000 13.960 295.600 14.640 ;
        RECT 4.400 13.240 295.600 13.960 ;
        RECT 4.400 12.560 296.000 13.240 ;
        RECT 4.000 11.920 296.000 12.560 ;
        RECT 4.000 10.560 295.600 11.920 ;
        RECT 4.400 10.520 295.600 10.560 ;
        RECT 4.400 9.200 296.000 10.520 ;
        RECT 4.400 9.160 295.600 9.200 ;
        RECT 4.000 7.800 295.600 9.160 ;
        RECT 4.000 6.480 296.000 7.800 ;
        RECT 4.000 5.615 295.600 6.480 ;
      LAYER met4 ;
        RECT 79.415 11.735 97.440 303.785 ;
        RECT 99.840 11.735 174.240 303.785 ;
        RECT 176.640 11.735 219.585 303.785 ;
  END
END multiplexer
END LIBRARY

