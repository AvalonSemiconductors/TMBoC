// This is the unpowered netlist.
module tune_player (OP,
    clk,
    rst);
 output OP;
 input clk;
 input rst;

 wire \LFSR[0] ;
 wire \LFSR[1] ;
 wire \LFSR[2] ;
 wire \LFSR[3] ;
 wire \LFSR[4] ;
 wire \LFSR[5] ;
 wire \LFSR[6] ;
 wire OP_reg;
 wire \PC[0] ;
 wire \PC[1] ;
 wire \PC[2] ;
 wire \PC[3] ;
 wire \PC[4] ;
 wire \PC[5] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire \clock_div[0] ;
 wire \clock_div[1] ;
 wire \clock_div[2] ;
 wire \clock_div[3] ;
 wire \clock_div[4] ;
 wire \clock_div[5] ;
 wire \clock_div[6] ;
 wire \clock_div[7] ;
 wire \clock_div[8] ;
 wire just_inc;
 wire just_rst;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire prev_clk_div;
 wire \rhythm_LFSR[0] ;
 wire \rhythm_LFSR[1] ;
 wire \rhythm_LFSR[2] ;
 wire \rhythm_LFSR[3] ;
 wire \tempo_LFSR[0] ;
 wire \tempo_LFSR[1] ;
 wire \tempo_LFSR[2] ;
 wire \tempo_LFSR[3] ;
 wire \tune_ROM[0] ;
 wire \tune_ROM[1] ;
 wire \tune_ROM[2] ;
 wire \tune_ROM[3] ;
 wire \tune_ROM[4] ;
 wire \tune_ROM[5] ;

 sky130_fd_sc_hd__decap_3 FILLER_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__inv_2 _199_ (.A(\tempo_LFSR[2] ),
    .Y(_181_));
 sky130_fd_sc_hd__inv_2 _200_ (.A(\PC[2] ),
    .Y(_182_));
 sky130_fd_sc_hd__inv_2 _201_ (.A(\PC[1] ),
    .Y(_183_));
 sky130_fd_sc_hd__clkinv_4 _202_ (.A(just_rst),
    .Y(_184_));
 sky130_fd_sc_hd__inv_2 _203_ (.A(\clock_div[7] ),
    .Y(_185_));
 sky130_fd_sc_hd__inv_2 _204_ (.A(prev_clk_div),
    .Y(_186_));
 sky130_fd_sc_hd__clkinv_4 _205_ (.A(net8),
    .Y(_187_));
 sky130_fd_sc_hd__inv_2 _206_ (.A(\tune_ROM[4] ),
    .Y(_188_));
 sky130_fd_sc_hd__and3_1 _207_ (.A(\clock_div[0] ),
    .B(\clock_div[2] ),
    .C(\clock_div[1] ),
    .X(_189_));
 sky130_fd_sc_hd__and4_4 _208_ (.A(\clock_div[0] ),
    .B(\clock_div[2] ),
    .C(\clock_div[3] ),
    .D(\clock_div[1] ),
    .X(_190_));
 sky130_fd_sc_hd__and2_2 _209_ (.A(\clock_div[4] ),
    .B(\clock_div[5] ),
    .X(_191_));
 sky130_fd_sc_hd__and2_1 _210_ (.A(_190_),
    .B(_191_),
    .X(_192_));
 sky130_fd_sc_hd__and3_1 _211_ (.A(\clock_div[6] ),
    .B(_190_),
    .C(_191_),
    .X(_193_));
 sky130_fd_sc_hd__a41o_1 _212_ (.A1(\clock_div[6] ),
    .A2(\clock_div[7] ),
    .A3(_190_),
    .A4(_191_),
    .B1(\clock_div[8] ),
    .X(_194_));
 sky130_fd_sc_hd__nand4_2 _213_ (.A(\clock_div[6] ),
    .B(\clock_div[8] ),
    .C(_190_),
    .D(_191_),
    .Y(_195_));
 sky130_fd_sc_hd__o211a_4 _214_ (.A1(_185_),
    .A2(_195_),
    .B1(_194_),
    .C1(_186_),
    .X(_196_));
 sky130_fd_sc_hd__nor2_2 _215_ (.A(just_rst),
    .B(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__or2_1 _216_ (.A(\rhythm_LFSR[1] ),
    .B(\rhythm_LFSR[0] ),
    .X(_198_));
 sky130_fd_sc_hd__or3b_2 _217_ (.A(_198_),
    .B(\rhythm_LFSR[2] ),
    .C_N(\rhythm_LFSR[3] ),
    .X(_039_));
 sky130_fd_sc_hd__inv_2 _218_ (.A(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__nor2_1 _219_ (.A(just_rst),
    .B(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__nand2_2 _220_ (.A(_184_),
    .B(_039_),
    .Y(_042_));
 sky130_fd_sc_hd__or4b_4 _221_ (.A(\tempo_LFSR[2] ),
    .B(\tempo_LFSR[1] ),
    .C(\tempo_LFSR[0] ),
    .D_N(\tempo_LFSR[3] ),
    .X(_043_));
 sky130_fd_sc_hd__inv_2 _222_ (.A(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__nand2_1 _223_ (.A(_184_),
    .B(_043_),
    .Y(_045_));
 sky130_fd_sc_hd__a31o_1 _224_ (.A1(_196_),
    .A2(_040_),
    .A3(_044_),
    .B1(just_rst),
    .X(_046_));
 sky130_fd_sc_hd__o2111a_4 _225_ (.A1(just_rst),
    .A2(_196_),
    .B1(_042_),
    .C1(_045_),
    .D1(\PC[0] ),
    .X(_047_));
 sky130_fd_sc_hd__xnor2_2 _226_ (.A(\PC[1] ),
    .B(_047_),
    .Y(_048_));
 sky130_fd_sc_hd__or2_4 _227_ (.A(net8),
    .B(_048_),
    .X(_049_));
 sky130_fd_sc_hd__inv_2 _228_ (.A(_049_),
    .Y(_011_));
 sky130_fd_sc_hd__nor2_1 _229_ (.A(\PC[2] ),
    .B(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__or3_2 _230_ (.A(\PC[2] ),
    .B(net8),
    .C(_048_),
    .X(_051_));
 sky130_fd_sc_hd__a311o_1 _231_ (.A1(_196_),
    .A2(_040_),
    .A3(_044_),
    .B1(just_rst),
    .C1(\PC[0] ),
    .X(_052_));
 sky130_fd_sc_hd__and2b_1 _232_ (.A_N(_047_),
    .B(_052_),
    .X(_053_));
 sky130_fd_sc_hd__nor3b_4 _233_ (.A(net8),
    .B(_047_),
    .C_N(_052_),
    .Y(_010_));
 sky130_fd_sc_hd__and2_2 _234_ (.A(_183_),
    .B(_010_),
    .X(_054_));
 sky130_fd_sc_hd__nor2_1 _235_ (.A(_050_),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__and3_1 _236_ (.A(\PC[2] ),
    .B(\PC[1] ),
    .C(_047_),
    .X(_056_));
 sky130_fd_sc_hd__and4_2 _237_ (.A(\PC[3] ),
    .B(\PC[2] ),
    .C(\PC[1] ),
    .D(_047_),
    .X(_057_));
 sky130_fd_sc_hd__xnor2_1 _238_ (.A(\PC[4] ),
    .B(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__or2_4 _239_ (.A(net9),
    .B(_058_),
    .X(_059_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(_059_),
    .Y(_014_));
 sky130_fd_sc_hd__and2_2 _241_ (.A(\PC[1] ),
    .B(_010_),
    .X(_060_));
 sky130_fd_sc_hd__nand2_2 _242_ (.A(\PC[1] ),
    .B(_010_),
    .Y(_061_));
 sky130_fd_sc_hd__a21oi_2 _243_ (.A1(\PC[1] ),
    .A2(_047_),
    .B1(\PC[2] ),
    .Y(_062_));
 sky130_fd_sc_hd__or2_4 _244_ (.A(_056_),
    .B(_062_),
    .X(_063_));
 sky130_fd_sc_hd__a31o_1 _245_ (.A1(\PC[2] ),
    .A2(\PC[1] ),
    .A3(_047_),
    .B1(\PC[3] ),
    .X(_064_));
 sky130_fd_sc_hd__nand2b_1 _246_ (.A_N(_057_),
    .B(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__or3b_4 _247_ (.A(net9),
    .B(_057_),
    .C_N(_064_),
    .X(_066_));
 sky130_fd_sc_hd__inv_2 _248_ (.A(_066_),
    .Y(_013_));
 sky130_fd_sc_hd__nand2_1 _249_ (.A(_063_),
    .B(net4),
    .Y(_067_));
 sky130_fd_sc_hd__and3_1 _250_ (.A(_061_),
    .B(_063_),
    .C(net4),
    .X(_068_));
 sky130_fd_sc_hd__a21oi_1 _251_ (.A1(\PC[4] ),
    .A2(_057_),
    .B1(\PC[5] ),
    .Y(_069_));
 sky130_fd_sc_hd__a31o_1 _252_ (.A1(\PC[5] ),
    .A2(\PC[4] ),
    .A3(_057_),
    .B1(net9),
    .X(_070_));
 sky130_fd_sc_hd__or2_4 _253_ (.A(_069_),
    .B(_070_),
    .X(_071_));
 sky130_fd_sc_hd__clkinv_4 _254_ (.A(_071_),
    .Y(_015_));
 sky130_fd_sc_hd__or3_4 _255_ (.A(net8),
    .B(_056_),
    .C(_062_),
    .X(_072_));
 sky130_fd_sc_hd__inv_2 _256_ (.A(_072_),
    .Y(_012_));
 sky130_fd_sc_hd__o21ai_1 _257_ (.A1(_060_),
    .A2(_072_),
    .B1(_051_),
    .Y(_073_));
 sky130_fd_sc_hd__a221o_1 _258_ (.A1(\PC[2] ),
    .A2(_054_),
    .B1(net4),
    .B2(_073_),
    .C1(_059_),
    .X(_074_));
 sky130_fd_sc_hd__o311a_1 _259_ (.A1(_055_),
    .A2(net3),
    .A3(_068_),
    .B1(_015_),
    .C1(_074_),
    .X(_075_));
 sky130_fd_sc_hd__or3_2 _260_ (.A(net8),
    .B(_048_),
    .C(_053_),
    .X(_076_));
 sky130_fd_sc_hd__or4_4 _261_ (.A(net8),
    .B(_053_),
    .C(_056_),
    .D(_062_),
    .X(_077_));
 sky130_fd_sc_hd__or2_4 _262_ (.A(_049_),
    .B(_077_),
    .X(_078_));
 sky130_fd_sc_hd__nand2_1 _263_ (.A(_060_),
    .B(_063_),
    .Y(_079_));
 sky130_fd_sc_hd__a21o_1 _264_ (.A1(_060_),
    .A2(_063_),
    .B1(_066_),
    .X(_080_));
 sky130_fd_sc_hd__and3b_1 _265_ (.A_N(_080_),
    .B(_049_),
    .C(_012_),
    .X(_081_));
 sky130_fd_sc_hd__a21oi_1 _266_ (.A1(_078_),
    .A2(_079_),
    .B1(net4),
    .Y(_082_));
 sky130_fd_sc_hd__or3_1 _267_ (.A(net3),
    .B(_081_),
    .C(_082_),
    .X(_083_));
 sky130_fd_sc_hd__nor2_1 _268_ (.A(_063_),
    .B(net4),
    .Y(_084_));
 sky130_fd_sc_hd__o31ai_1 _269_ (.A1(_011_),
    .A2(_010_),
    .A3(_084_),
    .B1(_014_),
    .Y(_085_));
 sky130_fd_sc_hd__a31o_1 _270_ (.A1(_071_),
    .A2(_083_),
    .A3(_085_),
    .B1(_075_),
    .X(_000_));
 sky130_fd_sc_hd__nor3_1 _271_ (.A(\PC[4] ),
    .B(_066_),
    .C(_079_),
    .Y(_086_));
 sky130_fd_sc_hd__o2111a_1 _272_ (.A1(\PC[2] ),
    .A2(net5),
    .B1(_183_),
    .C1(\PC[4] ),
    .D1(_010_),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _273_ (.A0(_060_),
    .A1(_054_),
    .S(_067_),
    .X(_088_));
 sky130_fd_sc_hd__nor2_2 _274_ (.A(_011_),
    .B(_077_),
    .Y(_089_));
 sky130_fd_sc_hd__nor2_1 _275_ (.A(net4),
    .B(_089_),
    .Y(_090_));
 sky130_fd_sc_hd__nor2_1 _276_ (.A(_182_),
    .B(_061_),
    .Y(_091_));
 sky130_fd_sc_hd__o221a_1 _277_ (.A1(net4),
    .A2(_089_),
    .B1(_091_),
    .B2(_065_),
    .C1(net3),
    .X(_092_));
 sky130_fd_sc_hd__a211o_1 _278_ (.A1(_059_),
    .A2(_088_),
    .B1(_092_),
    .C1(_071_),
    .X(_093_));
 sky130_fd_sc_hd__o31a_1 _279_ (.A1(_015_),
    .A2(_086_),
    .A3(_087_),
    .B1(_093_),
    .X(_001_));
 sky130_fd_sc_hd__nand2_1 _280_ (.A(_072_),
    .B(_076_),
    .Y(_094_));
 sky130_fd_sc_hd__nand2_1 _281_ (.A(\PC[2] ),
    .B(_011_),
    .Y(_095_));
 sky130_fd_sc_hd__o2bb2a_1 _282_ (.A1_N(_072_),
    .A2_N(_076_),
    .B1(_182_),
    .B2(_049_),
    .X(_096_));
 sky130_fd_sc_hd__a21oi_1 _283_ (.A1(_051_),
    .A2(_077_),
    .B1(_066_),
    .Y(_097_));
 sky130_fd_sc_hd__a21oi_1 _284_ (.A1(_066_),
    .A2(_096_),
    .B1(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__a2111o_1 _285_ (.A1(_049_),
    .A2(_072_),
    .B1(_015_),
    .C1(_066_),
    .D1(_060_),
    .X(_099_));
 sky130_fd_sc_hd__o211a_1 _286_ (.A1(_071_),
    .A2(_098_),
    .B1(_099_),
    .C1(_059_),
    .X(_100_));
 sky130_fd_sc_hd__a21oi_1 _287_ (.A1(_010_),
    .A2(_095_),
    .B1(_068_),
    .Y(_101_));
 sky130_fd_sc_hd__and3_1 _288_ (.A(_054_),
    .B(_063_),
    .C(net4),
    .X(_102_));
 sky130_fd_sc_hd__a211o_1 _289_ (.A1(_078_),
    .A2(_101_),
    .B1(_102_),
    .C1(_071_),
    .X(_103_));
 sky130_fd_sc_hd__nand2_1 _290_ (.A(_078_),
    .B(_094_),
    .Y(_104_));
 sky130_fd_sc_hd__a221o_1 _291_ (.A1(_061_),
    .A2(_090_),
    .B1(_104_),
    .B2(net4),
    .C1(_015_),
    .X(_105_));
 sky130_fd_sc_hd__a31o_1 _292_ (.A1(net3),
    .A2(_103_),
    .A3(_105_),
    .B1(_100_),
    .X(_002_));
 sky130_fd_sc_hd__and2b_1 _293_ (.A_N(_054_),
    .B(_072_),
    .X(_106_));
 sky130_fd_sc_hd__o21ai_1 _294_ (.A1(_066_),
    .A2(_096_),
    .B1(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__o31a_1 _295_ (.A1(_066_),
    .A2(_096_),
    .A3(_106_),
    .B1(_015_),
    .X(_108_));
 sky130_fd_sc_hd__o211a_1 _296_ (.A1(_011_),
    .A2(_010_),
    .B1(_066_),
    .C1(_077_),
    .X(_109_));
 sky130_fd_sc_hd__a31o_1 _297_ (.A1(_051_),
    .A2(net5),
    .A3(_078_),
    .B1(_015_),
    .X(_110_));
 sky130_fd_sc_hd__a2bb2o_1 _298_ (.A1_N(_110_),
    .A2_N(_109_),
    .B1(_108_),
    .B2(_107_),
    .X(_111_));
 sky130_fd_sc_hd__or3b_1 _299_ (.A(_102_),
    .B(_071_),
    .C_N(_076_),
    .X(_112_));
 sky130_fd_sc_hd__nor2_1 _300_ (.A(net4),
    .B(_106_),
    .Y(_113_));
 sky130_fd_sc_hd__o41a_1 _301_ (.A1(_050_),
    .A2(_015_),
    .A3(_091_),
    .A4(_113_),
    .B1(_059_),
    .X(_114_));
 sky130_fd_sc_hd__a22o_1 _302_ (.A1(_014_),
    .A2(_111_),
    .B1(_112_),
    .B2(_114_),
    .X(_003_));
 sky130_fd_sc_hd__o22a_1 _303_ (.A1(_011_),
    .A2(_010_),
    .B1(_060_),
    .B2(_072_),
    .X(_115_));
 sky130_fd_sc_hd__a211o_1 _304_ (.A1(net3),
    .A2(_067_),
    .B1(_113_),
    .C1(_115_),
    .X(_116_));
 sky130_fd_sc_hd__a21oi_1 _305_ (.A1(net3),
    .A2(_115_),
    .B1(_015_),
    .Y(_117_));
 sky130_fd_sc_hd__mux2_1 _306_ (.A0(\PC[3] ),
    .A1(_080_),
    .S(_078_),
    .X(_118_));
 sky130_fd_sc_hd__o21ai_1 _307_ (.A1(_061_),
    .A2(_067_),
    .B1(net3),
    .Y(_119_));
 sky130_fd_sc_hd__o22a_1 _308_ (.A1(net3),
    .A2(_118_),
    .B1(_119_),
    .B2(_089_),
    .X(_120_));
 sky130_fd_sc_hd__a2bb2o_1 _309_ (.A1_N(_071_),
    .A2_N(_120_),
    .B1(_117_),
    .B2(_116_),
    .X(_004_));
 sky130_fd_sc_hd__a2bb2o_1 _310_ (.A1_N(\PC[4] ),
    .A2_N(_115_),
    .B1(net3),
    .B2(_048_),
    .X(_121_));
 sky130_fd_sc_hd__nand2_1 _311_ (.A(net5),
    .B(_121_),
    .Y(_122_));
 sky130_fd_sc_hd__o211a_1 _312_ (.A1(\PC[3] ),
    .A2(_078_),
    .B1(_080_),
    .C1(_058_),
    .X(_123_));
 sky130_fd_sc_hd__o2bb2a_1 _313_ (.A1_N(_117_),
    .A2_N(_122_),
    .B1(_123_),
    .B2(_071_),
    .X(_005_));
 sky130_fd_sc_hd__and2_1 _314_ (.A(OP_reg),
    .B(just_inc),
    .X(net2));
 sky130_fd_sc_hd__nor2_4 _315_ (.A(net8),
    .B(_197_),
    .Y(_124_));
 sky130_fd_sc_hd__nand2_1 _316_ (.A(\tune_ROM[1] ),
    .B(_042_),
    .Y(_125_));
 sky130_fd_sc_hd__o21a_1 _317_ (.A1(\rhythm_LFSR[1] ),
    .A2(_042_),
    .B1(_125_),
    .X(_126_));
 sky130_fd_sc_hd__mux2_1 _318_ (.A0(\rhythm_LFSR[0] ),
    .A1(_126_),
    .S(_124_),
    .X(_006_));
 sky130_fd_sc_hd__nand2_1 _319_ (.A(\tune_ROM[0] ),
    .B(\tune_ROM[1] ),
    .Y(_127_));
 sky130_fd_sc_hd__or2_1 _320_ (.A(\tune_ROM[0] ),
    .B(\tune_ROM[1] ),
    .X(_128_));
 sky130_fd_sc_hd__a32o_1 _321_ (.A1(_042_),
    .A2(_127_),
    .A3(_128_),
    .B1(\rhythm_LFSR[2] ),
    .B2(_184_),
    .X(_129_));
 sky130_fd_sc_hd__mux2_1 _322_ (.A0(\rhythm_LFSR[1] ),
    .A1(_129_),
    .S(_124_),
    .X(_007_));
 sky130_fd_sc_hd__and2_2 _323_ (.A(_042_),
    .B(_124_),
    .X(_130_));
 sky130_fd_sc_hd__o22a_1 _324_ (.A1(just_rst),
    .A2(\rhythm_LFSR[3] ),
    .B1(\tune_ROM[0] ),
    .B2(_041_),
    .X(_131_));
 sky130_fd_sc_hd__mux2_1 _325_ (.A0(\rhythm_LFSR[2] ),
    .A1(_131_),
    .S(_124_),
    .X(_008_));
 sky130_fd_sc_hd__a21oi_1 _326_ (.A1(\rhythm_LFSR[1] ),
    .A2(\rhythm_LFSR[0] ),
    .B1(just_rst),
    .Y(_132_));
 sky130_fd_sc_hd__a2bb2o_1 _327_ (.A1_N(\tune_ROM[0] ),
    .A2_N(_125_),
    .B1(_132_),
    .B2(_198_),
    .X(_133_));
 sky130_fd_sc_hd__mux2_1 _328_ (.A0(\rhythm_LFSR[3] ),
    .A1(_133_),
    .S(_124_),
    .X(_009_));
 sky130_fd_sc_hd__o21ba_1 _329_ (.A1(_197_),
    .A2(_041_),
    .B1_N(just_inc),
    .X(_134_));
 sky130_fd_sc_hd__nor3_1 _330_ (.A(net8),
    .B(_046_),
    .C(_134_),
    .Y(_016_));
 sky130_fd_sc_hd__or2_1 _331_ (.A(\LFSR[1] ),
    .B(\LFSR[0] ),
    .X(_135_));
 sky130_fd_sc_hd__or4b_2 _332_ (.A(\LFSR[3] ),
    .B(_135_),
    .C(\LFSR[2] ),
    .D_N(\LFSR[6] ),
    .X(_136_));
 sky130_fd_sc_hd__o31ai_4 _333_ (.A1(\LFSR[5] ),
    .A2(\LFSR[4] ),
    .A3(_136_),
    .B1(_184_),
    .Y(_137_));
 sky130_fd_sc_hd__o21ai_1 _334_ (.A1(OP_reg),
    .A2(_137_),
    .B1(_187_),
    .Y(_138_));
 sky130_fd_sc_hd__a21oi_1 _335_ (.A1(OP_reg),
    .A2(_137_),
    .B1(_138_),
    .Y(_017_));
 sky130_fd_sc_hd__nor2_1 _336_ (.A(\tune_ROM[2] ),
    .B(\tune_ROM[3] ),
    .Y(_139_));
 sky130_fd_sc_hd__o21ai_1 _337_ (.A1(net6),
    .A2(_139_),
    .B1(\tune_ROM[4] ),
    .Y(_140_));
 sky130_fd_sc_hd__nand2_2 _338_ (.A(\tune_ROM[2] ),
    .B(\tune_ROM[3] ),
    .Y(_141_));
 sky130_fd_sc_hd__or2_2 _339_ (.A(\tune_ROM[4] ),
    .B(\tune_ROM[3] ),
    .X(_142_));
 sky130_fd_sc_hd__nand3_1 _340_ (.A(_140_),
    .B(_141_),
    .C(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__mux2_1 _341_ (.A0(\LFSR[1] ),
    .A1(_143_),
    .S(_137_),
    .X(_144_));
 sky130_fd_sc_hd__mux2_1 _342_ (.A0(\LFSR[0] ),
    .A1(_144_),
    .S(_187_),
    .X(_018_));
 sky130_fd_sc_hd__nor2_1 _343_ (.A(\tune_ROM[4] ),
    .B(_139_),
    .Y(_145_));
 sky130_fd_sc_hd__and2_1 _344_ (.A(\tune_ROM[4] ),
    .B(_139_),
    .X(_146_));
 sky130_fd_sc_hd__o21ai_1 _345_ (.A1(_145_),
    .A2(_146_),
    .B1(net6),
    .Y(_147_));
 sky130_fd_sc_hd__or2_1 _346_ (.A(net6),
    .B(_141_),
    .X(_148_));
 sky130_fd_sc_hd__a32o_1 _347_ (.A1(_137_),
    .A2(_147_),
    .A3(_148_),
    .B1(\LFSR[2] ),
    .B2(_184_),
    .X(_149_));
 sky130_fd_sc_hd__mux2_1 _348_ (.A0(\LFSR[1] ),
    .A1(_149_),
    .S(_187_),
    .X(_019_));
 sky130_fd_sc_hd__nand2_1 _349_ (.A(\tune_ROM[4] ),
    .B(\tune_ROM[3] ),
    .Y(_150_));
 sky130_fd_sc_hd__o21ai_1 _350_ (.A1(_188_),
    .A2(\tune_ROM[5] ),
    .B1(\tune_ROM[2] ),
    .Y(_151_));
 sky130_fd_sc_hd__o211ai_1 _351_ (.A1(net6),
    .A2(_142_),
    .B1(_150_),
    .C1(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__mux2_1 _352_ (.A0(\LFSR[3] ),
    .A1(_152_),
    .S(_137_),
    .X(_153_));
 sky130_fd_sc_hd__mux2_1 _353_ (.A0(\LFSR[2] ),
    .A1(_153_),
    .S(_187_),
    .X(_020_));
 sky130_fd_sc_hd__or2_1 _354_ (.A(\tune_ROM[4] ),
    .B(_141_),
    .X(_154_));
 sky130_fd_sc_hd__nand2_1 _355_ (.A(\tune_ROM[4] ),
    .B(_141_),
    .Y(_155_));
 sky130_fd_sc_hd__a22o_1 _356_ (.A1(net6),
    .A2(_141_),
    .B1(_154_),
    .B2(_155_),
    .X(_156_));
 sky130_fd_sc_hd__mux2_1 _357_ (.A0(\LFSR[4] ),
    .A1(_156_),
    .S(_137_),
    .X(_157_));
 sky130_fd_sc_hd__mux2_1 _358_ (.A0(\LFSR[3] ),
    .A1(_157_),
    .S(_187_),
    .X(_021_));
 sky130_fd_sc_hd__a21bo_1 _359_ (.A1(_188_),
    .A2(\tune_ROM[2] ),
    .B1_N(net6),
    .X(_158_));
 sky130_fd_sc_hd__a211o_1 _360_ (.A1(_142_),
    .A2(_155_),
    .B1(_146_),
    .C1(net6),
    .X(_159_));
 sky130_fd_sc_hd__o21ai_1 _361_ (.A1(_146_),
    .A2(_158_),
    .B1(_159_),
    .Y(_160_));
 sky130_fd_sc_hd__mux2_1 _362_ (.A0(\LFSR[5] ),
    .A1(_160_),
    .S(_137_),
    .X(_161_));
 sky130_fd_sc_hd__mux2_1 _363_ (.A0(\LFSR[4] ),
    .A1(_161_),
    .S(_187_),
    .X(_022_));
 sky130_fd_sc_hd__and4bb_1 _364_ (.A_N(net6),
    .B_N(_139_),
    .C(_142_),
    .D(_150_),
    .X(_162_));
 sky130_fd_sc_hd__a31o_1 _365_ (.A1(net6),
    .A2(_141_),
    .A3(_145_),
    .B1(_162_),
    .X(_163_));
 sky130_fd_sc_hd__nand2_1 _366_ (.A(_137_),
    .B(_163_),
    .Y(_164_));
 sky130_fd_sc_hd__o21a_1 _367_ (.A1(just_rst),
    .A2(\LFSR[6] ),
    .B1(_187_),
    .X(_165_));
 sky130_fd_sc_hd__a22o_1 _368_ (.A1(net7),
    .A2(\LFSR[5] ),
    .B1(_164_),
    .B2(_165_),
    .X(_023_));
 sky130_fd_sc_hd__nand3b_1 _369_ (.A_N(net6),
    .B(_154_),
    .C(_155_),
    .Y(_166_));
 sky130_fd_sc_hd__nand2_1 _370_ (.A(\LFSR[1] ),
    .B(\LFSR[0] ),
    .Y(_167_));
 sky130_fd_sc_hd__a21oi_1 _371_ (.A1(_135_),
    .A2(_167_),
    .B1(_137_),
    .Y(_168_));
 sky130_fd_sc_hd__a311o_1 _372_ (.A1(_137_),
    .A2(_158_),
    .A3(_166_),
    .B1(_168_),
    .C1(net7),
    .X(_169_));
 sky130_fd_sc_hd__a21bo_1 _373_ (.A1(net7),
    .A2(\LFSR[6] ),
    .B1_N(_169_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _374_ (.A0(\clock_div[8] ),
    .A1(prev_clk_div),
    .S(net9),
    .X(_025_));
 sky130_fd_sc_hd__nor2_1 _375_ (.A(\clock_div[0] ),
    .B(net7),
    .Y(_026_));
 sky130_fd_sc_hd__a21oi_1 _376_ (.A1(\clock_div[0] ),
    .A2(\clock_div[1] ),
    .B1(net7),
    .Y(_170_));
 sky130_fd_sc_hd__o21a_1 _377_ (.A1(\clock_div[0] ),
    .A2(\clock_div[1] ),
    .B1(_170_),
    .X(_027_));
 sky130_fd_sc_hd__a21oi_1 _378_ (.A1(\clock_div[0] ),
    .A2(\clock_div[1] ),
    .B1(\clock_div[2] ),
    .Y(_171_));
 sky130_fd_sc_hd__nor3_1 _379_ (.A(net7),
    .B(_189_),
    .C(_171_),
    .Y(_028_));
 sky130_fd_sc_hd__nor2_1 _380_ (.A(net7),
    .B(_190_),
    .Y(_172_));
 sky130_fd_sc_hd__o21a_1 _381_ (.A1(\clock_div[3] ),
    .A2(_189_),
    .B1(_172_),
    .X(_029_));
 sky130_fd_sc_hd__a21oi_1 _382_ (.A1(\clock_div[4] ),
    .A2(_190_),
    .B1(net7),
    .Y(_173_));
 sky130_fd_sc_hd__o21a_1 _383_ (.A1(\clock_div[4] ),
    .A2(_190_),
    .B1(_173_),
    .X(_030_));
 sky130_fd_sc_hd__a21oi_1 _384_ (.A1(\clock_div[4] ),
    .A2(_190_),
    .B1(\clock_div[5] ),
    .Y(_174_));
 sky130_fd_sc_hd__nor3_1 _385_ (.A(net7),
    .B(_192_),
    .C(_174_),
    .Y(_031_));
 sky130_fd_sc_hd__nor2_1 _386_ (.A(net9),
    .B(_193_),
    .Y(_175_));
 sky130_fd_sc_hd__o21a_1 _387_ (.A1(\clock_div[6] ),
    .A2(_192_),
    .B1(_175_),
    .X(_032_));
 sky130_fd_sc_hd__a21o_1 _388_ (.A1(\clock_div[7] ),
    .A2(_193_),
    .B1(net9),
    .X(_176_));
 sky130_fd_sc_hd__o21ba_1 _389_ (.A1(\clock_div[7] ),
    .A2(_193_),
    .B1_N(_176_),
    .X(_033_));
 sky130_fd_sc_hd__o211a_1 _390_ (.A1(_185_),
    .A2(_195_),
    .B1(_194_),
    .C1(_187_),
    .X(_034_));
 sky130_fd_sc_hd__or4_4 _391_ (.A(net8),
    .B(_197_),
    .C(_041_),
    .D(_045_),
    .X(_177_));
 sky130_fd_sc_hd__inv_2 _392_ (.A(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__o22a_1 _393_ (.A1(\tempo_LFSR[0] ),
    .A2(_130_),
    .B1(_177_),
    .B2(\tempo_LFSR[1] ),
    .X(_035_));
 sky130_fd_sc_hd__nor2_1 _394_ (.A(_181_),
    .B(just_rst),
    .Y(_179_));
 sky130_fd_sc_hd__mux2_1 _395_ (.A0(\tempo_LFSR[1] ),
    .A1(_179_),
    .S(_130_),
    .X(_036_));
 sky130_fd_sc_hd__a2bb2o_1 _396_ (.A1_N(_181_),
    .A2_N(_130_),
    .B1(_178_),
    .B2(\tempo_LFSR[3] ),
    .X(_037_));
 sky130_fd_sc_hd__xor2_1 _397_ (.A(\tempo_LFSR[1] ),
    .B(\tempo_LFSR[0] ),
    .X(_180_));
 sky130_fd_sc_hd__o22a_1 _398_ (.A1(\tempo_LFSR[3] ),
    .A2(_130_),
    .B1(_177_),
    .B2(_180_),
    .X(_038_));
 sky130_fd_sc_hd__dfxtp_1 _399_ (.CLK(clknet_2_2__leaf_clk),
    .D(_000_),
    .Q(\tune_ROM[0] ));
 sky130_fd_sc_hd__dfxtp_1 _400_ (.CLK(clknet_2_2__leaf_clk),
    .D(_001_),
    .Q(\tune_ROM[1] ));
 sky130_fd_sc_hd__dfxtp_2 _401_ (.CLK(clknet_2_3__leaf_clk),
    .D(_002_),
    .Q(\tune_ROM[2] ));
 sky130_fd_sc_hd__dfxtp_1 _402_ (.CLK(clknet_2_3__leaf_clk),
    .D(_003_),
    .Q(\tune_ROM[3] ));
 sky130_fd_sc_hd__dfxtp_4 _403_ (.CLK(clknet_2_3__leaf_clk),
    .D(_004_),
    .Q(\tune_ROM[4] ));
 sky130_fd_sc_hd__dfxtp_1 _404_ (.CLK(clknet_2_3__leaf_clk),
    .D(_005_),
    .Q(\tune_ROM[5] ));
 sky130_fd_sc_hd__dfxtp_1 _405_ (.CLK(clknet_2_0__leaf_clk),
    .D(_006_),
    .Q(\rhythm_LFSR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _406_ (.CLK(clknet_2_2__leaf_clk),
    .D(_007_),
    .Q(\rhythm_LFSR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _407_ (.CLK(clknet_2_2__leaf_clk),
    .D(_008_),
    .Q(\rhythm_LFSR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _408_ (.CLK(clknet_2_2__leaf_clk),
    .D(_009_),
    .Q(\rhythm_LFSR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _409_ (.CLK(clknet_2_2__leaf_clk),
    .D(_010_),
    .Q(\PC[0] ));
 sky130_fd_sc_hd__dfxtp_4 _410_ (.CLK(clknet_2_2__leaf_clk),
    .D(_011_),
    .Q(\PC[1] ));
 sky130_fd_sc_hd__dfxtp_4 _411_ (.CLK(clknet_2_2__leaf_clk),
    .D(_012_),
    .Q(\PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _412_ (.CLK(clknet_2_2__leaf_clk),
    .D(net5),
    .Q(\PC[3] ));
 sky130_fd_sc_hd__dfxtp_2 _413_ (.CLK(clknet_2_2__leaf_clk),
    .D(net3),
    .Q(\PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _414_ (.CLK(clknet_2_3__leaf_clk),
    .D(_015_),
    .Q(\PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _415_ (.CLK(clknet_2_2__leaf_clk),
    .D(_016_),
    .Q(just_inc));
 sky130_fd_sc_hd__dfxtp_1 _416_ (.CLK(clknet_2_1__leaf_clk),
    .D(_017_),
    .Q(OP_reg));
 sky130_fd_sc_hd__dfxtp_1 _417_ (.CLK(clknet_2_1__leaf_clk),
    .D(_018_),
    .Q(\LFSR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _418_ (.CLK(clknet_2_1__leaf_clk),
    .D(_019_),
    .Q(\LFSR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _419_ (.CLK(clknet_2_3__leaf_clk),
    .D(_020_),
    .Q(\LFSR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _420_ (.CLK(clknet_2_1__leaf_clk),
    .D(_021_),
    .Q(\LFSR[3] ));
 sky130_fd_sc_hd__dfxtp_2 _421_ (.CLK(clknet_2_1__leaf_clk),
    .D(_022_),
    .Q(\LFSR[4] ));
 sky130_fd_sc_hd__dfxtp_2 _422_ (.CLK(clknet_2_3__leaf_clk),
    .D(_023_),
    .Q(\LFSR[5] ));
 sky130_fd_sc_hd__dfxtp_1 _423_ (.CLK(clknet_2_0__leaf_clk),
    .D(_024_),
    .Q(\LFSR[6] ));
 sky130_fd_sc_hd__dfxtp_1 _424_ (.CLK(clknet_2_3__leaf_clk),
    .D(_025_),
    .Q(prev_clk_div));
 sky130_fd_sc_hd__dfxtp_2 _425_ (.CLK(clknet_2_0__leaf_clk),
    .D(_026_),
    .Q(\clock_div[0] ));
 sky130_fd_sc_hd__dfxtp_1 _426_ (.CLK(clknet_2_1__leaf_clk),
    .D(_027_),
    .Q(\clock_div[1] ));
 sky130_fd_sc_hd__dfxtp_1 _427_ (.CLK(clknet_2_0__leaf_clk),
    .D(_028_),
    .Q(\clock_div[2] ));
 sky130_fd_sc_hd__dfxtp_1 _428_ (.CLK(clknet_2_3__leaf_clk),
    .D(_029_),
    .Q(\clock_div[3] ));
 sky130_fd_sc_hd__dfxtp_1 _429_ (.CLK(clknet_2_1__leaf_clk),
    .D(_030_),
    .Q(\clock_div[4] ));
 sky130_fd_sc_hd__dfxtp_1 _430_ (.CLK(clknet_2_3__leaf_clk),
    .D(_031_),
    .Q(\clock_div[5] ));
 sky130_fd_sc_hd__dfxtp_1 _431_ (.CLK(clknet_2_3__leaf_clk),
    .D(_032_),
    .Q(\clock_div[6] ));
 sky130_fd_sc_hd__dfxtp_2 _432_ (.CLK(clknet_2_3__leaf_clk),
    .D(_033_),
    .Q(\clock_div[7] ));
 sky130_fd_sc_hd__dfxtp_1 _433_ (.CLK(clknet_2_3__leaf_clk),
    .D(_034_),
    .Q(\clock_div[8] ));
 sky130_fd_sc_hd__dfxtp_1 _434_ (.CLK(clknet_2_0__leaf_clk),
    .D(_035_),
    .Q(\tempo_LFSR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _435_ (.CLK(clknet_2_0__leaf_clk),
    .D(_036_),
    .Q(\tempo_LFSR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _436_ (.CLK(clknet_2_0__leaf_clk),
    .D(_037_),
    .Q(\tempo_LFSR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _437_ (.CLK(clknet_2_0__leaf_clk),
    .D(_038_),
    .Q(\tempo_LFSR[3] ));
 sky130_fd_sc_hd__dfxtp_4 _438_ (.CLK(clknet_2_0__leaf_clk),
    .D(net7),
    .Q(just_rst));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__buf_4 fanout3 (.A(_014_),
    .X(net3));
 sky130_fd_sc_hd__buf_4 fanout4 (.A(net5),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 fanout5 (.A(_013_),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 fanout6 (.A(\tune_ROM[5] ),
    .X(net6));
 sky130_fd_sc_hd__buf_4 fanout7 (.A(net9),
    .X(net7));
 sky130_fd_sc_hd__buf_6 fanout8 (.A(net9),
    .X(net8));
 sky130_fd_sc_hd__buf_4 fanout9 (.A(net1),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(rst),
    .X(net1));
 sky130_fd_sc_hd__buf_4 output2 (.A(net2),
    .X(OP));
endmodule

