* NGSPICE file created from tholin_avalonsemi_tbb1143.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

.subckt tholin_avalonsemi_tbb1143 clk io_in[0] io_in[1] io_in[2] io_in[3] io_in[4]
+ io_in[5] io_out[0] io_out[1] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ rst vccd1 vssd1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_432_ _000_ clknet_1_0__leaf__213_ vssd1 vssd1 vccd1 vccd1 _090_ sky130_fd_sc_hd__xor2_2
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_501_ clknet_1_0__leaf__262_ vssd1 vssd1 vccd1 vccd1 _263_ sky130_fd_sc_hd__buf_1
XFILLER_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_415_ _196_ _197_ _198_ _199_ vssd1 vssd1 vccd1 vccd1 _200_ sky130_fd_sc_hd__or4_1
XFILLER_33_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__401__A0 _188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_964_ net20 _176_ _099_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_3.input2 sky130_fd_sc_hd__dfrtp_1
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_895_ _042_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d _041_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__631__A0 _188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_680_ _328_ vssd1 vssd1 vccd1 vccd1 _134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_947_ _093_ CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d _092_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState sky130_fd_sc_hd__dfrtp_1
X_878_ _010_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock _009_
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_801_ _369_ vssd1 vssd1 vccd1 vccd1 _167_ sky130_fd_sc_hd__clkbuf_1
X_732_ _184_ CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2 _260_ vssd1 vssd1
+ vccd1 vccd1 _343_ sky130_fd_sc_hd__mux2_1
XFILLER_43_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_663_ _320_ _319_ vssd1 vssd1 vccd1 vccd1 _004_ sky130_fd_sc_hd__nand2_1
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_594_ CIRCUIT_2223.MEMORY_25.s_currentState vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_25.d
+ sky130_fd_sc_hd__clkinv_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout20_A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_715_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState vssd1 vssd1
+ vccd1 vccd1 _046_ sky130_fd_sc_hd__clkinv_2
X_646_ slow_clock\[3\] _309_ _311_ vssd1 vssd1 vccd1 vccd1 _125_ sky130_fd_sc_hd__o21a_1
X_577_ CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d sky130_fd_sc_hd__clkinv_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_500_ net27 _243_ _256_ _261_ _117_ vssd1 vssd1 vccd1 vccd1 _262_ sky130_fd_sc_hd__o32a_2
X_431_ _000_ clknet_1_0__leaf__213_ vssd1 vssd1 vccd1 vccd1 _092_ sky130_fd_sc_hd__xor2_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_629_ net2 net1 CIRCUIT_2223.GATES_1.input1\[0\] _257_ vssd1 vssd1 vccd1 vccd1 _301_
+ sky130_fd_sc_hd__and4_2
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__236_ clknet_0__236_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__236_
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__677__D net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_414_ CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_10.input2
+ vssd1 vssd1 vccd1 vccd1 _199_ sky130_fd_sc_hd__xor2_1
XFILLER_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__405__A _191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_963_ net20 _175_ _098_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_2.input2 sky130_fd_sc_hd__dfrtp_1
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_894_ _040_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d _039_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__395__A0 _184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_946_ _091_ CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d _090_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState sky130_fd_sc_hd__dfrtp_1
X_877_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_662_ _320_ _319_ vssd1 vssd1 vccd1 vccd1 _003_ sky130_fd_sc_hd__nand2_1
X_800_ net3 CIRCUIT_2223.tone_generator_2_2.GATES_11.input2 _368_ vssd1 vssd1 vccd1
+ vccd1 _369_ sky130_fd_sc_hd__mux2_1
X_731_ _342_ vssd1 vssd1 vccd1 vccd1 _146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_593_ CIRCUIT_2223.MEMORY_26.s_currentState vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_18.clock
+ sky130_fd_sc_hd__inv_2
XFILLER_6_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_929_ net25 _155_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__770__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__761__A0 _184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput10 net10 vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_2
Xoutput8 net8 vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_645_ _306_ _310_ vssd1 vssd1 vccd1 vccd1 _311_ sky130_fd_sc_hd__nor2_1
X_714_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState vssd1 vssd1
+ vccd1 vccd1 _044_ sky130_fd_sc_hd__clkinv_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_576_ CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d sky130_fd_sc_hd__clkinv_2
XFILLER_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__743__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_430_ _000_ clknet_1_0__leaf__213_ vssd1 vssd1 vccd1 vccd1 _094_ sky130_fd_sc_hd__xor2_2
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__734__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_628_ _243_ _256_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f__235_ clknet_0__235_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__235_
+ sky130_fd_sc_hd__clkbuf_16
X_559_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d sky130_fd_sc_hd__clkinv_2
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__511__A _191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_413_ CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_15.input2
+ vssd1 vssd1 vccd1 vccd1 _198_ sky130_fd_sc_hd__xor2_1
XFILLER_33_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__506__A _191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_962_ _097_ net3 vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_893_ CIRCUIT_2223.MEMORY_24.s_currentState CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d
+ _038_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_945_ _089_ CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d _088_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState sky130_fd_sc_hd__dfrtp_1
X_876_ net20 _141_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_1.input1\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_592_ CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock sky130_fd_sc_hd__clkinv_2
X_661_ net20 vssd1 vssd1 vccd1 vccd1 _320_ sky130_fd_sc_hd__buf_2
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_730_ _186_ CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2 _260_ vssd1 vssd1
+ vccd1 vccd1 _342_ sky130_fd_sc_hd__mux2_1
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_928_ net25 _154_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_859_ net16 CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState _003_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_19_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput11 net11 vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_2
Xoutput9 net9 vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_575_ CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d sky130_fd_sc_hd__clkinv_2
X_713_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState vssd1 vssd1
+ vccd1 vccd1 _042_ sky130_fd_sc_hd__clkinv_2
X_644_ slow_clock\[0\] slow_clock\[1\] slow_clock\[2\] slow_clock\[3\] vssd1 vssd1
+ vccd1 vccd1 _310_ sky130_fd_sc_hd__and4_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__509__A _191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_627_ CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.GATES_3.result sky130_fd_sc_hd__xor2_1
X_558_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d sky130_fd_sc_hd__clkinv_2
X_489_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2
+ vssd1 vssd1 vccd1 vccd1 _251_ sky130_fd_sc_hd__xor2_1
XFILLER_12_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_412_ CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_13.input2
+ vssd1 vssd1 vccd1 vccd1 _197_ sky130_fd_sc_hd__xor2_1
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__702__A _215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1_A CIRCUIT_2223.CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_961_ _096_ net3 vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__dfxtp_1
X_892_ _037_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d _036_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_9_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__432__A _000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_944_ _087_ CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d _086_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState sky130_fd_sc_hd__dfrtp_1
X_875_ net20 _140_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_1.input1\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_591_ CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_37.d sky130_fd_sc_hd__clkinv_2
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_660_ _179_ _319_ vssd1 vssd1 vccd1 vccd1 _002_ sky130_fd_sc_hd__nand2_1
XFILLER_6_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_927_ net24 _153_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2
+ sky130_fd_sc_hd__dfxtp_1
X_858_ net17 CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState _002_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState sky130_fd_sc_hd__dfstp_1
X_789_ CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState vssd1 vssd1 vccd1
+ vccd1 _091_ sky130_fd_sc_hd__clkinv_2
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput12 net12 vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_2
XFILLER_31_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_712_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState vssd1 vssd1
+ vccd1 vccd1 _040_ sky130_fd_sc_hd__clkinv_2
X_643_ _306_ _308_ _309_ vssd1 vssd1 vccd1 vccd1 _124_ sky130_fd_sc_hd__nor3_1
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_574_ CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d sky130_fd_sc_hd__clkinv_2
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_626_ CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.GATES_2.result sky130_fd_sc_hd__xor2_1
X_557_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock sky130_fd_sc_hd__clkinv_2
XANTENNA__435__A _191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_488_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2
+ vssd1 vssd1 vccd1 vccd1 _250_ sky130_fd_sc_hd__xor2_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_411_ CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_12.input2
+ vssd1 vssd1 vccd1 vccd1 _196_ sky130_fd_sc_hd__xor2_1
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_609_ _283_ _284_ _285_ vssd1 vssd1 vccd1 vccd1 _290_ sky130_fd_sc_hd__a21bo_1
XANTENNA__398__A0 _186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_960_ net24 _174_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_7.input2
+ sky130_fd_sc_hd__dfxtp_1
X_891_ _035_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d _034_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_1__f__282_ clknet_0__282_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__282_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_943_ _085_ CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d _084_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState sky130_fd_sc_hd__dfrtp_2
X_874_ net20 _139_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_1.input1\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__773__A0 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_590_ CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_36.d sky130_fd_sc_hd__clkinv_2
XFILLER_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__764__A0 _188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_788_ CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState vssd1 vssd1 vccd1
+ vccd1 _089_ sky130_fd_sc_hd__clkinv_2
X_926_ CIRCUIT_2223.tone_generator_2_1.GATES_27.result CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState
+ sky130_fd_sc_hd__dfxtp_1
X_857_ net17 CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState _001_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_13.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_34_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput13 net13 vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_642_ slow_clock\[0\] slow_clock\[1\] slow_clock\[2\] vssd1 vssd1 vccd1 vccd1 _309_
+ sky130_fd_sc_hd__and3_1
X_711_ _191_ clknet_1_1__leaf__262_ vssd1 vssd1 vccd1 vccd1 _038_ sky130_fd_sc_hd__xnor2_2
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_573_ CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d sky130_fd_sc_hd__inv_2
XANTENNA__737__A0 _188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_909_ net23 _147_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__728__A0 _188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__541__A _215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_625_ CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.GATES_1.result sky130_fd_sc_hd__xor2_1
XANTENNA__407__C1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_556_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock sky130_fd_sc_hd__clkinv_2
X_487_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2
+ vssd1 vssd1 vccd1 vccd1 _249_ sky130_fd_sc_hd__xor2_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_410_ clknet_1_1__leaf_clk CIRCUIT_2223.GATES_11.input2 vssd1 vssd1 vccd1 vccd1 _195_
+ sky130_fd_sc_hd__nand2_2
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_608_ _287_ _288_ vssd1 vssd1 vccd1 vccd1 _289_ sky130_fd_sc_hd__or2_1
X_539_ _215_ clknet_1_1__leaf__282_ vssd1 vssd1 vccd1 vccd1 _013_ sky130_fd_sc_hd__xor2_2
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__281_ clknet_0__281_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__281_
+ sky130_fd_sc_hd__clkbuf_16
X_890_ _033_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.d _032_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_873_ net19 _138_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_1.input1\[0\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__195_ clknet_0__195_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__195_
+ sky130_fd_sc_hd__clkbuf_16
X_942_ CIRCUIT_2223.MEMORY_18.s_currentState CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d
+ _083_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_925_ _074_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock _073_ vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState sky130_fd_sc_hd__dfrtp_1
X_787_ CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState vssd1 vssd1 vccd1
+ vccd1 _087_ sky130_fd_sc_hd__inv_2
XFILLER_34_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_856_ net17 CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState _000_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_12.s_currentState sky130_fd_sc_hd__dfstp_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput14 net14 vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_2
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_572_ CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d sky130_fd_sc_hd__clkinv_2
X_641_ slow_clock\[0\] slow_clock\[1\] slow_clock\[2\] vssd1 vssd1 vccd1 vccd1 _308_
+ sky130_fd_sc_hd__a21oi_1
X_710_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState vssd1 vssd1
+ vccd1 vccd1 _037_ sky130_fd_sc_hd__clkinv_2
XANTENNA__539__A _215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__673__A0 _184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_908_ net23 _146_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2
+ sky130_fd_sc_hd__dfxtp_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_839_ clknet_1_0__leaf_clk _124_ vssd1 vssd1 vccd1 vccd1 slow_clock\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_624_ _283_ _300_ vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__nor2_1
X_555_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d sky130_fd_sc_hd__clkinv_2
XFILLER_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_486_ _244_ _245_ _246_ _247_ vssd1 vssd1 vccd1 vccd1 _248_ sky130_fd_sc_hd__a22o_1
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_607_ CIRCUIT_2223.GATES_5.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState
+ CIRCUIT_2223.GATES_4.input1\[2\] CIRCUIT_2223.s_logisimNet48 vssd1 vssd1 vccd1 vccd1
+ _288_ sky130_fd_sc_hd__a22oi_1
XANTENNA__800__A0 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_538_ _215_ clknet_1_1__leaf__282_ vssd1 vssd1 vccd1 vccd1 _015_ sky130_fd_sc_hd__xor2_2
XFILLER_32_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_469_ _237_ clknet_1_1__leaf__236_ vssd1 vssd1 vccd1 vccd1 _065_ sky130_fd_sc_hd__xnor2_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_941_ _082_ CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d _081_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_1__f__263_ clknet_0__263_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__263_
+ sky130_fd_sc_hd__clkbuf_16
X_872_ net22 _137_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_924_ _072_ CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d _071_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState sky130_fd_sc_hd__dfrtp_1
X_786_ CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState vssd1 vssd1 vccd1
+ vccd1 _085_ sky130_fd_sc_hd__inv_2
X_855_ net17 CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_11.s_currentState sky130_fd_sc_hd__dfxtp_1
XFILLER_13_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__629__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__645__A _306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput15 net15 vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_640_ slow_clock\[0\] slow_clock\[1\] _307_ vssd1 vssd1 vccd1 vccd1 _123_ sky130_fd_sc_hd__o21a_1
X_571_ CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d sky130_fd_sc_hd__clkinv_2
XFILLER_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_838_ clknet_1_0__leaf_clk _123_ vssd1 vssd1 vccd1 vccd1 slow_clock\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_907_ net23 _145_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__465__A _215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_769_ _357_ vssd1 vssd1 vccd1 vccd1 _158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__822__B _319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_623_ CIRCUIT_2223.GATES_5.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState
+ CIRCUIT_2223.GATES_4.input1\[0\] CIRCUIT_2223.s_logisimNet48 vssd1 vssd1 vccd1 vccd1
+ _300_ sky130_fd_sc_hd__a22oi_1
X_554_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d sky130_fd_sc_hd__clkinv_2
XFILLER_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_485_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2
+ vssd1 vssd1 vccd1 vccd1 _247_ sky130_fd_sc_hd__or2_1
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input6_A io_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_606_ CIRCUIT_2223.s_logisimNet48 CIRCUIT_2223.GATES_5.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState
+ CIRCUIT_2223.GATES_4.input1\[2\] vssd1 vssd1 vccd1 vccd1 _287_ sky130_fd_sc_hd__and4_1
Xclkbuf_1_0__f__213_ clknet_0__213_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__213_
+ sky130_fd_sc_hd__clkbuf_16
X_537_ _214_ clknet_1_1__leaf__282_ vssd1 vssd1 vccd1 vccd1 _017_ sky130_fd_sc_hd__xor2_2
X_468_ _237_ clknet_1_1__leaf__236_ vssd1 vssd1 vccd1 vccd1 _067_ sky130_fd_sc_hd__xnor2_2
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_399_ _187_ vssd1 vssd1 vccd1 vccd1 _176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_3_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__648__A _306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_940_ _080_ CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d _079_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState sky130_fd_sc_hd__dfrtp_1
X_871_ net22 _136_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__262_ clknet_0__262_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__262_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__236_ _236_ vssd1 vssd1 vccd1 vccd1 clknet_0__236_ sky130_fd_sc_hd__clkbuf_16
X_854_ net16 CIRCUIT_2223.tone_generator_1.GATES_3.result vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_1.MEMORY_10.s_currentState sky130_fd_sc_hd__dfxtp_1
X_923_ _070_ CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d _069_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState sky130_fd_sc_hd__dfrtp_2
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_785_ _215_ clknet_1_0__leaf__212_ vssd1 vssd1 vccd1 vccd1 _083_ sky130_fd_sc_hd__xor2_2
XFILLER_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_570_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d sky130_fd_sc_hd__clkinv_2
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_906_ net25 _144_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_10.input2
+ sky130_fd_sc_hd__dfxtp_1
X_837_ clknet_1_0__leaf_clk _122_ vssd1 vssd1 vccd1 vccd1 slow_clock\[0\] sky130_fd_sc_hd__dfxtp_1
X_768_ _184_ CIRCUIT_2223.tone_generator_2_1.GATES_13.input2 _354_ vssd1 vssd1 vccd1
+ vccd1 _357_ sky130_fd_sc_hd__mux2_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_699_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState vssd1
+ vssd1 vccd1 vccd1 _016_ sky130_fd_sc_hd__clkinv_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_622_ _298_ _299_ _297_ vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__a21o_1
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_484_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_12.input2
+ vssd1 vssd1 vccd1 vccd1 _246_ sky130_fd_sc_hd__nand2_1
XFILLER_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_553_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.d sky130_fd_sc_hd__clkinv_2
XFILLER_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_605_ _283_ _286_ vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__xnor2_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_398_ _186_ CIRCUIT_2223.GATES_3.input2 _182_ vssd1 vssd1 vccd1 vccd1 _187_ sky130_fd_sc_hd__mux2_1
X_536_ _214_ clknet_1_0__leaf__282_ vssd1 vssd1 vccd1 vccd1 _019_ sky130_fd_sc_hd__xor2_2
X_467_ _190_ vssd1 vssd1 vccd1 vccd1 _237_ sky130_fd_sc_hd__buf_8
Xclkbuf_1_0__f__212_ clknet_0__212_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__212_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_519_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2
+ vssd1 vssd1 vccd1 vccd1 _271_ sky130_fd_sc_hd__nand2_1
XFILLER_18_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_870_ net22 _135_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__749__A _191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__694__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__235_ _235_ vssd1 vssd1 vccd1 vccd1 clknet_0__235_ sky130_fd_sc_hd__clkbuf_16
XANTENNA__394__A net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__685__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_784_ CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState vssd1 vssd1 vccd1
+ vccd1 _082_ sky130_fd_sc_hd__clkinv_2
X_853_ net16 CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_9.s_currentState sky130_fd_sc_hd__dfxtp_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_922_ _068_ CIRCUIT_2223.tone_generator_2_1.MEMORY_35.d _067_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_905_ net25 _143_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_9.input2
+ sky130_fd_sc_hd__dfxtp_1
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_767_ _356_ vssd1 vssd1 vccd1 vccd1 _157_ sky130_fd_sc_hd__clkbuf_1
X_836_ net23 _121_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_698_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState vssd1
+ vssd1 vccd1 vccd1 _014_ sky130_fd_sc_hd__clkinv_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_621_ _298_ _299_ vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__xor2_1
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_552_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d sky130_fd_sc_hd__clkinv_2
X_483_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2
+ vssd1 vssd1 vccd1 vccd1 _245_ sky130_fd_sc_hd__or2_1
XFILLER_16_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_819_ _181_ _301_ vssd1 vssd1 vccd1 vccd1 _379_ sky130_fd_sc_hd__and2_1
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_604_ _284_ _285_ vssd1 vssd1 vccd1 vccd1 _286_ sky130_fd_sc_hd__nand2_1
X_535_ _214_ clknet_1_1__leaf__282_ vssd1 vssd1 vccd1 vccd1 _022_ sky130_fd_sc_hd__xor2_2
XFILLER_17_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_397_ net4 vssd1 vssd1 vccd1 vccd1 _186_ sky130_fd_sc_hd__clkbuf_4
X_466_ _215_ clknet_1_1__leaf__236_ vssd1 vssd1 vccd1 vccd1 _069_ sky130_fd_sc_hd__xnor2_2
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__397__A net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_518_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2
+ vssd1 vssd1 vccd1 vccd1 _270_ sky130_fd_sc_hd__nand2_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_449_ CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_11.input2
+ vssd1 vssd1 vccd1 vccd1 _223_ sky130_fd_sc_hd__nand2_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__664__B _319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__659__B _319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_921_ _066_ CIRCUIT_2223.tone_generator_2_1.MEMORY_34.d _065_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState sky130_fd_sc_hd__dfrtp_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_783_ CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState vssd1 vssd1 vccd1
+ vccd1 _080_ sky130_fd_sc_hd__clkinv_2
X_852_ net16 CIRCUIT_2223.tone_generator_1.GATES_2.result vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_1.MEMORY_8.s_currentState sky130_fd_sc_hd__dfxtp_1
XFILLER_19_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__389__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_904_ net24 _142_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_8.input2
+ sky130_fd_sc_hd__dfxtp_1
X_697_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState vssd1
+ vssd1 vccd1 vccd1 _012_ sky130_fd_sc_hd__clkinv_2
X_766_ _186_ CIRCUIT_2223.tone_generator_2_1.GATES_12.input2 _354_ vssd1 vssd1 vccd1
+ vccd1 _356_ sky130_fd_sc_hd__mux2_1
X_835_ net22 _120_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2
+ sky130_fd_sc_hd__dfxtp_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_620_ _287_ _294_ _291_ _292_ vssd1 vssd1 vccd1 vccd1 _299_ sky130_fd_sc_hd__o31a_1
XFILLER_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_551_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d sky130_fd_sc_hd__clkinv_2
X_482_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2
+ vssd1 vssd1 vccd1 vccd1 _244_ sky130_fd_sc_hd__nand2_1
XFILLER_16_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_818_ _378_ vssd1 vssd1 vccd1 vccd1 _096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_749_ _191_ clknet_1_1__leaf__235_ vssd1 vssd1 vccd1 vccd1 _062_ sky130_fd_sc_hd__xnor2_2
XFILLER_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__667__B _319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__730__A0 _186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_603_ CIRCUIT_2223.s_logisimNet48 CIRCUIT_2223.GATES_5.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState
+ CIRCUIT_2223.GATES_4.input1\[1\] vssd1 vssd1 vccd1 vccd1 _285_ sky130_fd_sc_hd__nand4_1
XFILLER_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_534_ _214_ clknet_1_0__leaf__282_ vssd1 vssd1 vccd1 vccd1 _024_ sky130_fd_sc_hd__xor2_2
X_465_ _215_ clknet_1_0__leaf__236_ vssd1 vssd1 vccd1 vccd1 _071_ sky130_fd_sc_hd__xnor2_2
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__797__A0 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_396_ _185_ vssd1 vssd1 vccd1 vccd1 _177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A io_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__779__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout20 net21 vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_2
XFILLER_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_517_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2
+ vssd1 vssd1 vccd1 vccd1 _269_ sky130_fd_sc_hd__or2_1
X_448_ CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_17.input2
+ vssd1 vssd1 vccd1 vccd1 _222_ sky130_fd_sc_hd__nand2_1
XFILLER_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_851_ net16 CIRCUIT_2223.tone_generator_1.GATES_1.result vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_1.MEMORY_7.s_currentState sky130_fd_sc_hd__dfxtp_1
X_920_ _064_ CIRCUIT_2223.tone_generator_2_1.MEMORY_33.d _063_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_782_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState vssd1 vssd1 vccd1
+ vccd1 _078_ sky130_fd_sc_hd__clkinv_2
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout25_A CIRCUIT_2223.CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_903_ _053_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.clock vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState sky130_fd_sc_hd__dfxtp_1
X_834_ net22 _119_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2
+ sky130_fd_sc_hd__dfxtp_1
X_696_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState vssd1
+ vssd1 vccd1 vccd1 _010_ sky130_fd_sc_hd__clkinv_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_765_ _355_ vssd1 vssd1 vccd1 vccd1 _156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_550_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d sky130_fd_sc_hd__clkinv_2
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_481_ _238_ _239_ _240_ _241_ _242_ vssd1 vssd1 vccd1 vccd1 _243_ sky130_fd_sc_hd__a221o_1
XFILLER_8_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_817_ _181_ _326_ vssd1 vssd1 vccd1 vccd1 _378_ sky130_fd_sc_hd__and2_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_748_ CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState vssd1 vssd1 vccd1
+ vccd1 _061_ sky130_fd_sc_hd__clkinv_2
X_679_ _188_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2 _327_
+ vssd1 vssd1 vccd1 vccd1 _328_ sky130_fd_sc_hd__mux2_1
X_602_ CIRCUIT_2223.GATES_5.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState
+ CIRCUIT_2223.GATES_4.input1\[1\] CIRCUIT_2223.s_logisimNet48 vssd1 vssd1 vccd1 vccd1
+ _284_ sky130_fd_sc_hd__a22o_1
XFILLER_43_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_464_ _215_ clknet_1_0__leaf__236_ vssd1 vssd1 vccd1 vccd1 _073_ sky130_fd_sc_hd__xnor2_2
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_533_ _214_ clknet_1_0__leaf__282_ vssd1 vssd1 vccd1 vccd1 _026_ sky130_fd_sc_hd__xor2_2
XFILLER_43_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_395_ _184_ CIRCUIT_2223.GATES_5.input2 _182_ vssd1 vssd1 vccd1 vccd1 _185_ sky130_fd_sc_hd__mux2_1
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout21 net28 vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_447_ CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_17.input2
+ vssd1 vssd1 vccd1 vccd1 _221_ sky130_fd_sc_hd__or2_1
X_516_ _264_ _265_ _266_ _267_ vssd1 vssd1 vccd1 vccd1 _268_ sky130_fd_sc_hd__or4_1
XFILLER_9_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__688__A0 _188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__679__A0 _188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_781_ CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState vssd1 vssd1 vccd1
+ vccd1 _076_ sky130_fd_sc_hd__clkinv_2
X_850_ net16 CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_6.s_currentState sky130_fd_sc_hd__dfxtp_1
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout18_A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_902_ _052_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.clock vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState sky130_fd_sc_hd__dfxtp_1
XANTENNA__815__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_764_ _188_ CIRCUIT_2223.tone_generator_2_1.GATES_11.input2 _354_ vssd1 vssd1 vccd1
+ vccd1 _355_ sky130_fd_sc_hd__mux2_1
X_833_ CIRCUIT_2223.MEMORY_26.s_currentState vssd1 vssd1 vccd1 vccd1 _118_ sky130_fd_sc_hd__clkinv_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_695_ _336_ vssd1 vssd1 vccd1 vccd1 _141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__806__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_480_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2
+ vssd1 vssd1 vccd1 vccd1 _242_ sky130_fd_sc_hd__xor2_1
XFILLER_32_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_816_ _377_ vssd1 vssd1 vccd1 vccd1 _174_ sky130_fd_sc_hd__clkbuf_1
X_747_ CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState vssd1 vssd1 vccd1
+ vccd1 _059_ sky130_fd_sc_hd__clkinv_2
XANTENNA__400__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_678_ _259_ _326_ vssd1 vssd1 vccd1 vccd1 _327_ sky130_fd_sc_hd__nand2_1
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_601_ CIRCUIT_2223.s_logisimNet48 CIRCUIT_2223.GATES_5.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState
+ CIRCUIT_2223.GATES_4.input1\[0\] vssd1 vssd1 vccd1 vccd1 _283_ sky130_fd_sc_hd__and4_1
XFILLER_17_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_463_ clknet_1_0__leaf__235_ vssd1 vssd1 vccd1 vccd1 _236_ sky130_fd_sc_hd__buf_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_394_ net5 vssd1 vssd1 vccd1 vccd1 _184_ sky130_fd_sc_hd__clkbuf_4
X_532_ _000_ clknet_1_0__leaf__282_ vssd1 vssd1 vccd1 vccd1 _028_ sky130_fd_sc_hd__xor2_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout22 net23 vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_515_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2
+ vssd1 vssd1 vccd1 vccd1 _267_ sky130_fd_sc_hd__xor2_1
XFILLER_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_446_ _216_ _217_ _218_ _219_ vssd1 vssd1 vccd1 vccd1 _220_ sky130_fd_sc_hd__or4_1
XFILLER_10_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_429_ clknet_1_1__leaf__212_ vssd1 vssd1 vccd1 vccd1 _213_ sky130_fd_sc_hd__buf_1
XFILLER_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput1 io_in[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_4
XTAP_90 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_780_ _363_ vssd1 vssd1 vccd1 vccd1 _163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_42_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_901_ _051_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.d vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState sky130_fd_sc_hd__dfxtp_1
XFILLER_21_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_763_ _193_ _233_ vssd1 vssd1 vccd1 vccd1 _354_ sky130_fd_sc_hd__nand2_2
X_832_ CIRCUIT_2223.MEMORY_18.s_currentState vssd1 vssd1 vccd1 vccd1 _116_ sky130_fd_sc_hd__clkinv_2
X_694_ net6 CIRCUIT_2223.GATES_1.input1\[3\] _332_ vssd1 vssd1 vccd1 vccd1 _336_ sky130_fd_sc_hd__mux2_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_815_ net6 CIRCUIT_2223.tone_generator_2_2.GATES_7.input2 _373_ vssd1 vssd1 vccd1
+ vccd1 _377_ sky130_fd_sc_hd__mux2_1
X_746_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState vssd1 vssd1 vccd1
+ vccd1 _057_ sky130_fd_sc_hd__clkinv_2
X_677_ CIRCUIT_2223.GATES_1.input1\[0\] CIRCUIT_2223.GATES_1.input1\[1\] net2 net1
+ vssd1 vssd1 vccd1 vccd1 _326_ sky130_fd_sc_hd__and4b_2
XANTENNA__724__A0 _186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_600_ CIRCUIT_2223.MEMORY_18.s_currentState vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_18.d
+ sky130_fd_sc_hd__clkinv_2
XFILLER_27_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_531_ clknet_1_1__leaf__281_ vssd1 vssd1 vccd1 vccd1 _282_ sky130_fd_sc_hd__buf_1
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_393_ _183_ vssd1 vssd1 vccd1 vccd1 _178_ sky130_fd_sc_hd__clkbuf_1
X_462_ clknet_1_0__leaf__195_ CIRCUIT_2223.tone_generator_2_1.GATES_27.result _234_
+ vssd1 vssd1 vccd1 vccd1 _235_ sky130_fd_sc_hd__a21oi_2
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_729_ _341_ vssd1 vssd1 vccd1 vccd1 _145_ sky130_fd_sc_hd__clkbuf_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout23 CIRCUIT_2223.CLK vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_514_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2
+ vssd1 vssd1 vccd1 vccd1 _266_ sky130_fd_sc_hd__xor2_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_445_ CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_13.input2
+ vssd1 vssd1 vccd1 vccd1 _219_ sky130_fd_sc_hd__xor2_1
XANTENNA__961__D net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input2_A io_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_428_ net24 _192_ _194_ clknet_1_1__leaf__195_ CIRCUIT_2223.tone_generator_2_2.GATES_27.result
+ vssd1 vssd1 vccd1 vccd1 _212_ sky130_fd_sc_hd__a32o_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 io_in[1] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_4
XTAP_91 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__213_ _213_ vssd1 vssd1 vccd1 vccd1 clknet_0__213_ sky130_fd_sc_hd__clkbuf_16
X_900_ CIRCUIT_2223.triangle_wave_generator_1.GATES_27.result CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.d
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState
+ sky130_fd_sc_hd__dfxtp_1
X_831_ CIRCUIT_2223.MEMORY_19.s_currentState vssd1 vssd1 vccd1 vccd1 _114_ sky130_fd_sc_hd__clkinv_2
X_762_ _353_ vssd1 vssd1 vccd1 vccd1 _155_ sky130_fd_sc_hd__clkbuf_1
X_693_ _335_ vssd1 vssd1 vccd1 vccd1 _140_ sky130_fd_sc_hd__clkbuf_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout23_A CIRCUIT_2223.CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_814_ _376_ vssd1 vssd1 vccd1 vccd1 _173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_745_ CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState vssd1 vssd1 vccd1
+ vccd1 _055_ sky130_fd_sc_hd__inv_2
X_676_ _325_ vssd1 vssd1 vccd1 vccd1 _133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_461_ _180_ _233_ net19 vssd1 vssd1 vccd1 vccd1 _234_ sky130_fd_sc_hd__and3b_1
X_530_ clknet_1_1__leaf__195_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result
+ _280_ net24 vssd1 vssd1 vccd1 vccd1 _281_ sky130_fd_sc_hd__a22o_2
XFILLER_43_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_392_ net6 CIRCUIT_2223.s_logisimNet48 _182_ vssd1 vssd1 vccd1 vccd1 _183_ sky130_fd_sc_hd__mux2_1
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_728_ _188_ CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2 _260_ vssd1 vssd1
+ vccd1 vccd1 _341_ sky130_fd_sc_hd__mux2_1
X_659_ _179_ _319_ vssd1 vssd1 vccd1 vccd1 _001_ sky130_fd_sc_hd__nand2_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__633__A0 _186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout24 CIRCUIT_2223.CLK vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_513_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2
+ vssd1 vssd1 vccd1 vccd1 _265_ sky130_fd_sc_hd__xor2_1
X_444_ CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_15.input2
+ vssd1 vssd1 vccd1 vccd1 _218_ sky130_fd_sc_hd__xor2_1
XFILLER_13_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__507__A _191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_427_ _200_ _206_ _211_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_27.result
+ sky130_fd_sc_hd__nor3_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_92 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 io_in[2] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__buf_2
XFILLER_27_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__809__A0 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__212_ _212_ vssd1 vssd1 vccd1 vccd1 clknet_0__212_ sky130_fd_sc_hd__clkbuf_16
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_761_ _184_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_10.input2 _350_
+ vssd1 vssd1 vccd1 vccd1 _353_ sky130_fd_sc_hd__mux2_1
X_830_ CIRCUIT_2223.MEMORY_20.s_currentState vssd1 vssd1 vccd1 vccd1 _112_ sky130_fd_sc_hd__clkinv_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_692_ _184_ CIRCUIT_2223.GATES_1.input1\[2\] _332_ vssd1 vssd1 vccd1 vccd1 _335_
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__430__A _000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_959_ net24 _173_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_17.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_813_ net5 CIRCUIT_2223.tone_generator_2_2.GATES_17.input2 _373_ vssd1 vssd1 vccd1
+ vccd1 _376_ sky130_fd_sc_hd__mux2_1
X_744_ _349_ vssd1 vssd1 vccd1 vccd1 _152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_675_ net6 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2 _321_
+ vssd1 vssd1 vccd1 vccd1 _325_ sky130_fd_sc_hd__mux2_1
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__282_ clknet_0__282_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__282_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_460_ _232_ vssd1 vssd1 vccd1 vccd1 _233_ sky130_fd_sc_hd__clkbuf_2
XFILLER_27_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_391_ _180_ _181_ vssd1 vssd1 vccd1 vccd1 _182_ sky130_fd_sc_hd__nand2_2
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_727_ _340_ vssd1 vssd1 vccd1 vccd1 _144_ sky130_fd_sc_hd__clkbuf_1
X_589_ CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_35.d sky130_fd_sc_hd__clkinv_2
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_658_ net7 vssd1 vssd1 vccd1 vccd1 _319_ sky130_fd_sc_hd__buf_2
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout25 CIRCUIT_2223.CLK vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_443_ CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_10.input2
+ vssd1 vssd1 vccd1 vccd1 _217_ sky130_fd_sc_hd__xor2_1
X_512_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2
+ vssd1 vssd1 vccd1 vccd1 _264_ sky130_fd_sc_hd__xor2_1
XFILLER_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_426_ _207_ _208_ _209_ _210_ vssd1 vssd1 vccd1 vccd1 _211_ sky130_fd_sc_hd__or4_1
XANTENNA__433__A _000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput4 io_in[3] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_93 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_975_ _118_ CIRCUIT_2223.MEMORY_18.d _117_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_18.s_currentState
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_409_ CIRCUIT_2223.MEMORY_23.s_currentState vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_11.input2
+ sky130_fd_sc_hd__inv_2
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_760_ _352_ vssd1 vssd1 vccd1 vccd1 _154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_691_ _334_ vssd1 vssd1 vccd1 vccd1 _139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__711__A _191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_958_ net24 _172_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_16.input2
+ sky130_fd_sc_hd__dfxtp_1
X_889_ _031_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.d _030_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState sky130_fd_sc_hd__dfrtp_2
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_812_ _375_ vssd1 vssd1 vccd1 vccd1 _172_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__406__C1 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_743_ net6 CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2 _345_ vssd1 vssd1
+ vccd1 vccd1 _349_ sky130_fd_sc_hd__mux2_1
X_674_ _324_ vssd1 vssd1 vccd1 vccd1 _132_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__281_ clknet_0__281_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__281_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_390_ net2 net1 CIRCUIT_2223.GATES_1.input1\[2\] CIRCUIT_2223.GATES_1.input1\[3\]
+ vssd1 vssd1 vccd1 vccd1 _181_ sky130_fd_sc_hd__and4_1
XFILLER_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_726_ _184_ CIRCUIT_2223.tone_generator_2_2.GATES_10.input2 _337_ vssd1 vssd1 vccd1
+ vccd1 _340_ sky130_fd_sc_hd__mux2_1
X_657_ net18 _316_ _318_ vssd1 vssd1 vccd1 vccd1 _129_ sky130_fd_sc_hd__o21a_1
X_588_ CIRCUIT_2223.tone_generator_2_2.MEMORY_34.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_34.d sky130_fd_sc_hd__clkinv_2
Xclkbuf_1_0__f__195_ clknet_0__195_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__195_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_511_ _191_ clknet_1_1__leaf__263_ vssd1 vssd1 vccd1 vccd1 _030_ sky130_fd_sc_hd__xnor2_2
X_442_ CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_12.input2
+ vssd1 vssd1 vccd1 vccd1 _216_ sky130_fd_sc_hd__xor2_1
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_709_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState vssd1 vssd1
+ vccd1 vccd1 _035_ sky130_fd_sc_hd__clkinv_2
XFILLER_24_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_425_ CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_16.input2
+ vssd1 vssd1 vccd1 vccd1 _210_ sky130_fd_sc_hd__xor2_1
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 io_in[4] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__buf_2
XTAP_94 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_974_ _116_ CIRCUIT_2223.MEMORY_19.d _115_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_19.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_408_ _193_ vssd1 vssd1 vccd1 vccd1 _194_ sky130_fd_sc_hd__inv_2
XANTENNA__953__CLK net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__690__A0 _186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_690_ _186_ CIRCUIT_2223.GATES_1.input1\[1\] _332_ vssd1 vssd1 vccd1 vccd1 _334_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__681__A0 _186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_957_ net24 _171_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_15.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_888_ _029_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.d _028_ vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_811_ net4 CIRCUIT_2223.tone_generator_2_2.GATES_16.input2 _373_ vssd1 vssd1 vccd1
+ vccd1 _375_ sky130_fd_sc_hd__mux2_1
X_742_ _348_ vssd1 vssd1 vccd1 vccd1 _151_ sky130_fd_sc_hd__clkbuf_1
X_673_ _184_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2 _321_
+ vssd1 vssd1 vccd1 vccd1 _324_ sky130_fd_sc_hd__mux2_1
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_725_ _339_ vssd1 vssd1 vccd1 vccd1 _143_ sky130_fd_sc_hd__clkbuf_1
X_587_ CIRCUIT_2223.tone_generator_2_2.MEMORY_33.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_33.d sky130_fd_sc_hd__clkinv_2
X_656_ net18 _316_ _306_ vssd1 vssd1 vccd1 vccd1 _318_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__263_ clknet_0__263_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__263_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout16 net17 vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_441_ _190_ vssd1 vssd1 vccd1 vccd1 _215_ sky130_fd_sc_hd__clkbuf_16
X_510_ _191_ clknet_1_1__leaf__263_ vssd1 vssd1 vccd1 vccd1 _032_ sky130_fd_sc_hd__xnor2_2
XFILLER_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_639_ slow_clock\[0\] slow_clock\[1\] _306_ vssd1 vssd1 vccd1 vccd1 _307_ sky130_fd_sc_hd__a21oi_1
X_708_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState vssd1 vssd1
+ vccd1 vccd1 _033_ sky130_fd_sc_hd__clkinv_2
XFILLER_6_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_424_ CIRCUIT_2223.tone_generator_2_2.MEMORY_35.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_14.input2
+ vssd1 vssd1 vccd1 vccd1 _209_ sky130_fd_sc_hd__xor2_1
Xinput6 io_in[5] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_4
XFILLER_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_95 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_973_ _114_ CIRCUIT_2223.MEMORY_20.d _113_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_20.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_407_ CIRCUIT_2223.GATES_1.input1\[0\] CIRCUIT_2223.GATES_1.input1\[1\] net2 net1
+ vssd1 vssd1 vccd1 vccd1 _193_ sky130_fd_sc_hd__o211ai_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_956_ net21 _170_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_14.input2
+ sky130_fd_sc_hd__dfxtp_1
X_887_ _027_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.d _026_ vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_810_ _374_ vssd1 vssd1 vccd1 vccd1 _171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_672_ _323_ vssd1 vssd1 vccd1 vccd1 _131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_741_ _184_ CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2 _345_ vssd1 vssd1
+ vccd1 vccd1 _348_ sky130_fd_sc_hd__mux2_1
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_939_ _078_ CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d _077_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState sky130_fd_sc_hd__dfrtp_2
XFILLER_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_724_ _186_ CIRCUIT_2223.tone_generator_2_2.GATES_9.input2 _337_ vssd1 vssd1 vccd1
+ vccd1 _339_ sky130_fd_sc_hd__mux2_1
XFILLER_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_586_ CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_32.d sky130_fd_sc_hd__inv_2
X_655_ slow_clock\[6\] _314_ _317_ vssd1 vssd1 vccd1 vccd1 _128_ sky130_fd_sc_hd__o21a_1
XFILLER_16_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__262_ clknet_0__262_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__262_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__643__A _306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout17 CIRCUIT_2223.MEMORY_24.s_currentState vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_2
XFILLER_22_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_440_ _214_ clknet_1_1__leaf__213_ vssd1 vssd1 vccd1 vccd1 _075_ sky130_fd_sc_hd__xor2_2
XANTENNA__793__A0 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_707_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState vssd1 vssd1
+ vccd1 vccd1 _031_ sky130_fd_sc_hd__clkinv_2
X_569_ CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_39.d sky130_fd_sc_hd__clkinv_2
X_638_ slow_clock\[0\] _306_ vssd1 vssd1 vccd1 vccd1 _122_ sky130_fd_sc_hd__nor2_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__775__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_423_ CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_9.input2
+ vssd1 vssd1 vccd1 vccd1 _208_ sky130_fd_sc_hd__xor2_1
XANTENNA__766__A0 _186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__757__A0 _188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 rst vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XTAP_96 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_972_ _112_ CIRCUIT_2223.MEMORY_21.d _111_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_21.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__739__A0 _186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_406_ CIRCUIT_2223.GATES_1.input1\[2\] CIRCUIT_2223.GATES_1.input1\[3\] net2 net1
+ vssd1 vssd1 vccd1 vccd1 _192_ sky130_fd_sc_hd__o211ai_4
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__651__A _306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_955_ net21 _169_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_13.input2
+ sky130_fd_sc_hd__dfxtp_1
X_886_ _025_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.d _024_ vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_740_ _347_ vssd1 vssd1 vccd1 vccd1 _150_ sky130_fd_sc_hd__clkbuf_1
X_671_ _186_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2 _321_
+ vssd1 vssd1 vccd1 vccd1 _323_ sky130_fd_sc_hd__mux2_1
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_938_ _076_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d _075_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState sky130_fd_sc_hd__dfrtp_1
X_869_ net23 _134_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__466__A _215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__823__B _306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_723_ _338_ vssd1 vssd1 vccd1 vccd1 _142_ sky130_fd_sc_hd__clkbuf_1
X_654_ _306_ _316_ vssd1 vssd1 vccd1 vccd1 _317_ sky130_fd_sc_hd__nor2_1
X_585_ CIRCUIT_2223.tone_generator_2_2.MEMORY_31.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_31.d sky130_fd_sc_hd__clkinv_2
XFILLER_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout18 net21 vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__buf_2
XFILLER_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_706_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState vssd1
+ vssd1 vccd1 vccd1 _029_ sky130_fd_sc_hd__clkinv_2
X_637_ net7 vssd1 vssd1 vccd1 vccd1 _306_ sky130_fd_sc_hd__buf_2
XANTENNA__956__CLK net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_568_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock sky130_fd_sc_hd__clkinv_2
X_499_ _257_ _259_ _260_ vssd1 vssd1 vccd1 vccd1 _261_ sky130_fd_sc_hd__a21boi_1
XFILLER_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__654__A _306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__638__B _306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_422_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_7.input2
+ vssd1 vssd1 vccd1 vccd1 _207_ sky130_fd_sc_hd__xor2_1
XFILLER_5_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_97 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_971_ _110_ CIRCUIT_2223.MEMORY_22.d _109_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_22.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_405_ _191_ vssd1 vssd1 vccd1 vccd1 _000_ sky130_fd_sc_hd__buf_6
XFILLER_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__675__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_954_ net20 _168_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_12.input2
+ sky130_fd_sc_hd__dfxtp_1
X_885_ _023_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d _022_ vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__639__B1 _306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_670_ _322_ vssd1 vssd1 vccd1 vccd1 _130_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__811__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__802__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_799_ _192_ _301_ vssd1 vssd1 vccd1 vccd1 _368_ sky130_fd_sc_hd__nand2_1
X_937_ net18 _163_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_7.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_868_ net24 _133_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_722_ _188_ CIRCUIT_2223.tone_generator_2_2.GATES_8.input2 _337_ vssd1 vssd1 vccd1
+ vccd1 _338_ sky130_fd_sc_hd__mux2_1
X_653_ slow_clock\[6\] _314_ vssd1 vssd1 vccd1 vccd1 _316_ sky130_fd_sc_hd__and2_1
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_584_ CIRCUIT_2223.tone_generator_2_2.MEMORY_30.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_30.d sky130_fd_sc_hd__clkinv_2
XFILLER_31_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout19 net21 vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_705_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState vssd1
+ vssd1 vccd1 vccd1 _027_ sky130_fd_sc_hd__clkinv_2
X_567_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d sky130_fd_sc_hd__clkinv_2
X_636_ _305_ vssd1 vssd1 vccd1 vccd1 _121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_498_ _180_ _233_ vssd1 vssd1 vccd1 vccd1 _260_ sky130_fd_sc_hd__nand2_2
XFILLER_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_421_ _201_ _202_ _203_ _204_ _205_ vssd1 vssd1 vccd1 vccd1 _206_ sky130_fd_sc_hd__a221o_1
XFILLER_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_619_ _296_ _297_ vssd1 vssd1 vccd1 vccd1 _298_ sky130_fd_sc_hd__nor2_1
XFILLER_36_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_98 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_970_ _108_ CIRCUIT_2223.GATES_11.input2 _107_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_23.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_404_ _190_ vssd1 vssd1 vccd1 vccd1 _191_ sky130_fd_sc_hd__buf_8
XFILLER_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_953_ net21 _167_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.GATES_11.input2
+ sky130_fd_sc_hd__dfxtp_1
X_884_ CIRCUIT_2223.MEMORY_24.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d
+ _021_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__662__B _319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_936_ net18 _162_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_17.input2
+ sky130_fd_sc_hd__dfxtp_1
X_798_ _367_ vssd1 vssd1 vccd1 vccd1 _166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_867_ net24 _132_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_583_ CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_29.d sky130_fd_sc_hd__clkinv_2
X_721_ _180_ _192_ vssd1 vssd1 vccd1 vccd1 _337_ sky130_fd_sc_hd__nand2_1
X_652_ slow_clock\[5\] _312_ _315_ vssd1 vssd1 vccd1 vccd1 _127_ sky130_fd_sc_hd__o21a_1
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 CIRCUIT_2223.CLK vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dlygate4sd3_1
X_919_ CIRCUIT_2223.MEMORY_18.s_currentState CIRCUIT_2223.tone_generator_2_1.MEMORY_32.d
+ _062_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState
+ sky130_fd_sc_hd__dfrtp_2
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_704_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_29.s_currentState vssd1
+ vssd1 vccd1 vccd1 _025_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_566_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d sky130_fd_sc_hd__clkinv_2
X_635_ _184_ CIRCUIT_2223.triangle_wave_generator_1.GATES_10.input2 _302_ vssd1 vssd1
+ vccd1 vccd1 _305_ sky130_fd_sc_hd__mux2_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_497_ _258_ vssd1 vssd1 vccd1 vccd1 _259_ sky130_fd_sc_hd__clkbuf_2
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_420_ CIRCUIT_2223.tone_generator_2_2.MEMORY_32.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_11.input2
+ vssd1 vssd1 vccd1 vccd1 _205_ sky130_fd_sc_hd__xor2_1
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_549_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_31.d sky130_fd_sc_hd__clkinv_2
X_618_ CIRCUIT_2223.GATES_3.input2 CIRCUIT_2223.GATES_2.input2 CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState vssd1 vssd1 vccd1 vccd1
+ _297_ sky130_fd_sc_hd__and4_1
XTAP_99 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__665__B _319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0__282_ _282_ vssd1 vssd1 vccd1 vccd1 clknet_0__282_ sky130_fd_sc_hd__clkbuf_16
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_403_ net18 net7 vssd1 vssd1 vccd1 vccd1 _190_ sky130_fd_sc_hd__nand2_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_952_ net19 _166_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_10.input2
+ sky130_fd_sc_hd__dfxtp_1
X_883_ _020_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d _019_ vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_935_ net18 _161_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_16.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_866_ net25 _131_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2
+ sky130_fd_sc_hd__dfxtp_1
X_797_ net5 CIRCUIT_2223.tone_generator_2_1.GATES_10.input2 _364_ vssd1 vssd1 vccd1
+ vccd1 _367_ sky130_fd_sc_hd__mux2_1
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_720_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_39.s_currentState vssd1 vssd1
+ vccd1 vccd1 _053_ sky130_fd_sc_hd__clkinv_2
X_582_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_28.d sky130_fd_sc_hd__clkinv_2
X_651_ _306_ _314_ vssd1 vssd1 vccd1 vccd1 _315_ sky130_fd_sc_hd__nor2_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_849_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState CIRCUIT_2223.tone_generator_1.MEMORY_14.s_currentState
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_4.input1\[3\] sky130_fd_sc_hd__dfxtp_1
X_918_ _061_ CIRCUIT_2223.tone_generator_2_1.MEMORY_31.d _060_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_31.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_703_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState vssd1
+ vssd1 vccd1 vccd1 _023_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_634_ _304_ vssd1 vssd1 vccd1 vccd1 _120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_565_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d sky130_fd_sc_hd__clkinv_2
X_496_ CIRCUIT_2223.GATES_1.input1\[2\] CIRCUIT_2223.GATES_1.input1\[3\] net2 net1
+ vssd1 vssd1 vccd1 vccd1 _258_ sky130_fd_sc_hd__and4b_1
XFILLER_8_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_617_ CIRCUIT_2223.GATES_3.input2 CIRCUIT_2223.tone_generator_2_1.MEMORY_39.s_currentState
+ CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState CIRCUIT_2223.GATES_2.input2
+ vssd1 vssd1 vccd1 vccd1 _296_ sky130_fd_sc_hd__a22oi_1
X_548_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.d sky130_fd_sc_hd__clkinv_2
X_479_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2
+ vssd1 vssd1 vccd1 vccd1 _241_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__281_ _281_ vssd1 vssd1 vccd1 vccd1 clknet_0__281_ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__669__A0 _188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_402_ _189_ vssd1 vssd1 vccd1 vccd1 _175_ sky130_fd_sc_hd__clkbuf_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_0__195_ _195_ vssd1 vssd1 vccd1 vccd1 clknet_0__195_ sky130_fd_sc_hd__clkbuf_16
XFILLER_11_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_882_ _018_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d _017_ vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState
+ sky130_fd_sc_hd__dfrtp_2
X_951_ net18 _165_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_9.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__687__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_934_ net18 _160_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_15.input2
+ sky130_fd_sc_hd__dfxtp_1
X_796_ _366_ vssd1 vssd1 vccd1 vccd1 _165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_865_ net22 _130_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_650_ slow_clock\[4\] slow_clock\[5\] _310_ vssd1 vssd1 vccd1 vccd1 _314_ sky130_fd_sc_hd__and3_1
X_581_ CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d sky130_fd_sc_hd__clkinv_2
XFILLER_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_848_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_4.input1\[2\] sky130_fd_sc_hd__dfxtp_1
X_917_ _059_ CIRCUIT_2223.tone_generator_2_1.MEMORY_30.d _058_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState sky130_fd_sc_hd__dfrtp_2
X_779_ net6 CIRCUIT_2223.tone_generator_2_1.GATES_7.input2 _359_ vssd1 vssd1 vccd1
+ vccd1 _363_ sky130_fd_sc_hd__mux2_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_633_ _186_ CIRCUIT_2223.triangle_wave_generator_1.GATES_9.input2 _302_ vssd1 vssd1
+ vccd1 vccd1 _304_ sky130_fd_sc_hd__mux2_1
X_702_ _215_ clknet_1_0__leaf__281_ vssd1 vssd1 vccd1 vccd1 _021_ sky130_fd_sc_hd__xor2_2
X_564_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.d sky130_fd_sc_hd__clkinv_2
XFILLER_8_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_495_ CIRCUIT_2223.GATES_1.input1\[1\] vssd1 vssd1 vccd1 vccd1 _257_ sky130_fd_sc_hd__inv_2
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__785__A _215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input7_A rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_616_ _293_ _295_ vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__xnor2_1
X_547_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.d sky130_fd_sc_hd__inv_2
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_478_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2
+ vssd1 vssd1 vccd1 vccd1 _240_ sky130_fd_sc_hd__or2_1
XFILLER_35_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_401_ _188_ CIRCUIT_2223.GATES_2.input2 _182_ vssd1 vssd1 vccd1 vccd1 _189_ sky130_fd_sc_hd__mux2_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__263_ _263_ vssd1 vssd1 vccd1 vccd1 clknet_0__263_ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_950_ net18 _164_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_8.input2
+ sky130_fd_sc_hd__dfxtp_1
X_881_ _016_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d _015_ vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_36_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__741__A0 _184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__732__A0 _184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_933_ net19 _159_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_14.input2
+ sky130_fd_sc_hd__dfxtp_1
X_864_ net16 CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState _008_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState sky130_fd_sc_hd__dfrtp_2
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_795_ net4 CIRCUIT_2223.tone_generator_2_1.GATES_9.input2 _364_ vssd1 vssd1 vccd1
+ vccd1 _366_ sky130_fd_sc_hd__mux2_1
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_580_ CIRCUIT_2223.tone_generator_2_1.MEMORY_38.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_28.clock sky130_fd_sc_hd__clkinv_2
XFILLER_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_916_ _057_ CIRCUIT_2223.tone_generator_2_1.MEMORY_29.d _056_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState sky130_fd_sc_hd__dfrtp_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_847_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_4.input1\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_778_ _362_ vssd1 vssd1 vccd1 vccd1 _162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_701_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState vssd1
+ vssd1 vccd1 vccd1 _020_ sky130_fd_sc_hd__inv_2
XFILLER_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_563_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_33.d sky130_fd_sc_hd__clkinv_2
X_632_ _303_ vssd1 vssd1 vccd1 vccd1 _119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_494_ _248_ _249_ _250_ _255_ vssd1 vssd1 vccd1 vccd1 _256_ sky130_fd_sc_hd__or4_1
XFILLER_12_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_615_ _287_ _294_ vssd1 vssd1 vccd1 vccd1 _295_ sky130_fd_sc_hd__nor2_1
X_546_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_34.d sky130_fd_sc_hd__clkinv_2
X_477_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2
+ vssd1 vssd1 vccd1 vccd1 _239_ sky130_fd_sc_hd__or2_1
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_400_ net3 vssd1 vssd1 vccd1 vccd1 _188_ sky130_fd_sc_hd__buf_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_529_ _181_ _193_ _259_ CIRCUIT_2223.GATES_1.input1\[1\] vssd1 vssd1 vccd1 vccd1
+ _280_ sky130_fd_sc_hd__a22o_1
XFILLER_17_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__262_ _262_ vssd1 vssd1 vccd1 vccd1 clknet_0__262_ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_880_ _014_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d _013_ vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__496__D net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_863_ net16 CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState _007_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_19.s_currentState sky130_fd_sc_hd__dfstp_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_932_ net19 _158_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_13.input2
+ sky130_fd_sc_hd__dfxtp_1
X_794_ _365_ vssd1 vssd1 vccd1 vccd1 _164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_846_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_39.s_currentState CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_4.input1\[0\] sky130_fd_sc_hd__dfxtp_1
X_915_ _055_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.d _054_ vssd1 vssd1 vccd1 vccd1
+ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState sky130_fd_sc_hd__dfrtp_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_777_ net5 CIRCUIT_2223.tone_generator_2_1.GATES_17.input2 _359_ vssd1 vssd1 vccd1
+ vccd1 _362_ sky130_fd_sc_hd__mux2_1
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_700_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_33.s_currentState vssd1
+ vssd1 vccd1 vccd1 _018_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__502__A _215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_493_ _251_ _252_ _253_ _254_ vssd1 vssd1 vccd1 vccd1 _255_ sky130_fd_sc_hd__or4_1
X_631_ _188_ CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2 _302_ vssd1 vssd1
+ vccd1 vccd1 _303_ sky130_fd_sc_hd__mux2_1
X_562_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.d sky130_fd_sc_hd__clkinv_2
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_829_ CIRCUIT_2223.MEMORY_21.s_currentState vssd1 vssd1 vccd1 vccd1 _110_ sky130_fd_sc_hd__clkinv_2
XFILLER_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_614_ _289_ _290_ vssd1 vssd1 vccd1 vccd1 _294_ sky130_fd_sc_hd__and2b_1
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_476_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2
+ vssd1 vssd1 vccd1 vccd1 _238_ sky130_fd_sc_hd__nand2_1
X_545_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.d sky130_fd_sc_hd__clkinv_2
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__962__D net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_459_ CIRCUIT_2223.GATES_1.input1\[3\] CIRCUIT_2223.GATES_1.input1\[2\] net1 net2
+ vssd1 vssd1 vccd1 vccd1 _232_ sky130_fd_sc_hd__and4b_1
X_528_ _268_ _274_ _279_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_27.result
+ sky130_fd_sc_hd__nor3_1
XFILLER_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__510__A _191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_475__1 clknet_1_0__leaf__195_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__inv_2
XFILLER_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_862_ net16 CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState _006_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_18.s_currentState sky130_fd_sc_hd__dfstp_1
X_931_ net19 _157_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_12.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_793_ net3 CIRCUIT_2223.tone_generator_2_1.GATES_8.input2 _364_ vssd1 vssd1 vccd1
+ vccd1 _365_ sky130_fd_sc_hd__mux2_1
XFILLER_19_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__236_ clknet_0__236_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__236_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_845_ net16 CIRCUIT_2223.tone_generator_1.MEMORY_20.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_4.s_currentState sky130_fd_sc_hd__dfxtp_1
X_776_ _361_ vssd1 vssd1 vccd1 vccd1 _161_ sky130_fd_sc_hd__clkbuf_1
X_914_ net22 _152_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_7.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_630_ _259_ _301_ vssd1 vssd1 vccd1 vccd1 _302_ sky130_fd_sc_hd__nand2_1
X_492_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_34.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_13.input2
+ vssd1 vssd1 vccd1 vccd1 _254_ sky130_fd_sc_hd__xor2_1
X_561_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_31.d sky130_fd_sc_hd__clkinv_2
XFILLER_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_759_ _186_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2 _350_
+ vssd1 vssd1 vccd1 vccd1 _352_ sky130_fd_sc_hd__mux2_1
X_828_ CIRCUIT_2223.MEMORY_22.s_currentState vssd1 vssd1 vccd1 vccd1 _108_ sky130_fd_sc_hd__clkinv_2
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_613_ _291_ _292_ vssd1 vssd1 vccd1 vccd1 _293_ sky130_fd_sc_hd__and2b_1
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_544_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_36.d sky130_fd_sc_hd__clkinv_2
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_input5_A io_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__508__A _191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_527_ _275_ _276_ _277_ _278_ vssd1 vssd1 vccd1 vccd1 _279_ sky130_fd_sc_hd__or4_1
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_458_ _220_ _226_ _231_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_27.result
+ sky130_fd_sc_hd__nor3_1
X_389_ net2 net1 CIRCUIT_2223.GATES_1.input1\[0\] CIRCUIT_2223.GATES_1.input1\[1\]
+ vssd1 vssd1 vccd1 vccd1 _180_ sky130_fd_sc_hd__and4_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_475__2 clknet_1_1__leaf__195_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__inv_2
XFILLER_42_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__726__A0 _184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_930_ net19 _156_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_1.GATES_11.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_861_ net17 CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState _005_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_17.s_currentState sky130_fd_sc_hd__dfrtp_1
X_792_ _233_ _326_ vssd1 vssd1 vccd1 vccd1 _364_ sky130_fd_sc_hd__nand2_1
XFILLER_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__431__A _000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_913_ net22 _151_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_17.input2
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__235_ clknet_0__235_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__235_
+ sky130_fd_sc_hd__clkbuf_16
X_844_ clknet_1_1__leaf_clk _129_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.CLK sky130_fd_sc_hd__dfxtp_1
X_775_ net4 CIRCUIT_2223.tone_generator_2_1.GATES_16.input2 _359_ vssd1 vssd1 vccd1
+ vccd1 _361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_560_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.s_currentState vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_30.d sky130_fd_sc_hd__clkinv_2
XFILLER_44_98 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_491_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_32.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_11.input2
+ vssd1 vssd1 vccd1 vccd1 _253_ sky130_fd_sc_hd__xor2_1
XFILLER_5_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_758_ _351_ vssd1 vssd1 vccd1 vccd1 _153_ sky130_fd_sc_hd__clkbuf_1
X_827_ _179_ vssd1 vssd1 vccd1 vccd1 _106_ sky130_fd_sc_hd__inv_2
X_689_ _333_ vssd1 vssd1 vccd1 vccd1 _138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_612_ CIRCUIT_2223.GATES_5.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState
+ CIRCUIT_2223.GATES_4.input1\[3\] CIRCUIT_2223.s_logisimNet48 vssd1 vssd1 vccd1 vccd1
+ _292_ sky130_fd_sc_hd__a22o_1
X_543_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d sky130_fd_sc_hd__clkinv_2
X_474_ _237_ clknet_1_0__leaf__236_ vssd1 vssd1 vccd1 vccd1 _054_ sky130_fd_sc_hd__xnor2_2
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_526_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_16.input2
+ vssd1 vssd1 vccd1 vccd1 _278_ sky130_fd_sc_hd__xor2_1
XANTENNA__434__A _000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_457_ _227_ _228_ _229_ _230_ vssd1 vssd1 vccd1 vccd1 _231_ sky130_fd_sc_hd__or4_1
X_388_ _179_ vssd1 vssd1 vccd1 vccd1 _102_ sky130_fd_sc_hd__inv_2
XFILLER_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__671__A0 _186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_509_ _191_ clknet_1_1__leaf__263_ vssd1 vssd1 vccd1 vccd1 _034_ sky130_fd_sc_hd__xnor2_2
XFILLER_9_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_791_ CIRCUIT_2223.tone_generator_2_2.MEMORY_37.s_currentState vssd1 vssd1 vccd1
+ vccd1 _095_ sky130_fd_sc_hd__clkinv_2
X_860_ net17 CIRCUIT_2223.tone_generator_1.MEMORY_15.s_currentState _004_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.tone_generator_1.MEMORY_16.s_currentState sky130_fd_sc_hd__dfstp_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__635__A0 _184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__532__A _000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout19_A net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_843_ clknet_1_1__leaf_clk _128_ vssd1 vssd1 vccd1 vccd1 slow_clock\[6\] sky130_fd_sc_hd__dfxtp_1
X_912_ net22 _150_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2
+ sky130_fd_sc_hd__dfxtp_1
X_774_ _360_ vssd1 vssd1 vccd1 vccd1 _160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_490_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_29.s_currentState CIRCUIT_2223.triangle_wave_generator_1.GATES_8.input2
+ vssd1 vssd1 vccd1 vccd1 _252_ sky130_fd_sc_hd__xor2_1
X_826_ net17 vssd1 vssd1 vccd1 vccd1 _105_ sky130_fd_sc_hd__clkinv_2
X_757_ _188_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_8.input2 _350_
+ vssd1 vssd1 vccd1 vccd1 _351_ sky130_fd_sc_hd__mux2_1
X_688_ _188_ CIRCUIT_2223.GATES_1.input1\[0\] _332_ vssd1 vssd1 vccd1 vccd1 _333_
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_611_ CIRCUIT_2223.s_logisimNet48 CIRCUIT_2223.GATES_5.input2 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_40.s_currentState
+ CIRCUIT_2223.GATES_4.input1\[3\] vssd1 vssd1 vccd1 vccd1 _291_ sky130_fd_sc_hd__and4_1
X_542_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.clock
+ sky130_fd_sc_hd__clkinv_2
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_473_ _237_ clknet_1_0__leaf__236_ vssd1 vssd1 vccd1 vccd1 _056_ sky130_fd_sc_hd__xnor2_2
XFILLER_4_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_809_ net3 CIRCUIT_2223.tone_generator_2_2.GATES_15.input2 _373_ vssd1 vssd1 vccd1
+ vccd1 _374_ sky130_fd_sc_hd__mux2_1
XFILLER_35_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__540__A _215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_456_ CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_14.input2
+ vssd1 vssd1 vccd1 vccd1 _230_ sky130_fd_sc_hd__xor2_1
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_525_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_35.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2
+ vssd1 vssd1 vccd1 vccd1 _277_ sky130_fd_sc_hd__xor2_1
XFILLER_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_387_ _179_ vssd1 vssd1 vccd1 vccd1 _104_ sky130_fd_sc_hd__inv_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_439_ _214_ clknet_1_1__leaf__213_ vssd1 vssd1 vccd1 vccd1 _077_ sky130_fd_sc_hd__xor2_2
XFILLER_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_508_ _191_ clknet_1_1__leaf__263_ vssd1 vssd1 vccd1 vccd1 _036_ sky130_fd_sc_hd__xnor2_2
XFILLER_36_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_790_ CIRCUIT_2223.tone_generator_2_2.MEMORY_36.s_currentState vssd1 vssd1 vccd1
+ vccd1 _093_ sky130_fd_sc_hd__clkinv_2
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_842_ clknet_1_0__leaf_clk _127_ vssd1 vssd1 vccd1 vccd1 slow_clock\[5\] sky130_fd_sc_hd__dfxtp_1
X_911_ net22 _149_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_773_ net3 CIRCUIT_2223.tone_generator_2_1.GATES_15.input2 _359_ vssd1 vssd1 vccd1
+ vccd1 _360_ sky130_fd_sc_hd__mux2_1
XFILLER_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_756_ _181_ _193_ vssd1 vssd1 vccd1 vccd1 _350_ sky130_fd_sc_hd__nand2_1
X_825_ CIRCUIT_2223.MEMORY_25.s_currentState vssd1 vssd1 vccd1 vccd1 _103_ sky130_fd_sc_hd__clkinv_2
X_687_ net1 net2 vssd1 vssd1 vccd1 vccd1 _332_ sky130_fd_sc_hd__or2b_1
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_610_ _289_ _290_ vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__xnor2_1
XFILLER_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_541_ _215_ clknet_1_1__leaf__282_ vssd1 vssd1 vccd1 vccd1 _009_ sky130_fd_sc_hd__xor2_2
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_472_ _237_ clknet_1_0__leaf__236_ vssd1 vssd1 vccd1 vccd1 _058_ sky130_fd_sc_hd__xnor2_2
XANTENNA__538__A _215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_808_ _192_ _326_ vssd1 vssd1 vccd1 vccd1 _373_ sky130_fd_sc_hd__nand2_2
X_739_ _186_ CIRCUIT_2223.triangle_wave_generator_1.GATES_16.input2 _345_ vssd1 vssd1
+ vccd1 vccd1 _347_ sky130_fd_sc_hd__mux2_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_524_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_30.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_9.input2
+ vssd1 vssd1 vccd1 vccd1 _276_ sky130_fd_sc_hd__xor2_1
X_455_ CIRCUIT_2223.tone_generator_2_1.MEMORY_28.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_7.input2
+ vssd1 vssd1 vccd1 vccd1 _229_ sky130_fd_sc_hd__xor2_1
X_386_ _179_ vssd1 vssd1 vccd1 vccd1 _107_ sky130_fd_sc_hd__inv_2
XANTENNA__856__SET_B _000_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input3_A io_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_438_ _214_ clknet_1_1__leaf__213_ vssd1 vssd1 vccd1 vccd1 _079_ sky130_fd_sc_hd__xor2_2
X_507_ _191_ clknet_1_0__leaf__263_ vssd1 vssd1 vccd1 vccd1 _039_ sky130_fd_sc_hd__xnor2_2
XFILLER_9_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_841_ clknet_1_0__leaf_clk _126_ vssd1 vssd1 vccd1 vccd1 slow_clock\[4\] sky130_fd_sc_hd__dfxtp_1
X_910_ net23 _148_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2
+ sky130_fd_sc_hd__dfxtp_1
X_772_ _233_ _301_ vssd1 vssd1 vccd1 vccd1 _359_ sky130_fd_sc_hd__nand2_2
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout24_A CIRCUIT_2223.CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_755_ CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState vssd1 vssd1 vccd1
+ vccd1 _074_ sky130_fd_sc_hd__clkinv_2
X_824_ _320_ _306_ vssd1 vssd1 vccd1 vccd1 _101_ sky130_fd_sc_hd__nand2_1
X_686_ _331_ vssd1 vssd1 vccd1 vccd1 _137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__955__CLK net21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_540_ _215_ clknet_1_1__leaf__282_ vssd1 vssd1 vccd1 vccd1 _011_ sky130_fd_sc_hd__xor2_2
XFILLER_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_471_ _237_ clknet_1_1__leaf__236_ vssd1 vssd1 vccd1 vccd1 _060_ sky130_fd_sc_hd__xnor2_2
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_807_ _372_ vssd1 vssd1 vccd1 vccd1 _170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_738_ _346_ vssd1 vssd1 vccd1 vccd1 _149_ sky130_fd_sc_hd__clkbuf_1
X_669_ _188_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_15.input2 _321_
+ vssd1 vssd1 vccd1 vccd1 _322_ sky130_fd_sc_hd__mux2_1
XANTENNA__464__A _215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__692__A0 _184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__821__B _319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__683__A0 _184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_523_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_28.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_7.input2
+ vssd1 vssd1 vccd1 vccd1 _275_ sky130_fd_sc_hd__xor2_1
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_454_ CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_16.input2
+ vssd1 vssd1 vccd1 vccd1 _228_ sky130_fd_sc_hd__xor2_1
X_385_ _179_ vssd1 vssd1 vccd1 vccd1 _109_ sky130_fd_sc_hd__inv_2
XFILLER_23_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__656__B1 _306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_506_ _191_ clknet_1_0__leaf__263_ vssd1 vssd1 vccd1 vccd1 _041_ sky130_fd_sc_hd__xnor2_2
X_437_ _214_ clknet_1_1__leaf__213_ vssd1 vssd1 vccd1 vccd1 _081_ sky130_fd_sc_hd__xor2_2
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_840_ clknet_1_0__leaf_clk _125_ vssd1 vssd1 vccd1 vccd1 slow_clock\[3\] sky130_fd_sc_hd__dfxtp_1
X_771_ _358_ vssd1 vssd1 vccd1 vccd1 _159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_969_ net26 CIRCUIT_2223.MEMORY_24.d _106_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_24.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__824__B _306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_823_ _320_ _306_ vssd1 vssd1 vccd1 vccd1 _100_ sky130_fd_sc_hd__nand2_1
X_754_ CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState vssd1 vssd1 vccd1
+ vccd1 _072_ sky130_fd_sc_hd__clkinv_2
X_685_ net6 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_14.input2 _327_
+ vssd1 vssd1 vccd1 vccd1 _331_ sky130_fd_sc_hd__mux2_1
XFILLER_34_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_470_ _237_ clknet_1_1__leaf__236_ vssd1 vssd1 vccd1 vccd1 _063_ sky130_fd_sc_hd__xnor2_2
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_806_ net6 CIRCUIT_2223.tone_generator_2_2.GATES_14.input2 _368_ vssd1 vssd1 vccd1
+ vccd1 _372_ sky130_fd_sc_hd__mux2_1
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_737_ _188_ CIRCUIT_2223.triangle_wave_generator_1.GATES_15.input2 _345_ vssd1 vssd1
+ vccd1 vccd1 _346_ sky130_fd_sc_hd__mux2_1
X_668_ _180_ _259_ vssd1 vssd1 vccd1 vccd1 _321_ sky130_fd_sc_hd__nand2_2
X_599_ CIRCUIT_2223.MEMORY_19.s_currentState vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_19.d
+ sky130_fd_sc_hd__clkinv_2
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_453_ CIRCUIT_2223.tone_generator_2_1.MEMORY_30.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_9.input2
+ vssd1 vssd1 vccd1 vccd1 _227_ sky130_fd_sc_hd__xor2_1
XFILLER_17_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_522_ _269_ _270_ _271_ _272_ _273_ vssd1 vssd1 vccd1 vccd1 _274_ sky130_fd_sc_hd__a221o_1
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_384_ _179_ vssd1 vssd1 vccd1 vccd1 _111_ sky130_fd_sc_hd__inv_2
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_436_ _214_ clknet_1_1__leaf__213_ vssd1 vssd1 vccd1 vccd1 _084_ sky130_fd_sc_hd__xor2_2
X_505_ _237_ clknet_1_0__leaf__263_ vssd1 vssd1 vccd1 vccd1 _043_ sky130_fd_sc_hd__xnor2_2
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_419_ CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_8.input2
+ vssd1 vssd1 vccd1 vccd1 _204_ sky130_fd_sc_hd__nand2_1
XFILLER_24_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__795__A0 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_770_ net6 CIRCUIT_2223.tone_generator_2_1.GATES_14.input2 _354_ vssd1 vssd1 vccd1
+ vccd1 _358_ sky130_fd_sc_hd__mux2_1
X_968_ _105_ CIRCUIT_2223.MEMORY_25.d _104_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_25.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_899_ _050_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_28.clock _049_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_38.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__777__A0 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__213_ clknet_0__213_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__213_
+ sky130_fd_sc_hd__clkbuf_16
X_822_ _320_ _319_ vssd1 vssd1 vccd1 vccd1 _099_ sky130_fd_sc_hd__nand2_1
XANTENNA__768__A0 _184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_753_ CIRCUIT_2223.tone_generator_2_1.MEMORY_35.s_currentState vssd1 vssd1 vccd1
+ vccd1 _070_ sky130_fd_sc_hd__clkinv_2
XFILLER_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_684_ _330_ vssd1 vssd1 vccd1 vccd1 _136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__759__A0 _186_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__660__B _319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_805_ _371_ vssd1 vssd1 vccd1 vccd1 _169_ sky130_fd_sc_hd__clkbuf_1
X_736_ _193_ _259_ vssd1 vssd1 vccd1 vccd1 _345_ sky130_fd_sc_hd__nand2_1
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_667_ _320_ _319_ vssd1 vssd1 vccd1 vccd1 _008_ sky130_fd_sc_hd__nand2_1
X_598_ CIRCUIT_2223.MEMORY_20.s_currentState vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_20.d
+ sky130_fd_sc_hd__clkinv_2
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__390__B net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_452_ _221_ _222_ _223_ _224_ _225_ vssd1 vssd1 vccd1 vccd1 _226_ sky130_fd_sc_hd__a221o_1
X_383_ _179_ vssd1 vssd1 vccd1 vccd1 _113_ sky130_fd_sc_hd__inv_2
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_521_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_38.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_17.input2
+ vssd1 vssd1 vccd1 vccd1 _273_ sky130_fd_sc_hd__xor2_1
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_719_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_42.s_currentState vssd1 vssd1
+ vccd1 vccd1 _052_ sky130_fd_sc_hd__clkinv_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__459__C net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_504_ _237_ clknet_1_0__leaf__263_ vssd1 vssd1 vccd1 vccd1 _045_ sky130_fd_sc_hd__xnor2_2
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_435_ _191_ vssd1 vssd1 vccd1 vccd1 _214_ sky130_fd_sc_hd__buf_8
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input1_A io_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_418_ CIRCUIT_2223.tone_generator_2_2.MEMORY_29.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_8.input2
+ vssd1 vssd1 vccd1 vccd1 _203_ sky130_fd_sc_hd__or2_1
XANTENNA__663__B _319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_898_ _048_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.d _047_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_967_ _103_ CIRCUIT_2223.MEMORY_18.clock _102_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_26.s_currentState
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__212_ clknet_0__212_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__212_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_821_ _320_ _319_ vssd1 vssd1 vccd1 vccd1 _098_ sky130_fd_sc_hd__nand2_1
X_752_ CIRCUIT_2223.tone_generator_2_1.MEMORY_34.s_currentState vssd1 vssd1 vccd1
+ vccd1 _068_ sky130_fd_sc_hd__clkinv_2
X_683_ _184_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_13.input2 _327_
+ vssd1 vssd1 vccd1 vccd1 _330_ sky130_fd_sc_hd__mux2_1
XFILLER_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_804_ net5 CIRCUIT_2223.tone_generator_2_2.GATES_13.input2 _368_ vssd1 vssd1 vccd1
+ vccd1 _371_ sky130_fd_sc_hd__mux2_1
XFILLER_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_735_ _344_ vssd1 vssd1 vccd1 vccd1 _148_ sky130_fd_sc_hd__clkbuf_1
X_666_ _320_ _319_ vssd1 vssd1 vccd1 vccd1 _007_ sky130_fd_sc_hd__nand2_1
X_597_ CIRCUIT_2223.MEMORY_21.s_currentState vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_21.d
+ sky130_fd_sc_hd__clkinv_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_520_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_32.s_currentState CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_11.input2
+ vssd1 vssd1 vccd1 vccd1 _272_ sky130_fd_sc_hd__or2_1
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_451_ CIRCUIT_2223.tone_generator_2_1.MEMORY_29.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_8.input2
+ vssd1 vssd1 vccd1 vccd1 _225_ sky130_fd_sc_hd__xor2_1
X_382_ _179_ vssd1 vssd1 vccd1 vccd1 _115_ sky130_fd_sc_hd__inv_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_718_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_41.s_currentState vssd1 vssd1
+ vccd1 vccd1 _051_ sky130_fd_sc_hd__clkinv_2
X_649_ slow_clock\[4\] _310_ _313_ vssd1 vssd1 vccd1 vccd1 _126_ sky130_fd_sc_hd__o21a_1
XFILLER_36_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__666__B _319_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__813__A0 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_503_ _237_ clknet_1_0__leaf__263_ vssd1 vssd1 vccd1 vccd1 _047_ sky130_fd_sc_hd__xnor2_2
X_434_ _000_ clknet_1_0__leaf__213_ vssd1 vssd1 vccd1 vccd1 _086_ sky130_fd_sc_hd__xor2_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__804__A0 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_417_ CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_17.input2
+ vssd1 vssd1 vccd1 vccd1 _202_ sky130_fd_sc_hd__nand2_1
XFILLER_23_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_966_ net20 _178_ _101_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.s_logisimNet48 sky130_fd_sc_hd__dfrtp_2
X_897_ _046_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.d _045_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_820_ _379_ vssd1 vssd1 vccd1 vccd1 _097_ sky130_fd_sc_hd__clkbuf_1
X_751_ CIRCUIT_2223.tone_generator_2_1.MEMORY_33.s_currentState vssd1 vssd1 vccd1
+ vccd1 _066_ sky130_fd_sc_hd__clkinv_2
XFILLER_18_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_682_ _329_ vssd1 vssd1 vccd1 vccd1 _135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_18_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_949_ CIRCUIT_2223.tone_generator_2_2.GATES_27.result CIRCUIT_2223.tone_generator_2_2.MEMORY_39.d
+ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_39.s_currentState
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__392__A0 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_803_ _370_ vssd1 vssd1 vccd1 vccd1 _168_ sky130_fd_sc_hd__clkbuf_1
X_665_ _320_ _319_ vssd1 vssd1 vccd1 vccd1 _006_ sky130_fd_sc_hd__nand2_1
XFILLER_28_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_734_ net6 CIRCUIT_2223.triangle_wave_generator_1.GATES_14.input2 _260_ vssd1 vssd1
+ vccd1 vccd1 _344_ sky130_fd_sc_hd__mux2_1
X_596_ CIRCUIT_2223.MEMORY_22.s_currentState vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_22.d
+ sky130_fd_sc_hd__clkinv_2
XFILLER_6_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_450_ CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState CIRCUIT_2223.tone_generator_2_1.GATES_11.input2
+ vssd1 vssd1 vccd1 vccd1 _224_ sky130_fd_sc_hd__or2_1
X_381_ net20 vssd1 vssd1 vccd1 vccd1 _179_ sky130_fd_sc_hd__clkbuf_4
XFILLER_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_648_ _306_ _312_ vssd1 vssd1 vccd1 vccd1 _313_ sky130_fd_sc_hd__nor2_1
X_717_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_37.s_currentState vssd1 vssd1
+ vccd1 vccd1 _050_ sky130_fd_sc_hd__clkinv_2
X_579_ CIRCUIT_2223.tone_generator_2_1.MEMORY_37.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_37.d sky130_fd_sc_hd__clkinv_2
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_433_ _000_ clknet_1_0__leaf__213_ vssd1 vssd1 vccd1 vccd1 _088_ sky130_fd_sc_hd__xor2_2
X_502_ _215_ clknet_1_1__leaf__263_ vssd1 vssd1 vccd1 vccd1 _049_ sky130_fd_sc_hd__xnor2_2
XFILLER_26_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_416_ CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState CIRCUIT_2223.tone_generator_2_2.GATES_17.input2
+ vssd1 vssd1 vccd1 vccd1 _201_ sky130_fd_sc_hd__or2_1
XFILLER_18_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__722__A0 _188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_965_ net20 _177_ _100_ vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.GATES_5.input2 sky130_fd_sc_hd__dfrtp_2
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_896_ _044_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.d _043_ vssd1 vssd1
+ vccd1 vccd1 CIRCUIT_2223.triangle_wave_generator_1.MEMORY_35.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_750_ CIRCUIT_2223.tone_generator_2_1.MEMORY_32.s_currentState vssd1 vssd1 vccd1
+ vccd1 _064_ sky130_fd_sc_hd__clkinv_2
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_681_ _186_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.GATES_12.input2 _327_
+ vssd1 vssd1 vccd1 vccd1 _329_ sky130_fd_sc_hd__mux2_1
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_948_ _095_ CIRCUIT_2223.tone_generator_2_2.MEMORY_28.clock _094_ vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_2.MEMORY_38.s_currentState sky130_fd_sc_hd__dfrtp_1
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_879_ _012_ CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.d _011_ vssd1
+ vssd1 vccd1 vccd1 CIRCUIT_2223.tone_generator_1.tone_generator_2_1.MEMORY_37.s_currentState
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_802_ net4 CIRCUIT_2223.tone_generator_2_2.GATES_12.input2 _368_ vssd1 vssd1 vccd1
+ vccd1 _370_ sky130_fd_sc_hd__mux2_1
XFILLER_29_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_664_ _320_ _319_ vssd1 vssd1 vccd1 vccd1 _005_ sky130_fd_sc_hd__nand2_1
X_733_ _343_ vssd1 vssd1 vccd1 vccd1 _147_ sky130_fd_sc_hd__clkbuf_1
X_595_ net17 vssd1 vssd1 vccd1 vccd1 CIRCUIT_2223.MEMORY_24.d sky130_fd_sc_hd__clkinv_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_380_ net18 vssd1 vssd1 vccd1 vccd1 _117_ sky130_fd_sc_hd__inv_2
X_716_ CIRCUIT_2223.triangle_wave_generator_1.MEMORY_36.s_currentState vssd1 vssd1
+ vccd1 vccd1 _048_ sky130_fd_sc_hd__clkinv_2
X_647_ slow_clock\[4\] _310_ vssd1 vssd1 vccd1 vccd1 _312_ sky130_fd_sc_hd__and2_1
X_578_ CIRCUIT_2223.tone_generator_2_1.MEMORY_36.s_currentState vssd1 vssd1 vccd1
+ vccd1 CIRCUIT_2223.tone_generator_2_1.MEMORY_36.d sky130_fd_sc_hd__clkinv_2
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

