magic
tech sky130B
magscale 1 2
timestamp 1680007705
<< obsli1 >>
rect 1104 2159 68816 67473
<< obsm1 >>
rect 934 2128 69078 67504
<< obsm2 >>
rect 938 2139 69074 67493
<< metal3 >>
rect 0 62568 800 62688
rect 69200 60936 70000 61056
rect 0 48696 800 48816
rect 69200 43528 70000 43648
rect 0 34824 800 34944
rect 69200 26120 70000 26240
rect 0 20952 800 21072
rect 69200 8712 70000 8832
rect 0 7080 800 7200
<< obsm3 >>
rect 800 62768 69200 67489
rect 880 62488 69200 62768
rect 800 61136 69200 62488
rect 800 60856 69120 61136
rect 800 48896 69200 60856
rect 880 48616 69200 48896
rect 800 43728 69200 48616
rect 800 43448 69120 43728
rect 800 35024 69200 43448
rect 880 34744 69200 35024
rect 800 26320 69200 34744
rect 800 26040 69120 26320
rect 800 21152 69200 26040
rect 880 20872 69200 21152
rect 800 8912 69200 20872
rect 800 8632 69120 8912
rect 800 7280 69200 8632
rect 880 7000 69200 7280
rect 800 2143 69200 7000
<< metal4 >>
rect 4208 2128 4528 67504
rect 19568 2128 19888 67504
rect 34928 2128 35248 67504
rect 50288 2128 50608 67504
rect 65648 2128 65968 67504
<< obsm4 >>
rect 7235 3979 19488 57357
rect 19968 3979 34848 57357
rect 35328 3979 50208 57357
rect 50688 3979 65568 57357
rect 66048 3979 67101 57357
<< labels >>
rlabel metal3 s 0 48696 800 48816 6 clk
port 1 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 io_in[0]
port 2 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 69200 8712 70000 8832 6 io_out[0]
port 5 nsew signal output
rlabel metal3 s 69200 26120 70000 26240 6 io_out[1]
port 6 nsew signal output
rlabel metal3 s 69200 43528 70000 43648 6 io_out[2]
port 7 nsew signal output
rlabel metal3 s 69200 60936 70000 61056 6 io_out[3]
port 8 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 rst
port 9 nsew signal input
rlabel metal4 s 4208 2128 4528 67504 6 vccd1
port 10 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 67504 6 vccd1
port 10 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 67504 6 vccd1
port 10 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 67504 6 vssd1
port 11 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 67504 6 vssd1
port 11 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 70000 70000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11873386
string GDS_FILE /run/media/tholin/e6042058-84c8-448b-be8a-b40bc065b34b/TMBoC/openlane/PositUnit/runs/23_03_28_14_44/results/signoff/posit_unit.magic.gds
string GDS_START 1534712
<< end >>

